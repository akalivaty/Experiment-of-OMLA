//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936;
  XNOR2_X1  g000(.A(G169gat), .B(G197gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OR3_X1    g010(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT92), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT93), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n214), .A2(KEYINPUT92), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(KEYINPUT92), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT93), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n213), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OR3_X1    g022(.A1(new_n209), .A2(KEYINPUT94), .A3(new_n210), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n215), .A2(new_n212), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT94), .B1(new_n209), .B2(new_n210), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n209), .A2(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT17), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(G1gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G1gat), .B2(new_n231), .ZN(new_n234));
  INV_X1    g033(.A(G8gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n236), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n229), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n238), .B(new_n229), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n240), .B(KEYINPUT13), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(new_n237), .B2(new_n241), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n208), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT96), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n237), .A2(new_n241), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n247), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n253), .A2(new_n245), .A3(new_n242), .A4(new_n207), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(KEYINPUT96), .B(new_n208), .C1(new_n246), .C2(new_n249), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT89), .ZN(new_n258));
  XOR2_X1   g057(.A(G127gat), .B(G134gat), .Z(new_n259));
  INV_X1    g058(.A(G113gat), .ZN(new_n260));
  INV_X1    g059(.A(G120gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G113gat), .A2(G120gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n259), .A2(new_n264), .A3(KEYINPUT1), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G113gat), .A2(G120gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(G113gat), .A2(G120gat), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT68), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n262), .A2(new_n270), .A3(new_n263), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n273), .A2(KEYINPUT69), .A3(new_n259), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT69), .B1(new_n273), .B2(new_n259), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n266), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT24), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(G183gat), .A3(G190gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G183gat), .B(G190gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n278), .ZN(new_n281));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT23), .ZN(new_n283));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT23), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n277), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n281), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n283), .A2(KEYINPUT25), .A3(new_n286), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n291), .A2(new_n292), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(KEYINPUT64), .B(new_n277), .C1(new_n281), .C2(new_n287), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n283), .A4(new_n286), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT66), .B1(new_n300), .B2(new_n281), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n290), .A2(new_n298), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n284), .ZN(new_n306));
  INV_X1    g105(.A(G183gat), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT27), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G183gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(KEYINPUT27), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n313), .A2(KEYINPUT28), .A3(new_n308), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(KEYINPUT67), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  AOI21_X1  g115(.A(G190gat), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT28), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  OAI221_X1 g117(.A(new_n306), .B1(new_n307), .B2(new_n308), .C1(new_n314), .C2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n276), .B1(new_n302), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n276), .A3(new_n319), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n321), .A2(G227gat), .A3(G233gat), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT32), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT33), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G15gat), .B(G43gat), .Z(new_n327));
  XNOR2_X1  g126(.A(G71gat), .B(G99gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n322), .ZN(new_n331));
  INV_X1    g130(.A(G227gat), .ZN(new_n332));
  INV_X1    g131(.A(G233gat), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n331), .A2(new_n320), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT34), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI221_X1 g135(.A(KEYINPUT34), .B1(new_n332), .B2(new_n333), .C1(new_n331), .C2(new_n320), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n329), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n323), .B(KEYINPUT32), .C1(new_n325), .C2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n330), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n330), .B2(new_n340), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n258), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n330), .A2(new_n340), .ZN(new_n345));
  INV_X1    g144(.A(new_n338), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(KEYINPUT89), .A3(new_n341), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n350), .A2(KEYINPUT72), .ZN(new_n351));
  XNOR2_X1  g150(.A(G197gat), .B(G204gat), .ZN(new_n352));
  AND2_X1   g151(.A1(G211gat), .A2(G218gat), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n352), .B1(KEYINPUT22), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n351), .B(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(KEYINPUT29), .ZN(new_n356));
  INV_X1    g155(.A(G141gat), .ZN(new_n357));
  INV_X1    g156(.A(G148gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G141gat), .A2(G148gat), .ZN(new_n360));
  AND2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n359), .B(new_n360), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G162gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT77), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G162gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G155gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n369), .B2(KEYINPUT2), .ZN(new_n370));
  NAND2_X1  g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT2), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(new_n359), .A3(new_n360), .ZN(new_n373));
  INV_X1    g172(.A(G155gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n364), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n371), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT76), .B1(new_n361), .B2(new_n362), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n373), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n356), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(new_n370), .B2(new_n379), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(KEYINPUT83), .A3(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(G228gat), .A2(G233gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n375), .A2(new_n371), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n359), .A2(new_n360), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n374), .B1(new_n365), .B2(new_n367), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT2), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n378), .A3(new_n377), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n355), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n397), .B(new_n381), .C1(new_n356), .C2(KEYINPUT3), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n384), .A2(new_n385), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n370), .B2(new_n379), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n390), .A2(KEYINPUT79), .A3(new_n392), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT29), .B1(new_n354), .B2(new_n350), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n350), .B2(new_n354), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n406), .A2(KEYINPUT82), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT3), .B1(new_n406), .B2(KEYINPUT82), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n355), .B2(new_n395), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n399), .B1(new_n410), .B2(new_n385), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G22gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  MUX2_X1   g215(.A(G22gat), .B(new_n413), .S(new_n416), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n411), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n349), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n421), .B(KEYINPUT73), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n302), .A2(new_n319), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(new_n394), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n302), .B2(new_n319), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n355), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n426), .ZN(new_n428));
  INV_X1    g227(.A(new_n355), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(new_n302), .B2(new_n319), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n428), .B(new_n429), .C1(new_n430), .C2(new_n423), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(G64gat), .ZN(new_n434));
  INV_X1    g233(.A(G92gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(KEYINPUT74), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT30), .B1(new_n432), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n432), .A2(new_n441), .A3(KEYINPUT30), .A4(new_n436), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n427), .A2(new_n431), .A3(KEYINPUT30), .A4(new_n436), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT75), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n437), .A2(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT90), .B(KEYINPUT35), .Z(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G1gat), .B(G29gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(KEYINPUT0), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(G57gat), .ZN(new_n450));
  INV_X1    g249(.A(G85gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT85), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n450), .B(G85gat), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT5), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n276), .B(new_n381), .ZN(new_n458));
  NAND2_X1  g257(.A1(G225gat), .A2(G233gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n273), .A2(new_n259), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n273), .A2(KEYINPUT69), .A3(new_n259), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n265), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n383), .A2(new_n393), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n276), .A2(KEYINPUT78), .A3(new_n393), .A4(new_n383), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT4), .B1(new_n403), .B2(new_n276), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT4), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n468), .A2(new_n474), .A3(new_n380), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n476), .A3(new_n459), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT80), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT80), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n476), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n462), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n404), .A2(new_n468), .A3(new_n474), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT4), .B1(new_n276), .B2(new_n381), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n479), .A2(new_n485), .A3(new_n457), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n453), .B(new_n456), .C1(new_n482), .C2(new_n487), .ZN(new_n488));
  AND4_X1   g287(.A1(new_n480), .A2(new_n472), .A3(new_n476), .A4(new_n459), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n480), .B1(new_n479), .B2(new_n476), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n461), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n452), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT6), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n452), .B1(new_n491), .B2(new_n486), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n488), .A2(new_n494), .B1(new_n495), .B2(KEYINPUT6), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n447), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n420), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT6), .B(new_n454), .C1(new_n482), .C2(new_n487), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n482), .B2(new_n492), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n501), .B2(new_n495), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT81), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n502), .A2(new_n503), .A3(new_n445), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n502), .B2(new_n445), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n347), .A2(KEYINPUT70), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT70), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n343), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n506), .A2(new_n508), .A3(new_n418), .A4(new_n341), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n498), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n427), .A2(new_n431), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT37), .ZN(new_n515));
  INV_X1    g314(.A(new_n436), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n514), .B2(KEYINPUT37), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT37), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n427), .A2(new_n431), .A3(KEYINPUT87), .A4(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n517), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT38), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n521), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n516), .A3(new_n515), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(KEYINPUT88), .A3(KEYINPUT38), .ZN(new_n527));
  AOI211_X1 g326(.A(KEYINPUT38), .B(new_n439), .C1(new_n514), .C2(KEYINPUT37), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n525), .A2(new_n528), .B1(new_n436), .B2(new_n432), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n524), .A2(new_n527), .A3(new_n496), .A4(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT86), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n453), .A2(new_n456), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n459), .B1(new_n485), .B2(new_n472), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT39), .B1(new_n458), .B2(new_n460), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI211_X1 g334(.A(KEYINPUT39), .B(new_n459), .C1(new_n485), .C2(new_n472), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n531), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT40), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT40), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n531), .B(new_n539), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n538), .A2(new_n488), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n445), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n419), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n530), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n419), .B1(new_n504), .B2(new_n505), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n341), .A2(KEYINPUT36), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n506), .A2(new_n546), .A3(new_n508), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT71), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n506), .A2(new_n546), .A3(new_n549), .A4(new_n508), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT36), .B1(new_n347), .B2(new_n341), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n544), .A2(new_n545), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n257), .B1(new_n512), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT101), .B(G183gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT100), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n563));
  INV_X1    g362(.A(G57gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(G64gat), .ZN(new_n565));
  INV_X1    g364(.A(G64gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(G57gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n563), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(new_n569), .B2(new_n568), .ZN(new_n571));
  XOR2_X1   g370(.A(G71gat), .B(G78gat), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n563), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n572), .B1(KEYINPUT99), .B2(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n565), .A2(KEYINPUT98), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n565), .A2(KEYINPUT98), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n567), .A3(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n574), .A2(KEYINPUT99), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G127gat), .B(G155gat), .ZN(new_n582));
  OR3_X1    g381(.A1(new_n581), .A2(KEYINPUT21), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G211gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n581), .B2(KEYINPUT21), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n584), .B1(new_n583), .B2(new_n585), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n562), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n238), .B1(new_n581), .B2(KEYINPUT21), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n583), .A2(new_n585), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(G211gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n561), .A3(new_n586), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n589), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n591), .B1(new_n589), .B2(new_n594), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n557), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(new_n556), .A3(new_n595), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT7), .ZN(new_n603));
  INV_X1    g402(.A(G99gat), .ZN(new_n604));
  INV_X1    g403(.A(G106gat), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT8), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT104), .B(G85gat), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n603), .B(new_n606), .C1(G92gat), .C2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G99gat), .B(G106gat), .Z(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT105), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n230), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n610), .A2(new_n611), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n617), .B2(new_n229), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n615), .A2(new_n620), .A3(new_n618), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT106), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT102), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n625), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n625), .A2(new_n626), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n622), .A2(KEYINPUT106), .A3(new_n624), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n630), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G230gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n333), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n617), .A2(new_n581), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n573), .A2(new_n580), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n612), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n581), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(new_n643), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n647), .B2(new_n639), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G176gat), .ZN(new_n650));
  INV_X1    g449(.A(G204gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n646), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(new_n639), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n601), .A2(new_n637), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n555), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n502), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g460(.A1(new_n659), .A2(new_n445), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT16), .B(G8gat), .Z(new_n663));
  AND2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n665), .B(new_n666), .C1(new_n235), .C2(new_n662), .ZN(G1325gat));
  OAI21_X1  g466(.A(G15gat), .B1(new_n659), .B2(new_n553), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n349), .A2(G15gat), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n659), .B2(new_n669), .ZN(G1326gat));
  NOR2_X1   g469(.A1(new_n659), .A2(new_n418), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT43), .B(G22gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  AOI21_X1  g472(.A(new_n636), .B1(new_n512), .B2(new_n554), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n636), .B(new_n678), .C1(new_n512), .C2(new_n554), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n502), .ZN(new_n682));
  INV_X1    g481(.A(new_n657), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n601), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n257), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n681), .A2(KEYINPUT109), .A3(new_n682), .A4(new_n685), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(G29gat), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n684), .A2(new_n636), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n555), .A2(new_n217), .A3(new_n682), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT107), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT45), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n690), .A2(new_n695), .A3(new_n696), .ZN(G1328gat));
  NAND4_X1  g496(.A1(new_n555), .A2(new_n218), .A3(new_n542), .A4(new_n691), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT46), .Z(new_n699));
  AND3_X1   g498(.A1(new_n681), .A2(new_n542), .A3(new_n685), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(new_n218), .ZN(G1329gat));
  XNOR2_X1  g500(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n553), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n512), .A2(new_n554), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n675), .B1(new_n705), .B2(new_n637), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n704), .B(new_n685), .C1(new_n706), .C2(new_n679), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n707), .A2(G43gat), .ZN(new_n708));
  INV_X1    g507(.A(G43gat), .ZN(new_n709));
  INV_X1    g508(.A(new_n349), .ZN(new_n710));
  AND4_X1   g509(.A1(new_n709), .A2(new_n555), .A3(new_n710), .A4(new_n691), .ZN(new_n711));
  OAI211_X1 g510(.A(KEYINPUT111), .B(new_n703), .C1(new_n708), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n707), .B2(G43gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT47), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n713), .B2(new_n702), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n712), .A2(new_n714), .A3(new_n716), .ZN(G1330gat));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n419), .B(new_n685), .C1(new_n706), .C2(new_n679), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(G50gat), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n418), .A2(G50gat), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n555), .A2(new_n691), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n719), .B2(G50gat), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI221_X4 g524(.A(new_n722), .B1(new_n718), .B2(KEYINPUT48), .C1(new_n719), .C2(G50gat), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n598), .A2(new_n600), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n636), .ZN(new_n729));
  INV_X1    g528(.A(new_n257), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n683), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT113), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n729), .A2(KEYINPUT113), .A3(new_n731), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n705), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n502), .B(KEYINPUT114), .Z(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n564), .ZN(G1332gat));
  AOI211_X1 g536(.A(new_n445), .B(new_n734), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n734), .B2(new_n553), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n742));
  INV_X1    g541(.A(G71gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n710), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n741), .B(new_n742), .C1(new_n734), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n733), .A2(new_n732), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n512), .B2(new_n554), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n743), .B1(new_n747), .B2(new_n704), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n734), .A2(new_n744), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT115), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n747), .A2(new_n419), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n730), .A2(new_n728), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n657), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n681), .A2(new_n682), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT116), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n607), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(KEYINPUT116), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n705), .A2(new_n637), .A3(new_n755), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT51), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n674), .A2(new_n764), .A3(new_n755), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n657), .A3(new_n765), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n502), .A2(new_n607), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n760), .A2(new_n761), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  OR3_X1    g567(.A1(new_n766), .A2(G92gat), .A3(new_n445), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n681), .A2(new_n542), .A3(new_n757), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n756), .B1(new_n676), .B2(new_n680), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n435), .B1(new_n774), .B2(new_n542), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n766), .A2(G92gat), .A3(new_n445), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT52), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(new_n604), .B1(new_n766), .B2(new_n349), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n681), .A2(G99gat), .A3(new_n704), .A4(new_n757), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(KEYINPUT117), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1338gat));
  OAI211_X1 g584(.A(new_n419), .B(new_n757), .C1(new_n706), .C2(new_n679), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n786), .A2(G106gat), .B1(KEYINPUT118), .B2(KEYINPUT53), .ZN(new_n787));
  OR2_X1    g586(.A1(KEYINPUT118), .A2(KEYINPUT53), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n418), .A2(G106gat), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n763), .A2(new_n657), .A3(new_n765), .A4(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n787), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(G1339gat));
  NAND4_X1  g592(.A1(new_n728), .A2(new_n636), .A3(new_n257), .A4(new_n683), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n240), .B1(new_n237), .B2(new_n239), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n243), .A2(new_n244), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n206), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n657), .A2(new_n254), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n644), .A2(new_n645), .A3(new_n639), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n652), .B1(new_n646), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n656), .A3(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n636), .B(new_n798), .C1(new_n257), .C2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n254), .A2(new_n797), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n601), .B1(new_n811), .B2(new_n636), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n794), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n808), .B(new_n601), .C1(new_n636), .C2(new_n811), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(KEYINPUT119), .A3(new_n794), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n542), .A2(new_n502), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n420), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n821), .A2(new_n260), .A3(new_n257), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n818), .A2(new_n735), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n509), .A2(new_n542), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n730), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n822), .B1(new_n827), .B2(new_n260), .ZN(G1340gat));
  NOR3_X1   g627(.A1(new_n821), .A2(new_n261), .A3(new_n683), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n826), .A2(new_n657), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n261), .ZN(G1341gat));
  OAI21_X1  g630(.A(G127gat), .B1(new_n821), .B2(new_n601), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n601), .A2(G127gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n825), .B2(new_n833), .ZN(G1342gat));
  OR2_X1    g633(.A1(new_n636), .A2(G134gat), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n825), .A2(KEYINPUT56), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n821), .B2(new_n636), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT56), .B1(new_n825), .B2(new_n835), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(G1343gat));
  NOR3_X1   g638(.A1(new_n704), .A2(new_n542), .A3(new_n418), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n823), .A2(new_n357), .A3(new_n730), .A4(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n816), .A2(new_n842), .B1(new_n658), .B2(new_n257), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n842), .B2(new_n816), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n418), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n815), .A2(new_n419), .A3(new_n817), .ZN(new_n847));
  XNOR2_X1  g646(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n844), .A2(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n553), .A2(new_n820), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n849), .A2(new_n257), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n841), .B1(new_n851), .B2(new_n357), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n841), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OAI221_X1 g655(.A(new_n841), .B1(new_n854), .B2(new_n853), .C1(new_n851), .C2(new_n357), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1344gat));
  AND2_X1   g657(.A1(new_n823), .A2(new_n840), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n358), .A3(new_n657), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n813), .A2(new_n419), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n845), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n847), .B2(new_n848), .ZN(new_n864));
  INV_X1    g663(.A(new_n850), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n657), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n358), .B1(new_n866), .B2(KEYINPUT123), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n864), .A2(new_n868), .A3(new_n657), .A4(new_n865), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n861), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n849), .A2(new_n683), .A3(new_n850), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(KEYINPUT59), .A3(new_n358), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n860), .B1(new_n870), .B2(new_n872), .ZN(G1345gat));
  NAND3_X1  g672(.A1(new_n859), .A2(new_n374), .A3(new_n728), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n849), .A2(new_n601), .A3(new_n850), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n374), .ZN(G1346gat));
  NAND4_X1  g675(.A1(new_n859), .A2(new_n365), .A3(new_n367), .A4(new_n637), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n849), .A2(new_n636), .A3(new_n850), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n368), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(G1347gat));
  AND2_X1   g681(.A1(new_n735), .A2(new_n542), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n815), .A2(new_n420), .A3(new_n817), .A4(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(G169gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(new_n257), .ZN(new_n886));
  INV_X1    g685(.A(new_n509), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n682), .A2(new_n445), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n815), .A2(new_n887), .A3(new_n817), .A4(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n730), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n886), .B1(new_n891), .B2(new_n885), .ZN(G1348gat));
  OAI21_X1  g691(.A(G176gat), .B1(new_n884), .B2(new_n683), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n683), .A2(G176gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT125), .ZN(G1349gat));
  NAND2_X1  g695(.A1(new_n728), .A2(new_n313), .ZN(new_n897));
  OR3_X1    g696(.A1(new_n889), .A2(KEYINPUT126), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G183gat), .B1(new_n884), .B2(new_n601), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT126), .B1(new_n889), .B2(new_n897), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n902));
  OR2_X1    g701(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1350gat));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n308), .A3(new_n637), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n884), .A2(new_n636), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(G190gat), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n908), .B2(G190gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(G1351gat));
  NOR2_X1   g712(.A1(new_n704), .A2(new_n418), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n819), .A2(new_n914), .A3(new_n888), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916), .B2(new_n730), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n883), .A2(new_n553), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n864), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n730), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  NOR3_X1   g721(.A1(new_n915), .A2(G204gat), .A3(new_n683), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n864), .A2(new_n657), .A3(new_n919), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n925), .B(new_n926), .C1(new_n651), .C2(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n916), .A2(new_n584), .A3(new_n728), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n864), .A2(new_n728), .A3(new_n919), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  AOI21_X1  g732(.A(G218gat), .B1(new_n916), .B2(new_n637), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n637), .A2(G218gat), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n920), .B2(new_n936), .ZN(G1355gat));
endmodule


