

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781;

  XNOR2_X1 U366 ( .A(n347), .B(n346), .ZN(n378) );
  INV_X1 U367 ( .A(n379), .ZN(n346) );
  NOR2_X4 U368 ( .A1(n719), .A2(n567), .ZN(n568) );
  XNOR2_X2 U369 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X2 U370 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U371 ( .A1(n747), .A2(G472), .ZN(n347) );
  AND2_X2 U372 ( .A1(n747), .A2(G475), .ZN(n674) );
  NAND2_X2 U373 ( .A1(n530), .A2(G214), .ZN(n716) );
  XNOR2_X2 U374 ( .A(G902), .B(KEYINPUT15), .ZN(n594) );
  AND2_X2 U375 ( .A1(n348), .A2(n458), .ZN(n359) );
  NAND2_X1 U376 ( .A1(n670), .A2(n468), .ZN(n348) );
  AND2_X1 U377 ( .A1(n477), .A2(n478), .ZN(n349) );
  NOR2_X2 U378 ( .A1(n682), .A2(n755), .ZN(n683) );
  NOR2_X2 U379 ( .A1(n657), .A2(n755), .ZN(n659) );
  XNOR2_X2 U380 ( .A(n356), .B(KEYINPUT45), .ZN(n644) );
  NAND2_X2 U381 ( .A1(n357), .A2(n593), .ZN(n356) );
  NAND2_X1 U382 ( .A1(n457), .A2(n455), .ZN(n358) );
  NOR2_X1 U383 ( .A1(n592), .A2(n665), .ZN(n593) );
  XNOR2_X1 U384 ( .A(n614), .B(KEYINPUT42), .ZN(n780) );
  XNOR2_X1 U385 ( .A(n607), .B(KEYINPUT40), .ZN(n453) );
  NAND2_X1 U386 ( .A1(n485), .A2(n484), .ZN(n483) );
  XNOR2_X1 U387 ( .A(n620), .B(n605), .ZN(n717) );
  INV_X1 U388 ( .A(n624), .ZN(n350) );
  AND2_X1 U389 ( .A1(n440), .A2(n439), .ZN(n419) );
  XNOR2_X2 U390 ( .A(n521), .B(n520), .ZN(n764) );
  XNOR2_X2 U391 ( .A(n352), .B(n351), .ZN(n521) );
  XNOR2_X2 U392 ( .A(n354), .B(G113), .ZN(n351) );
  XNOR2_X2 U393 ( .A(n353), .B(n355), .ZN(n352) );
  XNOR2_X2 U394 ( .A(G119), .B(G116), .ZN(n353) );
  XNOR2_X2 U395 ( .A(G101), .B(KEYINPUT3), .ZN(n354) );
  XNOR2_X2 U396 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n355) );
  NAND2_X1 U397 ( .A1(n359), .A2(n358), .ZN(n357) );
  INV_X1 U398 ( .A(n360), .ZN(n591) );
  NAND2_X1 U399 ( .A1(n575), .A2(n360), .ZN(n576) );
  XNOR2_X2 U400 ( .A(n570), .B(n569), .ZN(n360) );
  NAND2_X1 U401 ( .A1(n360), .A2(n578), .ZN(n663) );
  XNOR2_X1 U402 ( .A(n398), .B(n374), .ZN(n397) );
  NAND2_X1 U403 ( .A1(n453), .A2(n780), .ZN(n398) );
  NAND2_X1 U404 ( .A1(n407), .A2(n406), .ZN(n408) );
  BUF_X1 U405 ( .A(n764), .Z(n361) );
  NAND2_X1 U406 ( .A1(n465), .A2(n462), .ZN(n362) );
  NAND2_X1 U407 ( .A1(n465), .A2(n462), .ZN(n670) );
  INV_X1 U408 ( .A(n716), .ZN(n427) );
  NAND2_X1 U409 ( .A1(n442), .A2(n366), .ZN(n400) );
  XNOR2_X1 U410 ( .A(n504), .B(KEYINPUT68), .ZN(n706) );
  NOR2_X1 U411 ( .A1(n699), .A2(n567), .ZN(n504) );
  NAND2_X1 U412 ( .A1(n699), .A2(n609), .ZN(n617) );
  AND2_X1 U413 ( .A1(n706), .A2(n624), .ZN(n601) );
  INV_X1 U414 ( .A(KEYINPUT44), .ZN(n468) );
  XNOR2_X1 U415 ( .A(n396), .B(KEYINPUT48), .ZN(n482) );
  XNOR2_X1 U416 ( .A(n400), .B(n630), .ZN(n399) );
  XNOR2_X1 U417 ( .A(n425), .B(n424), .ZN(n560) );
  INV_X1 U418 ( .A(KEYINPUT8), .ZN(n424) );
  NAND2_X1 U419 ( .A1(n508), .A2(G234), .ZN(n425) );
  XNOR2_X1 U420 ( .A(G122), .B(KEYINPUT99), .ZN(n553) );
  XNOR2_X1 U421 ( .A(G116), .B(G107), .ZN(n556) );
  XNOR2_X1 U422 ( .A(G113), .B(G122), .ZN(n540) );
  XNOR2_X1 U423 ( .A(G143), .B(G104), .ZN(n543) );
  XNOR2_X1 U424 ( .A(G146), .B(G125), .ZN(n524) );
  XNOR2_X1 U425 ( .A(n470), .B(n469), .ZN(n526) );
  XNOR2_X1 U426 ( .A(KEYINPUT88), .B(KEYINPUT18), .ZN(n469) );
  XNOR2_X1 U427 ( .A(n471), .B(KEYINPUT17), .ZN(n470) );
  XNOR2_X1 U428 ( .A(KEYINPUT82), .B(KEYINPUT90), .ZN(n471) );
  XNOR2_X1 U429 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n505) );
  NAND2_X1 U430 ( .A1(n421), .A2(n420), .ZN(n571) );
  XNOR2_X1 U431 ( .A(KEYINPUT16), .B(G122), .ZN(n520) );
  XNOR2_X1 U432 ( .A(n524), .B(n426), .ZN(n770) );
  XNOR2_X1 U433 ( .A(G140), .B(KEYINPUT10), .ZN(n426) );
  XNOR2_X1 U434 ( .A(n472), .B(n512), .ZN(n654) );
  XNOR2_X1 U435 ( .A(G101), .B(G140), .ZN(n510) );
  XNOR2_X1 U436 ( .A(n613), .B(n410), .ZN(n734) );
  XNOR2_X1 U437 ( .A(n612), .B(KEYINPUT110), .ZN(n410) );
  NOR2_X1 U438 ( .A1(n720), .A2(n719), .ZN(n613) );
  XNOR2_X1 U439 ( .A(n408), .B(n606), .ZN(n632) );
  AND2_X1 U440 ( .A1(n454), .A2(n717), .ZN(n407) );
  NAND2_X1 U441 ( .A1(n449), .A2(n450), .ZN(n392) );
  INV_X1 U442 ( .A(n617), .ZN(n431) );
  OR2_X1 U443 ( .A1(n752), .A2(G902), .ZN(n404) );
  NAND2_X1 U444 ( .A1(KEYINPUT1), .A2(n418), .ZN(n417) );
  INV_X1 U445 ( .A(n436), .ZN(n418) );
  NOR2_X1 U446 ( .A1(n461), .A2(n468), .ZN(n456) );
  INV_X1 U447 ( .A(G237), .ZN(n528) );
  NAND2_X1 U448 ( .A1(n438), .A2(n437), .ZN(n436) );
  INV_X1 U449 ( .A(G469), .ZN(n438) );
  NAND2_X1 U450 ( .A1(n414), .A2(n412), .ZN(n411) );
  NAND2_X1 U451 ( .A1(KEYINPUT1), .A2(n413), .ZN(n412) );
  OR2_X1 U452 ( .A1(n654), .A2(n417), .ZN(n414) );
  INV_X1 U453 ( .A(n439), .ZN(n413) );
  NOR2_X1 U454 ( .A1(n440), .A2(n416), .ZN(n415) );
  XNOR2_X1 U455 ( .A(n548), .B(n506), .ZN(n428) );
  XNOR2_X1 U456 ( .A(G137), .B(G134), .ZN(n506) );
  NAND2_X1 U457 ( .A1(G234), .A2(G237), .ZN(n533) );
  NAND2_X1 U458 ( .A1(n539), .A2(n371), .ZN(n487) );
  AND2_X1 U459 ( .A1(n571), .A2(n706), .ZN(n517) );
  NAND2_X1 U460 ( .A1(G902), .A2(G469), .ZN(n439) );
  XNOR2_X1 U461 ( .A(n448), .B(n447), .ZN(n566) );
  INV_X1 U462 ( .A(G478), .ZN(n447) );
  OR2_X1 U463 ( .A1(n749), .A2(G902), .ZN(n448) );
  INV_X1 U464 ( .A(n641), .ZN(n480) );
  XNOR2_X1 U465 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U466 ( .A(n556), .B(n555), .ZN(n557) );
  INV_X1 U467 ( .A(KEYINPUT98), .ZN(n555) );
  NOR2_X1 U468 ( .A1(G953), .A2(G237), .ZN(n547) );
  INV_X1 U469 ( .A(KEYINPUT11), .ZN(n542) );
  XNOR2_X1 U470 ( .A(n384), .B(n383), .ZN(n677) );
  XNOR2_X1 U471 ( .A(n764), .B(n527), .ZN(n384) );
  NAND2_X1 U472 ( .A1(n450), .A2(n367), .ZN(n633) );
  XNOR2_X1 U473 ( .A(n601), .B(n600), .ZN(n406) );
  XNOR2_X1 U474 ( .A(n552), .B(G475), .ZN(n445) );
  OR2_X1 U475 ( .A1(n672), .A2(G902), .ZN(n446) );
  INV_X1 U476 ( .A(n566), .ZN(n584) );
  NAND2_X1 U477 ( .A1(n601), .A2(n433), .ZN(n580) );
  AND2_X1 U478 ( .A1(n566), .A2(n444), .ZN(n616) );
  XNOR2_X1 U479 ( .A(n405), .B(n495), .ZN(n752) );
  XNOR2_X1 U480 ( .A(n423), .B(n770), .ZN(n405) );
  XOR2_X1 U481 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n493) );
  INV_X2 U482 ( .A(G953), .ZN(n508) );
  NAND2_X1 U483 ( .A1(n734), .A2(n452), .ZN(n614) );
  NOR2_X1 U484 ( .A1(n627), .A2(n350), .ZN(n452) );
  XNOR2_X1 U485 ( .A(n389), .B(KEYINPUT112), .ZN(n442) );
  AND2_X1 U486 ( .A1(n422), .A2(n370), .ZN(n363) );
  INV_X1 U487 ( .A(n699), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n446), .B(n445), .ZN(n585) );
  INV_X1 U489 ( .A(n585), .ZN(n444) );
  NOR2_X1 U490 ( .A1(n617), .A2(n427), .ZN(n489) );
  NAND2_X1 U491 ( .A1(n641), .A2(n481), .ZN(n364) );
  OR2_X1 U492 ( .A1(n451), .A2(n636), .ZN(n365) );
  AND2_X1 U493 ( .A1(n664), .A2(n629), .ZN(n366) );
  AND2_X1 U494 ( .A1(n618), .A2(n489), .ZN(n367) );
  AND2_X1 U495 ( .A1(n381), .A2(n479), .ZN(n368) );
  AND2_X1 U496 ( .A1(n517), .A2(n376), .ZN(n369) );
  AND2_X1 U497 ( .A1(n416), .A2(n439), .ZN(n370) );
  INV_X1 U498 ( .A(G902), .ZN(n437) );
  INV_X1 U499 ( .A(n660), .ZN(n618) );
  XNOR2_X1 U500 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n371) );
  XNOR2_X1 U501 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n372) );
  XOR2_X1 U502 ( .A(KEYINPUT101), .B(KEYINPUT6), .Z(n373) );
  INV_X1 U503 ( .A(KEYINPUT34), .ZN(n479) );
  XOR2_X1 U504 ( .A(n615), .B(KEYINPUT64), .Z(n374) );
  NAND2_X1 U505 ( .A1(n642), .A2(n595), .ZN(n375) );
  INV_X1 U506 ( .A(KEYINPUT84), .ZN(n595) );
  XNOR2_X2 U507 ( .A(n385), .B(KEYINPUT65), .ZN(n747) );
  INV_X1 U508 ( .A(n433), .ZN(n376) );
  XNOR2_X1 U509 ( .A(n377), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U510 ( .A1(n378), .A2(n651), .ZN(n377) );
  INV_X1 U511 ( .A(n648), .ZN(n379) );
  OR2_X1 U512 ( .A1(n654), .A2(n436), .ZN(n422) );
  XNOR2_X2 U513 ( .A(n380), .B(n645), .ZN(n702) );
  NOR2_X1 U514 ( .A1(n647), .A2(G902), .ZN(n380) );
  BUF_X2 U515 ( .A(n571), .Z(n705) );
  NOR2_X1 U516 ( .A1(n415), .A2(n411), .ZN(n421) );
  XNOR2_X1 U517 ( .A(n519), .B(n518), .ZN(n733) );
  NAND2_X1 U518 ( .A1(n486), .A2(n483), .ZN(n381) );
  NAND2_X1 U519 ( .A1(n486), .A2(n483), .ZN(n434) );
  BUF_X1 U520 ( .A(n747), .Z(n751) );
  NAND2_X1 U521 ( .A1(n434), .A2(n568), .ZN(n570) );
  NOR2_X1 U522 ( .A1(n364), .A2(n482), .ZN(n394) );
  BUF_X1 U523 ( .A(n644), .Z(n756) );
  XNOR2_X2 U524 ( .A(n382), .B(n529), .ZN(n619) );
  NAND2_X1 U525 ( .A1(n677), .A2(n594), .ZN(n382) );
  XNOR2_X1 U526 ( .A(n435), .B(n522), .ZN(n383) );
  NAND2_X1 U527 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U528 ( .A(n740), .ZN(n386) );
  XNOR2_X1 U529 ( .A(n388), .B(KEYINPUT66), .ZN(n387) );
  NAND2_X1 U530 ( .A1(n393), .A2(n643), .ZN(n388) );
  NOR2_X2 U531 ( .A1(n409), .A2(n737), .ZN(n740) );
  NAND2_X1 U532 ( .A1(n390), .A2(n705), .ZN(n389) );
  XNOR2_X1 U533 ( .A(n392), .B(n391), .ZN(n390) );
  INV_X1 U534 ( .A(KEYINPUT36), .ZN(n391) );
  NAND2_X1 U535 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U536 ( .A1(n402), .A2(n401), .ZN(n395) );
  NAND2_X1 U537 ( .A1(n399), .A2(n397), .ZN(n396) );
  NAND2_X1 U538 ( .A1(n644), .A2(n375), .ZN(n401) );
  NAND2_X1 U539 ( .A1(n403), .A2(n595), .ZN(n402) );
  INV_X1 U540 ( .A(n644), .ZN(n403) );
  XNOR2_X2 U541 ( .A(n404), .B(n500), .ZN(n699) );
  AND2_X1 U542 ( .A1(n454), .A2(n406), .ZN(n623) );
  NAND2_X1 U543 ( .A1(n771), .A2(KEYINPUT2), .ZN(n409) );
  INV_X1 U544 ( .A(n621), .ZN(n478) );
  INV_X1 U545 ( .A(n663), .ZN(n461) );
  NAND2_X1 U546 ( .A1(n464), .A2(n463), .ZN(n462) );
  NAND2_X2 U547 ( .A1(n619), .A2(n716), .ZN(n532) );
  NAND2_X1 U548 ( .A1(n581), .A2(KEYINPUT34), .ZN(n477) );
  INV_X1 U549 ( .A(KEYINPUT1), .ZN(n416) );
  NAND2_X1 U550 ( .A1(n363), .A2(n440), .ZN(n420) );
  NAND2_X1 U551 ( .A1(n419), .A2(n422), .ZN(n624) );
  INV_X1 U552 ( .A(n442), .ZN(n443) );
  NAND2_X1 U553 ( .A1(n560), .A2(G221), .ZN(n423) );
  XNOR2_X2 U554 ( .A(n435), .B(n428), .ZN(n769) );
  XNOR2_X2 U555 ( .A(n429), .B(G131), .ZN(n548) );
  XNOR2_X2 U556 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n429) );
  XNOR2_X2 U557 ( .A(n563), .B(n505), .ZN(n435) );
  XNOR2_X2 U558 ( .A(n430), .B(G128), .ZN(n563) );
  XNOR2_X2 U559 ( .A(G143), .B(KEYINPUT83), .ZN(n430) );
  AND2_X1 U560 ( .A1(n702), .A2(n431), .ZN(n611) );
  OR2_X1 U561 ( .A1(n702), .A2(n432), .ZN(n577) );
  XNOR2_X1 U562 ( .A(n702), .B(n373), .ZN(n588) );
  INV_X1 U563 ( .A(n702), .ZN(n433) );
  INV_X1 U564 ( .A(n381), .ZN(n581) );
  NAND2_X1 U565 ( .A1(n369), .A2(n381), .ZN(n579) );
  NAND2_X1 U566 ( .A1(n654), .A2(G469), .ZN(n440) );
  BUF_X1 U567 ( .A(n733), .Z(n441) );
  XNOR2_X1 U568 ( .A(n443), .B(n666), .ZN(G27) );
  NOR2_X1 U569 ( .A1(n660), .A2(n365), .ZN(n449) );
  INV_X1 U570 ( .A(n588), .ZN(n450) );
  INV_X1 U571 ( .A(n489), .ZN(n451) );
  INV_X1 U572 ( .A(n734), .ZN(n714) );
  XNOR2_X1 U573 ( .A(n453), .B(G131), .ZN(G33) );
  AND2_X1 U574 ( .A1(n604), .A2(n608), .ZN(n454) );
  NAND2_X1 U575 ( .A1(n668), .A2(n663), .ZN(n459) );
  XNOR2_X2 U576 ( .A(n576), .B(KEYINPUT32), .ZN(n668) );
  AND2_X1 U577 ( .A1(n668), .A2(n456), .ZN(n455) );
  INV_X1 U578 ( .A(n362), .ZN(n457) );
  NAND2_X1 U579 ( .A1(n459), .A2(n468), .ZN(n458) );
  INV_X1 U580 ( .A(n474), .ZN(n463) );
  NOR2_X1 U581 ( .A1(n473), .A2(n372), .ZN(n464) );
  AND2_X2 U582 ( .A1(n467), .A2(n466), .ZN(n465) );
  NAND2_X1 U583 ( .A1(n473), .A2(n372), .ZN(n466) );
  NAND2_X1 U584 ( .A1(n474), .A2(n372), .ZN(n467) );
  AND2_X2 U585 ( .A1(n488), .A2(n487), .ZN(n486) );
  XNOR2_X1 U586 ( .A(n472), .B(n490), .ZN(n647) );
  XNOR2_X2 U587 ( .A(n769), .B(G146), .ZN(n472) );
  AND2_X1 U588 ( .A1(n733), .A2(n368), .ZN(n473) );
  NAND2_X1 U589 ( .A1(n475), .A2(n349), .ZN(n474) );
  NAND2_X1 U590 ( .A1(n476), .A2(KEYINPUT34), .ZN(n475) );
  INV_X1 U591 ( .A(n733), .ZN(n476) );
  NOR2_X2 U592 ( .A1(n482), .A2(n480), .ZN(n771) );
  NAND2_X1 U593 ( .A1(n594), .A2(KEYINPUT84), .ZN(n481) );
  NOR2_X1 U594 ( .A1(n539), .A2(n371), .ZN(n484) );
  INV_X1 U595 ( .A(n625), .ZN(n485) );
  NAND2_X1 U596 ( .A1(n625), .A2(n371), .ZN(n488) );
  XNOR2_X2 U597 ( .A(n532), .B(n531), .ZN(n625) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U599 ( .A(n521), .B(n516), .Z(n490) );
  XNOR2_X1 U600 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U601 ( .A(n545), .B(n544), .ZN(n546) );
  INV_X1 U602 ( .A(KEYINPUT107), .ZN(n600) );
  BUF_X1 U603 ( .A(n677), .Z(n679) );
  INV_X1 U604 ( .A(n755), .ZN(n651) );
  INV_X1 U605 ( .A(KEYINPUT121), .ZN(n658) );
  XOR2_X1 U606 ( .A(G110), .B(G128), .Z(n492) );
  XNOR2_X1 U607 ( .A(G119), .B(G137), .ZN(n491) );
  XNOR2_X1 U608 ( .A(n492), .B(n491), .ZN(n494) );
  XOR2_X1 U609 ( .A(KEYINPUT81), .B(KEYINPUT25), .Z(n499) );
  XOR2_X1 U610 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n497) );
  NAND2_X1 U611 ( .A1(G234), .A2(n594), .ZN(n496) );
  XNOR2_X1 U612 ( .A(n497), .B(n496), .ZN(n501) );
  NAND2_X1 U613 ( .A1(G217), .A2(n501), .ZN(n498) );
  XNOR2_X1 U614 ( .A(n499), .B(n498), .ZN(n500) );
  AND2_X1 U615 ( .A1(n501), .A2(G221), .ZN(n503) );
  XNOR2_X1 U616 ( .A(KEYINPUT94), .B(KEYINPUT21), .ZN(n502) );
  XNOR2_X1 U617 ( .A(n503), .B(n502), .ZN(n700) );
  INV_X1 U618 ( .A(n700), .ZN(n567) );
  XOR2_X1 U619 ( .A(G104), .B(G110), .Z(n507) );
  XNOR2_X1 U620 ( .A(n507), .B(G107), .ZN(n762) );
  XNOR2_X1 U621 ( .A(n762), .B(KEYINPUT75), .ZN(n522) );
  NAND2_X1 U622 ( .A1(n508), .A2(G227), .ZN(n509) );
  XNOR2_X1 U623 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U624 ( .A(n522), .B(n511), .ZN(n512) );
  NAND2_X1 U625 ( .A1(n547), .A2(G210), .ZN(n513) );
  XNOR2_X1 U626 ( .A(n513), .B(KEYINPUT5), .ZN(n515) );
  XNOR2_X1 U627 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n514) );
  XNOR2_X1 U628 ( .A(n515), .B(n514), .ZN(n516) );
  INV_X1 U629 ( .A(G472), .ZN(n645) );
  INV_X1 U630 ( .A(n588), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n573), .A2(n517), .ZN(n519) );
  XNOR2_X1 U632 ( .A(KEYINPUT76), .B(KEYINPUT33), .ZN(n518) );
  NAND2_X1 U633 ( .A1(G224), .A2(n508), .ZN(n523) );
  XNOR2_X1 U634 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U635 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U636 ( .A1(n437), .A2(n528), .ZN(n530) );
  AND2_X1 U637 ( .A1(n530), .A2(G210), .ZN(n529) );
  INV_X1 U638 ( .A(KEYINPUT19), .ZN(n531) );
  XNOR2_X1 U639 ( .A(n533), .B(KEYINPUT14), .ZN(n537) );
  NAND2_X1 U640 ( .A1(G902), .A2(n537), .ZN(n534) );
  XNOR2_X1 U641 ( .A(KEYINPUT91), .B(n534), .ZN(n535) );
  NAND2_X1 U642 ( .A1(n535), .A2(G953), .ZN(n596) );
  NOR2_X1 U643 ( .A1(G898), .A2(n596), .ZN(n536) );
  XNOR2_X1 U644 ( .A(n536), .B(KEYINPUT92), .ZN(n538) );
  NAND2_X1 U645 ( .A1(G952), .A2(n537), .ZN(n731) );
  NOR2_X1 U646 ( .A1(n731), .A2(G953), .ZN(n598) );
  NOR2_X1 U647 ( .A1(n538), .A2(n598), .ZN(n539) );
  XNOR2_X1 U648 ( .A(KEYINPUT13), .B(KEYINPUT96), .ZN(n552) );
  XOR2_X1 U649 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n541) );
  XNOR2_X1 U650 ( .A(n541), .B(n540), .ZN(n545) );
  XNOR2_X1 U651 ( .A(n546), .B(n770), .ZN(n551) );
  NAND2_X1 U652 ( .A1(n547), .A2(G214), .ZN(n549) );
  XOR2_X1 U653 ( .A(n549), .B(n548), .Z(n550) );
  XNOR2_X1 U654 ( .A(n551), .B(n550), .ZN(n672) );
  XOR2_X1 U655 ( .A(KEYINPUT7), .B(KEYINPUT97), .Z(n554) );
  XNOR2_X1 U656 ( .A(n554), .B(n553), .ZN(n558) );
  XOR2_X1 U657 ( .A(n559), .B(KEYINPUT9), .Z(n565) );
  NAND2_X1 U658 ( .A1(n560), .A2(G217), .ZN(n561) );
  XNOR2_X1 U659 ( .A(n561), .B(G134), .ZN(n562) );
  XNOR2_X1 U660 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U661 ( .A(n565), .B(n564), .ZN(n749) );
  NAND2_X1 U662 ( .A1(n444), .A2(n584), .ZN(n621) );
  NAND2_X1 U663 ( .A1(n585), .A2(n566), .ZN(n719) );
  XOR2_X1 U664 ( .A(KEYINPUT78), .B(KEYINPUT22), .Z(n569) );
  NAND2_X1 U665 ( .A1(n705), .A2(n699), .ZN(n572) );
  XNOR2_X1 U666 ( .A(n572), .B(KEYINPUT102), .ZN(n574) );
  NOR2_X1 U667 ( .A1(n574), .A2(n450), .ZN(n575) );
  NOR2_X1 U668 ( .A1(n705), .A2(n577), .ZN(n578) );
  XOR2_X1 U669 ( .A(KEYINPUT31), .B(n579), .Z(n695) );
  INV_X1 U670 ( .A(n695), .ZN(n582) );
  NOR2_X1 U671 ( .A1(n581), .A2(n580), .ZN(n684) );
  NOR2_X1 U672 ( .A1(n582), .A2(n684), .ZN(n587) );
  NAND2_X1 U673 ( .A1(n585), .A2(n584), .ZN(n583) );
  XNOR2_X1 U674 ( .A(n583), .B(KEYINPUT100), .ZN(n696) );
  INV_X1 U675 ( .A(n616), .ZN(n586) );
  AND2_X1 U676 ( .A1(n696), .A2(n586), .ZN(n721) );
  NOR2_X1 U677 ( .A1(n587), .A2(n721), .ZN(n592) );
  NOR2_X1 U678 ( .A1(n705), .A2(n699), .ZN(n589) );
  NAND2_X1 U679 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U680 ( .A1(n591), .A2(n590), .ZN(n665) );
  INV_X1 U681 ( .A(n594), .ZN(n642) );
  XNOR2_X1 U682 ( .A(KEYINPUT104), .B(n596), .ZN(n597) );
  NOR2_X1 U683 ( .A1(G900), .A2(n597), .ZN(n599) );
  OR2_X1 U684 ( .A1(n599), .A2(n598), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n702), .A2(n716), .ZN(n603) );
  XOR2_X1 U686 ( .A(KEYINPUT108), .B(KEYINPUT30), .Z(n602) );
  XNOR2_X1 U687 ( .A(n603), .B(n602), .ZN(n604) );
  INV_X1 U688 ( .A(KEYINPUT38), .ZN(n605) );
  XOR2_X1 U689 ( .A(KEYINPUT77), .B(KEYINPUT39), .Z(n606) );
  NAND2_X1 U690 ( .A1(n632), .A2(n616), .ZN(n607) );
  AND2_X1 U691 ( .A1(n700), .A2(n608), .ZN(n609) );
  XNOR2_X1 U692 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n610) );
  XNOR2_X1 U693 ( .A(n611), .B(n610), .ZN(n627) );
  NAND2_X1 U694 ( .A1(n717), .A2(n716), .ZN(n720) );
  XNOR2_X1 U695 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n612) );
  XOR2_X1 U696 ( .A(KEYINPUT46), .B(KEYINPUT87), .Z(n615) );
  XNOR2_X1 U697 ( .A(n616), .B(KEYINPUT103), .ZN(n660) );
  BUF_X1 U698 ( .A(n619), .Z(n620) );
  INV_X1 U699 ( .A(n620), .ZN(n636) );
  NOR2_X1 U700 ( .A1(n621), .A2(n636), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n664) );
  OR2_X1 U702 ( .A1(n625), .A2(n350), .ZN(n626) );
  OR2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n690) );
  NOR2_X1 U704 ( .A1(n721), .A2(n690), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n628), .B(KEYINPUT47), .ZN(n629) );
  INV_X1 U706 ( .A(KEYINPUT72), .ZN(n630) );
  INV_X1 U707 ( .A(n696), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n698) );
  NOR2_X1 U709 ( .A1(n633), .A2(n705), .ZN(n635) );
  XNOR2_X1 U710 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n635), .B(n634), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n639) );
  INV_X1 U713 ( .A(KEYINPUT106), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n639), .B(n638), .ZN(n779) );
  INV_X1 U715 ( .A(n779), .ZN(n640) );
  AND2_X1 U716 ( .A1(n698), .A2(n640), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(KEYINPUT2), .ZN(n643) );
  INV_X1 U718 ( .A(n756), .ZN(n737) );
  XNOR2_X1 U719 ( .A(KEYINPUT113), .B(KEYINPUT62), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n648) );
  INV_X1 U721 ( .A(G952), .ZN(n650) );
  AND2_X1 U722 ( .A1(n650), .A2(G953), .ZN(n755) );
  NAND2_X1 U723 ( .A1(n747), .A2(G469), .ZN(n656) );
  XOR2_X1 U724 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n652) );
  XNOR2_X1 U725 ( .A(n652), .B(KEYINPUT58), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(G54) );
  NOR2_X1 U728 ( .A1(n660), .A2(n690), .ZN(n662) );
  XNOR2_X1 U729 ( .A(G146), .B(KEYINPUT115), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n662), .B(n661), .ZN(G48) );
  XNOR2_X1 U731 ( .A(n663), .B(G110), .ZN(G12) );
  XNOR2_X1 U732 ( .A(n664), .B(G143), .ZN(G45) );
  XOR2_X1 U733 ( .A(G101), .B(n665), .Z(G3) );
  XNOR2_X1 U734 ( .A(G125), .B(KEYINPUT37), .ZN(n666) );
  XNOR2_X1 U735 ( .A(G119), .B(KEYINPUT126), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(G21) );
  XNOR2_X1 U737 ( .A(G122), .B(KEYINPUT125), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n362), .B(n669), .ZN(G24) );
  XOR2_X1 U739 ( .A(KEYINPUT89), .B(KEYINPUT59), .Z(n671) );
  XNOR2_X1 U740 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U741 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U742 ( .A1(n675), .A2(n755), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n676), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U744 ( .A1(n747), .A2(G210), .ZN(n681) );
  XNOR2_X1 U745 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U747 ( .A(n683), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U748 ( .A(n684), .ZN(n686) );
  NOR2_X1 U749 ( .A1(n686), .A2(n660), .ZN(n685) );
  XOR2_X1 U750 ( .A(G104), .B(n685), .Z(G6) );
  NOR2_X1 U751 ( .A1(n686), .A2(n696), .ZN(n688) );
  XNOR2_X1 U752 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n687) );
  XNOR2_X1 U753 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U754 ( .A(G107), .B(n689), .ZN(G9) );
  NOR2_X1 U755 ( .A1(n690), .A2(n696), .ZN(n692) );
  XNOR2_X1 U756 ( .A(KEYINPUT114), .B(KEYINPUT29), .ZN(n691) );
  XNOR2_X1 U757 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U758 ( .A(G128), .B(n693), .ZN(G30) );
  NOR2_X1 U759 ( .A1(n660), .A2(n695), .ZN(n694) );
  XOR2_X1 U760 ( .A(G113), .B(n694), .Z(G15) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U762 ( .A(G116), .B(n697), .Z(G18) );
  XNOR2_X1 U763 ( .A(G134), .B(n698), .ZN(G36) );
  NOR2_X1 U764 ( .A1(n700), .A2(n432), .ZN(n701) );
  XOR2_X1 U765 ( .A(KEYINPUT49), .B(n701), .Z(n703) );
  NOR2_X1 U766 ( .A1(n703), .A2(n376), .ZN(n704) );
  XOR2_X1 U767 ( .A(n704), .B(KEYINPUT116), .Z(n709) );
  NOR2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U769 ( .A(n707), .B(KEYINPUT50), .ZN(n708) );
  NOR2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U771 ( .A(n710), .B(KEYINPUT117), .ZN(n712) );
  INV_X1 U772 ( .A(n369), .ZN(n711) );
  NAND2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U774 ( .A(KEYINPUT51), .B(n713), .ZN(n715) );
  NOR2_X1 U775 ( .A1(n715), .A2(n714), .ZN(n728) );
  NOR2_X1 U776 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U777 ( .A1(n719), .A2(n718), .ZN(n724) );
  NOR2_X1 U778 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U779 ( .A(n722), .B(KEYINPUT118), .ZN(n723) );
  NOR2_X1 U780 ( .A1(n724), .A2(n723), .ZN(n726) );
  INV_X1 U781 ( .A(n441), .ZN(n725) );
  NOR2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U783 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U784 ( .A(n729), .B(KEYINPUT52), .ZN(n730) );
  NOR2_X1 U785 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U786 ( .A(n732), .B(KEYINPUT119), .ZN(n736) );
  NAND2_X1 U787 ( .A1(n734), .A2(n441), .ZN(n735) );
  NAND2_X1 U788 ( .A1(n736), .A2(n735), .ZN(n744) );
  INV_X1 U789 ( .A(n771), .ZN(n738) );
  NOR2_X1 U790 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U791 ( .A1(n739), .A2(KEYINPUT2), .ZN(n741) );
  NOR2_X1 U792 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U793 ( .A(KEYINPUT85), .B(n742), .Z(n743) );
  NOR2_X1 U794 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U795 ( .A1(n508), .A2(n745), .ZN(n746) );
  XOR2_X1 U796 ( .A(KEYINPUT53), .B(n746), .Z(G75) );
  NAND2_X1 U797 ( .A1(n751), .A2(G478), .ZN(n748) );
  XNOR2_X1 U798 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U799 ( .A1(n755), .A2(n750), .ZN(G63) );
  NAND2_X1 U800 ( .A1(n751), .A2(G217), .ZN(n753) );
  XNOR2_X1 U801 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U802 ( .A1(n755), .A2(n754), .ZN(G66) );
  NAND2_X1 U803 ( .A1(n756), .A2(n508), .ZN(n761) );
  NAND2_X1 U804 ( .A1(G224), .A2(G953), .ZN(n757) );
  XNOR2_X1 U805 ( .A(n757), .B(KEYINPUT122), .ZN(n758) );
  XNOR2_X1 U806 ( .A(KEYINPUT61), .B(n758), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n759), .A2(G898), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(n768) );
  XOR2_X1 U809 ( .A(n762), .B(KEYINPUT123), .Z(n763) );
  XNOR2_X1 U810 ( .A(n361), .B(n763), .ZN(n766) );
  NOR2_X1 U811 ( .A1(G898), .A2(n508), .ZN(n765) );
  NOR2_X1 U812 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U813 ( .A(n768), .B(n767), .ZN(G69) );
  XOR2_X1 U814 ( .A(n769), .B(n770), .Z(n773) );
  XNOR2_X1 U815 ( .A(n771), .B(n773), .ZN(n772) );
  NAND2_X1 U816 ( .A1(n772), .A2(n508), .ZN(n778) );
  XOR2_X1 U817 ( .A(G227), .B(n773), .Z(n774) );
  XNOR2_X1 U818 ( .A(n774), .B(KEYINPUT124), .ZN(n775) );
  NAND2_X1 U819 ( .A1(n775), .A2(G900), .ZN(n776) );
  NAND2_X1 U820 ( .A1(G953), .A2(n776), .ZN(n777) );
  NAND2_X1 U821 ( .A1(n778), .A2(n777), .ZN(G72) );
  XOR2_X1 U822 ( .A(G140), .B(n779), .Z(G42) );
  XOR2_X1 U823 ( .A(G137), .B(n780), .Z(n781) );
  XNOR2_X1 U824 ( .A(KEYINPUT127), .B(n781), .ZN(G39) );
endmodule

