

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593;

  XOR2_X2 U322 ( .A(n331), .B(n319), .Z(n373) );
  XNOR2_X1 U323 ( .A(n400), .B(n399), .ZN(n405) );
  XNOR2_X1 U324 ( .A(KEYINPUT95), .B(n483), .ZN(n575) );
  XOR2_X1 U325 ( .A(n336), .B(n301), .Z(n290) );
  XOR2_X1 U326 ( .A(G92GAT), .B(G64GAT), .Z(n387) );
  INV_X1 U327 ( .A(KEYINPUT102), .ZN(n481) );
  INV_X1 U328 ( .A(KEYINPUT98), .ZN(n397) );
  OR2_X1 U329 ( .A1(n576), .A2(n447), .ZN(n449) );
  NOR2_X1 U330 ( .A1(n382), .A2(n381), .ZN(n383) );
  XNOR2_X1 U331 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U332 ( .A(n492), .B(KEYINPUT105), .ZN(n493) );
  XNOR2_X1 U333 ( .A(n494), .B(n493), .ZN(n530) );
  XNOR2_X1 U334 ( .A(n463), .B(KEYINPUT121), .ZN(n572) );
  XOR2_X1 U335 ( .A(n461), .B(n460), .Z(n540) );
  XNOR2_X1 U336 ( .A(n496), .B(n495), .ZN(n516) );
  XNOR2_X1 U337 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U338 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U339 ( .A(n467), .B(n466), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  INV_X1 U341 ( .A(KEYINPUT54), .ZN(n407) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(KEYINPUT68), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n291), .B(G29GAT), .ZN(n292) );
  XOR2_X1 U344 ( .A(n292), .B(KEYINPUT7), .Z(n294) );
  XNOR2_X1 U345 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n293) );
  XOR2_X1 U346 ( .A(n294), .B(n293), .Z(n331) );
  XOR2_X1 U347 ( .A(G85GAT), .B(KEYINPUT73), .Z(n336) );
  INV_X1 U348 ( .A(KEYINPUT78), .ZN(n295) );
  NAND2_X1 U349 ( .A1(n295), .A2(KEYINPUT11), .ZN(n298) );
  INV_X1 U350 ( .A(KEYINPUT11), .ZN(n296) );
  NAND2_X1 U351 ( .A1(n296), .A2(KEYINPUT78), .ZN(n297) );
  NAND2_X1 U352 ( .A1(n298), .A2(n297), .ZN(n300) );
  XNOR2_X1 U353 ( .A(G218GAT), .B(G106GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n301) );
  NAND2_X1 U355 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n290), .B(n302), .ZN(n306) );
  XOR2_X1 U357 ( .A(KEYINPUT65), .B(G162GAT), .Z(n304) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(G134GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n314) );
  XOR2_X1 U361 ( .A(G92GAT), .B(KEYINPUT10), .Z(n308) );
  XNOR2_X1 U362 ( .A(KEYINPUT9), .B(KEYINPUT79), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U364 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n310) );
  XNOR2_X1 U365 ( .A(G190GAT), .B(G99GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U367 ( .A(n312), .B(n311), .Z(n313) );
  NAND2_X1 U368 ( .A1(n314), .A2(n313), .ZN(n318) );
  INV_X1 U369 ( .A(n313), .ZN(n316) );
  INV_X1 U370 ( .A(n314), .ZN(n315) );
  NAND2_X1 U371 ( .A1(n316), .A2(n315), .ZN(n317) );
  NAND2_X1 U372 ( .A1(n318), .A2(n317), .ZN(n319) );
  XOR2_X1 U373 ( .A(G169GAT), .B(G8GAT), .Z(n388) );
  XOR2_X1 U374 ( .A(G22GAT), .B(G1GAT), .Z(n354) );
  XOR2_X1 U375 ( .A(n388), .B(n354), .Z(n321) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U378 ( .A(G43GAT), .B(G15GAT), .Z(n455) );
  XOR2_X1 U379 ( .A(n322), .B(n455), .Z(n330) );
  XOR2_X1 U380 ( .A(KEYINPUT30), .B(G197GAT), .Z(n324) );
  XNOR2_X1 U381 ( .A(G113GAT), .B(G141GAT), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U383 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n326) );
  XNOR2_X1 U384 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n579) );
  XOR2_X1 U389 ( .A(G71GAT), .B(G120GAT), .Z(n334) );
  XNOR2_X1 U390 ( .A(G99GAT), .B(G176GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n450) );
  XNOR2_X1 U392 ( .A(G106GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n335), .B(G204GAT), .ZN(n435) );
  XNOR2_X1 U394 ( .A(n450), .B(n435), .ZN(n349) );
  XOR2_X1 U395 ( .A(n387), .B(n336), .Z(n338) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U398 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n340) );
  XNOR2_X1 U399 ( .A(KEYINPUT75), .B(KEYINPUT72), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U401 ( .A(n342), .B(n341), .Z(n347) );
  XOR2_X1 U402 ( .A(G148GAT), .B(G57GAT), .Z(n411) );
  XOR2_X1 U403 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n344) );
  XNOR2_X1 U404 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n411), .B(n345), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n583) );
  XNOR2_X1 U409 ( .A(KEYINPUT41), .B(n583), .ZN(n562) );
  NAND2_X1 U410 ( .A1(n579), .A2(n562), .ZN(n350) );
  XNOR2_X1 U411 ( .A(KEYINPUT46), .B(n350), .ZN(n369) );
  XOR2_X1 U412 ( .A(G71GAT), .B(G127GAT), .Z(n352) );
  XNOR2_X1 U413 ( .A(G15GAT), .B(G183GAT), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U415 ( .A(n354), .B(n353), .Z(n356) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U418 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n358) );
  XNOR2_X1 U419 ( .A(KEYINPUT80), .B(KEYINPUT15), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U421 ( .A(n360), .B(n359), .Z(n368) );
  XOR2_X1 U422 ( .A(G64GAT), .B(G78GAT), .Z(n362) );
  XNOR2_X1 U423 ( .A(G155GAT), .B(G211GAT), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U425 ( .A(KEYINPUT81), .B(KEYINPUT13), .Z(n364) );
  XNOR2_X1 U426 ( .A(G8GAT), .B(G57GAT), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n549) );
  NAND2_X1 U430 ( .A1(n369), .A2(n549), .ZN(n370) );
  NOR2_X1 U431 ( .A1(n373), .A2(n370), .ZN(n371) );
  XOR2_X1 U432 ( .A(KEYINPUT47), .B(n371), .Z(n382) );
  INV_X1 U433 ( .A(KEYINPUT104), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n374), .B(KEYINPUT36), .ZN(n590) );
  NOR2_X1 U436 ( .A1(n590), .A2(n549), .ZN(n376) );
  XOR2_X1 U437 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n579), .B(KEYINPUT70), .ZN(n570) );
  INV_X1 U440 ( .A(n583), .ZN(n377) );
  NOR2_X1 U441 ( .A1(n570), .A2(n377), .ZN(n378) );
  AND2_X1 U442 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n380), .B(KEYINPUT114), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n383), .B(KEYINPUT64), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n384), .B(KEYINPUT48), .ZN(n558) );
  XOR2_X1 U446 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n386) );
  XNOR2_X1 U447 ( .A(G204GAT), .B(KEYINPUT80), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n386), .B(n385), .ZN(n392) );
  XOR2_X1 U449 ( .A(n387), .B(G176GAT), .Z(n390) );
  XNOR2_X1 U450 ( .A(G36GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U452 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n400) );
  XOR2_X1 U455 ( .A(G211GAT), .B(KEYINPUT21), .Z(n396) );
  XNOR2_X1 U456 ( .A(G197GAT), .B(G218GAT), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n437) );
  XNOR2_X1 U458 ( .A(n437), .B(KEYINPUT99), .ZN(n398) );
  XNOR2_X1 U459 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n401), .B(KEYINPUT84), .ZN(n402) );
  XOR2_X1 U461 ( .A(n402), .B(KEYINPUT18), .Z(n404) );
  XNOR2_X1 U462 ( .A(G183GAT), .B(G190GAT), .ZN(n403) );
  XOR2_X1 U463 ( .A(n404), .B(n403), .Z(n461) );
  XNOR2_X1 U464 ( .A(n405), .B(n461), .ZN(n477) );
  NOR2_X1 U465 ( .A1(n558), .A2(n477), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n576) );
  XOR2_X1 U467 ( .A(KEYINPUT92), .B(KEYINPUT1), .Z(n409) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G120GAT), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U470 ( .A(n410), .B(G85GAT), .Z(n413) );
  XNOR2_X1 U471 ( .A(G29GAT), .B(n411), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n419) );
  XOR2_X1 U473 ( .A(G127GAT), .B(KEYINPUT0), .Z(n415) );
  XNOR2_X1 U474 ( .A(G113GAT), .B(G134GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n451) );
  XOR2_X1 U476 ( .A(n451), .B(KEYINPUT5), .Z(n417) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U479 ( .A(n419), .B(n418), .Z(n429) );
  XOR2_X1 U480 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n421) );
  XNOR2_X1 U481 ( .A(G162GAT), .B(KEYINPUT88), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U483 ( .A(n422), .B(KEYINPUT2), .Z(n424) );
  XNOR2_X1 U484 ( .A(G141GAT), .B(G155GAT), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n445) );
  XOR2_X1 U486 ( .A(KEYINPUT4), .B(KEYINPUT94), .Z(n426) );
  XNOR2_X1 U487 ( .A(KEYINPUT6), .B(KEYINPUT93), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n445), .B(n427), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n483) );
  XOR2_X1 U491 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n431) );
  XNOR2_X1 U492 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U494 ( .A(G50GAT), .B(KEYINPUT90), .Z(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n441) );
  XNOR2_X1 U496 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n434), .B(G148GAT), .ZN(n436) );
  XOR2_X1 U498 ( .A(n436), .B(n435), .Z(n439) );
  XNOR2_X1 U499 ( .A(G22GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n443) );
  NAND2_X1 U502 ( .A1(G228GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n486) );
  INV_X1 U505 ( .A(n486), .ZN(n446) );
  OR2_X1 U506 ( .A1(n575), .A2(n446), .ZN(n447) );
  XNOR2_X1 U507 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n462) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n459) );
  XOR2_X1 U510 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n453) );
  XNOR2_X1 U511 ( .A(G169GAT), .B(KEYINPUT83), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U513 ( .A(n455), .B(n454), .Z(n457) );
  NAND2_X1 U514 ( .A1(G227GAT), .A2(G233GAT), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n462), .A2(n540), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n572), .A2(n373), .ZN(n467) );
  XOR2_X1 U519 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n465) );
  INV_X1 U520 ( .A(G190GAT), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT109), .B(n562), .Z(n544) );
  NAND2_X1 U522 ( .A1(n572), .A2(n544), .ZN(n473) );
  XOR2_X1 U523 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n469) );
  XNOR2_X1 U524 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n468) );
  XNOR2_X1 U525 ( .A(n469), .B(n468), .ZN(n471) );
  XOR2_X1 U526 ( .A(G176GAT), .B(KEYINPUT56), .Z(n470) );
  XNOR2_X1 U527 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n473), .B(n472), .ZN(G1349GAT) );
  INV_X1 U529 ( .A(n477), .ZN(n533) );
  AND2_X1 U530 ( .A1(n540), .A2(n533), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(KEYINPUT101), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n475), .A2(n486), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(KEYINPUT25), .ZN(n480) );
  XOR2_X1 U534 ( .A(n477), .B(KEYINPUT27), .Z(n485) );
  NOR2_X1 U535 ( .A1(n540), .A2(n486), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT26), .B(n478), .ZN(n578) );
  AND2_X1 U537 ( .A1(n485), .A2(n578), .ZN(n479) );
  NOR2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n484) );
  NAND2_X1 U540 ( .A1(n484), .A2(n483), .ZN(n490) );
  NAND2_X1 U541 ( .A1(n485), .A2(n575), .ZN(n556) );
  XOR2_X1 U542 ( .A(KEYINPUT28), .B(n486), .Z(n537) );
  NOR2_X1 U543 ( .A1(n556), .A2(n537), .ZN(n541) );
  XNOR2_X1 U544 ( .A(KEYINPUT100), .B(n541), .ZN(n488) );
  XNOR2_X1 U545 ( .A(n540), .B(KEYINPUT85), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n489) );
  NAND2_X1 U547 ( .A1(n490), .A2(n489), .ZN(n502) );
  NAND2_X1 U548 ( .A1(n549), .A2(n502), .ZN(n491) );
  NOR2_X1 U549 ( .A1(n590), .A2(n491), .ZN(n494) );
  INV_X1 U550 ( .A(KEYINPUT37), .ZN(n492) );
  NAND2_X1 U551 ( .A1(n583), .A2(n570), .ZN(n504) );
  NOR2_X1 U552 ( .A1(n530), .A2(n504), .ZN(n496) );
  XNOR2_X1 U553 ( .A(KEYINPUT38), .B(KEYINPUT106), .ZN(n495) );
  NAND2_X1 U554 ( .A1(n516), .A2(n575), .ZN(n500) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT107), .Z(n498) );
  XOR2_X1 U556 ( .A(KEYINPUT39), .B(KEYINPUT108), .Z(n497) );
  XNOR2_X1 U557 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n506) );
  NOR2_X1 U558 ( .A1(n549), .A2(n373), .ZN(n501) );
  XNOR2_X1 U559 ( .A(n501), .B(KEYINPUT16), .ZN(n503) );
  NAND2_X1 U560 ( .A1(n503), .A2(n502), .ZN(n519) );
  NOR2_X1 U561 ( .A1(n504), .A2(n519), .ZN(n511) );
  NAND2_X1 U562 ( .A1(n511), .A2(n575), .ZN(n505) );
  XNOR2_X1 U563 ( .A(n506), .B(n505), .ZN(G1324GAT) );
  NAND2_X1 U564 ( .A1(n533), .A2(n511), .ZN(n507) );
  XNOR2_X1 U565 ( .A(n507), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n509) );
  NAND2_X1 U567 ( .A1(n511), .A2(n540), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U569 ( .A(G15GAT), .B(n510), .Z(G1326GAT) );
  NAND2_X1 U570 ( .A1(n537), .A2(n511), .ZN(n512) );
  XNOR2_X1 U571 ( .A(n512), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U572 ( .A1(n533), .A2(n516), .ZN(n513) );
  XNOR2_X1 U573 ( .A(n513), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U574 ( .A1(n540), .A2(n516), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n514), .B(KEYINPUT40), .ZN(n515) );
  XNOR2_X1 U576 ( .A(G43GAT), .B(n515), .ZN(G1330GAT) );
  NAND2_X1 U577 ( .A1(n537), .A2(n516), .ZN(n517) );
  XNOR2_X1 U578 ( .A(n517), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U579 ( .A(n579), .ZN(n518) );
  NAND2_X1 U580 ( .A1(n518), .A2(n544), .ZN(n529) );
  NOR2_X1 U581 ( .A1(n529), .A2(n519), .ZN(n520) );
  XNOR2_X1 U582 ( .A(KEYINPUT110), .B(n520), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n575), .A2(n526), .ZN(n521) );
  XNOR2_X1 U584 ( .A(KEYINPUT42), .B(n521), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G57GAT), .B(n522), .ZN(G1332GAT) );
  NAND2_X1 U586 ( .A1(n526), .A2(n533), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U588 ( .A(G71GAT), .B(KEYINPUT111), .Z(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n540), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .Z(n528) );
  NAND2_X1 U592 ( .A1(n526), .A2(n537), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n532) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n536), .A2(n575), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1336GAT) );
  NAND2_X1 U598 ( .A1(n533), .A2(n536), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n540), .A2(n536), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n538), .B(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U606 ( .A1(n558), .A2(n542), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n570), .A2(n552), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n543), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n546) );
  NAND2_X1 U610 ( .A1(n552), .A2(n544), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U612 ( .A(G120GAT), .B(KEYINPUT115), .Z(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  INV_X1 U614 ( .A(n549), .ZN(n587) );
  NAND2_X1 U615 ( .A1(n587), .A2(n552), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT50), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n554) );
  NAND2_X1 U619 ( .A1(n552), .A2(n373), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(G134GAT), .B(n555), .Z(G1343GAT) );
  INV_X1 U622 ( .A(n556), .ZN(n557) );
  NAND2_X1 U623 ( .A1(n578), .A2(n557), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n568) );
  AND2_X1 U625 ( .A1(n579), .A2(n568), .ZN(n560) );
  XOR2_X1 U626 ( .A(G141GAT), .B(n560), .Z(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT118), .B(n561), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n564) );
  NAND2_X1 U629 ( .A1(n568), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(n565), .ZN(G1345GAT) );
  XOR2_X1 U632 ( .A(G155GAT), .B(KEYINPUT119), .Z(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n587), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n373), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(G169GAT), .B(n571), .ZN(G1348GAT) );
  XOR2_X1 U639 ( .A(G183GAT), .B(KEYINPUT125), .Z(n574) );
  NAND2_X1 U640 ( .A1(n572), .A2(n587), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(G1350GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n581) );
  NOR2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n589) );
  INV_X1 U645 ( .A(n589), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n586), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  OR2_X1 U650 ( .A1(n589), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

