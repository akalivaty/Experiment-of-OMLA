//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G113gat), .B2(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT69), .B(G120gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT70), .B(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  OAI22_X1  g009(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT71), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n202), .B(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n206), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT79), .B1(new_n217), .B2(G148gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(G141gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n218), .B(new_n221), .C1(G141gat), .C2(new_n220), .ZN(new_n222));
  XNOR2_X1  g021(.A(G155gat), .B(G162gat), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  INV_X1    g023(.A(G162gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT2), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n223), .ZN(new_n228));
  XNOR2_X1  g027(.A(G141gat), .B(G148gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(KEYINPUT2), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT80), .B1(new_n216), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n227), .A2(new_n230), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n202), .B(KEYINPUT71), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(new_n212), .A3(new_n211), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n233), .A2(new_n235), .A3(new_n236), .A4(new_n206), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n231), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT84), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT84), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n233), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT3), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n216), .A3(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n237), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n211), .A2(new_n212), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n250), .A2(new_n234), .B1(new_n203), .B2(new_n205), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .A4(new_n233), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n233), .A2(new_n235), .A3(new_n253), .A4(new_n206), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT82), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n248), .B1(new_n249), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n244), .B1(new_n258), .B2(new_n241), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n243), .B(KEYINPUT39), .C1(new_n259), .C2(new_n242), .ZN(new_n260));
  XNOR2_X1  g059(.A(G1gat), .B(G29gat), .ZN(new_n261));
  INV_X1    g060(.A(G85gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G57gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT39), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n258), .A2(new_n266), .A3(new_n241), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n260), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT40), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT77), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT22), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT76), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(KEYINPUT76), .ZN(new_n278));
  INV_X1    g077(.A(G211gat), .ZN(new_n279));
  INV_X1    g078(.A(G218gat), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n275), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G226gat), .A2(G233gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT23), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n291), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT66), .B(G190gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(G183gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n293), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT25), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n297), .A2(KEYINPUT64), .ZN(new_n303));
  INV_X1    g102(.A(new_n296), .ZN(new_n304));
  OR2_X1    g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(KEYINPUT64), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT25), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n293), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT26), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n290), .B1(new_n287), .B2(new_n310), .ZN(new_n311));
  NOR3_X1   g110(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n294), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT68), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT66), .B(G190gat), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(G183gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT27), .B(G183gat), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n315), .B(new_n318), .C1(new_n316), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n299), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n320), .A2(new_n321), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n302), .B(new_n309), .C1(new_n314), .C2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n286), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n307), .A2(new_n308), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n327), .A2(new_n293), .B1(new_n301), .B2(KEYINPUT25), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT68), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n313), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n320), .A2(new_n321), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(new_n319), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n285), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n284), .B1(new_n326), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n324), .A2(new_n286), .ZN(new_n337));
  INV_X1    g136(.A(new_n284), .ZN(new_n338));
  XOR2_X1   g137(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(new_n328), .B2(new_n334), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n337), .B(new_n338), .C1(new_n340), .C2(new_n286), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n273), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n341), .A3(new_n273), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(KEYINPUT30), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n336), .A2(new_n341), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n347));
  INV_X1    g146(.A(new_n273), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n232), .A2(new_n253), .A3(new_n237), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n216), .A2(new_n231), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n241), .B1(new_n353), .B2(KEYINPUT4), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n354), .A3(new_n248), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n239), .A2(new_n241), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n241), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n248), .B(new_n359), .C1(new_n249), .C2(new_n257), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n265), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT85), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n260), .A2(KEYINPUT40), .A3(new_n265), .A4(new_n267), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n270), .A2(new_n351), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n339), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n284), .B1(new_n246), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(G228gat), .B2(G233gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT3), .B1(new_n284), .B2(new_n365), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n233), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n284), .A2(new_n325), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n233), .B1(new_n370), .B2(new_n245), .ZN(new_n371));
  OAI211_X1 g170(.A(G228gat), .B(G233gat), .C1(new_n371), .C2(new_n366), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G78gat), .B(G106gat), .Z(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(G22gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT31), .B(G50gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n373), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n358), .A2(new_n360), .A3(new_n265), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n361), .A2(KEYINPUT85), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n361), .A2(KEYINPUT85), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n361), .A2(KEYINPUT6), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT37), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n348), .B1(new_n346), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n386), .B2(new_n346), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n342), .B1(new_n388), .B2(KEYINPUT38), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT38), .ZN(new_n390));
  OR3_X1    g189(.A1(new_n326), .A2(new_n335), .A3(new_n284), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n337), .B1(new_n340), .B2(new_n286), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n284), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n393), .A3(KEYINPUT37), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n384), .A2(new_n385), .A3(new_n389), .A4(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n364), .A2(new_n379), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT75), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT36), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(KEYINPUT75), .A2(KEYINPUT36), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n324), .A2(new_n216), .ZN(new_n402));
  INV_X1    g201(.A(G227gat), .ZN(new_n403));
  INV_X1    g202(.A(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n328), .A2(new_n334), .A3(new_n251), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT74), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n408), .A2(KEYINPUT34), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n408), .A2(KEYINPUT74), .A3(new_n409), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n402), .A2(new_n407), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n405), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT32), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G15gat), .B(G43gat), .ZN(new_n423));
  INV_X1    g222(.A(G71gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT72), .B(G99gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n418), .A4(new_n414), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n420), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n420), .B2(new_n430), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n400), .B(new_n401), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n420), .A2(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n428), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n429), .A3(new_n430), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n435), .A2(new_n398), .A3(new_n399), .A4(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n381), .A2(new_n380), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n385), .B1(new_n439), .B2(new_n361), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n440), .A2(KEYINPUT83), .A3(new_n350), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT83), .B1(new_n440), .B2(new_n350), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n378), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n397), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n431), .A2(new_n432), .A3(new_n378), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT35), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n384), .A2(new_n385), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n350), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n435), .A2(new_n379), .A3(new_n436), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n449), .A2(new_n441), .A3(new_n442), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n450), .B2(new_n446), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT88), .ZN(new_n455));
  AND2_X1   g254(.A1(G15gat), .A2(G22gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(G15gat), .A2(G22gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G1gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G15gat), .B(G22gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n455), .A3(G1gat), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT16), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G8gat), .ZN(new_n466));
  INV_X1    g265(.A(G8gat), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n460), .A2(new_n462), .A3(new_n467), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G183gat), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT21), .ZN(new_n472));
  XOR2_X1   g271(.A(G57gat), .B(G64gat), .Z(new_n473));
  INV_X1    g272(.A(KEYINPUT9), .ZN(new_n474));
  INV_X1    g273(.A(G78gat), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n474), .B1(new_n424), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G71gat), .B(G78gat), .Z(new_n478));
  OR2_X1    g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n472), .ZN(new_n483));
  OAI21_X1  g282(.A(G183gat), .B1(new_n483), .B2(new_n469), .ZN(new_n484));
  NAND2_X1  g283(.A1(G231gat), .A2(G233gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n485), .B(KEYINPUT91), .Z(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n482), .B2(new_n484), .ZN(new_n490));
  INV_X1    g289(.A(new_n481), .ZN(new_n491));
  OAI22_X1  g290(.A1(new_n489), .A2(new_n490), .B1(KEYINPUT21), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n490), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(KEYINPUT21), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n488), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n454), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(G211gat), .ZN(new_n499));
  XOR2_X1   g298(.A(G127gat), .B(G155gat), .Z(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n492), .A2(new_n495), .A3(new_n454), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n497), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n501), .ZN(new_n504));
  INV_X1    g303(.A(new_n502), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(new_n496), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G134gat), .B(G162gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT95), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT41), .ZN(new_n510));
  INV_X1    g309(.A(G232gat), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(new_n404), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n509), .B(new_n512), .Z(new_n513));
  NAND2_X1  g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514));
  INV_X1    g313(.A(G92gat), .ZN(new_n515));
  AOI22_X1  g314(.A1(KEYINPUT8), .A2(new_n514), .B1(new_n262), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT7), .ZN(new_n517));
  OAI22_X1  g316(.A1(new_n262), .A2(new_n515), .B1(new_n517), .B2(KEYINPUT94), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G99gat), .B(G106gat), .Z(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G50gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G43gat), .ZN(new_n532));
  INV_X1    g331(.A(G43gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G50gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT15), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n532), .A2(new_n534), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT15), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n535), .A3(new_n526), .ZN(new_n541));
  NOR4_X1   g340(.A1(KEYINPUT86), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT86), .ZN(new_n543));
  NOR2_X1   g342(.A1(G29gat), .A2(G36gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n542), .A2(new_n546), .A3(new_n528), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n537), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT87), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT87), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n550), .B(new_n537), .C1(new_n541), .C2(new_n547), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT17), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n548), .A2(KEYINPUT17), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n525), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n551), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n525), .ZN(new_n557));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n513), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n513), .A3(new_n560), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n479), .A2(new_n523), .A3(new_n480), .A4(new_n524), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT10), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n481), .A2(new_n525), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n566), .A3(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n568), .B2(new_n565), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n570), .A2(new_n571), .B1(KEYINPUT96), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G120gat), .B(G148gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n572), .A2(KEYINPUT96), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n573), .B2(new_n578), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n507), .A2(new_n564), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n549), .A2(new_n469), .A3(new_n551), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT89), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n549), .A2(new_n469), .A3(KEYINPUT89), .A4(new_n551), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n470), .B1(new_n552), .B2(new_n553), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT18), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G197gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT11), .B(G169gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT12), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n588), .A2(new_n590), .A3(KEYINPUT18), .A4(new_n589), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n556), .A2(new_n470), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n588), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n589), .B(KEYINPUT13), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n600), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n588), .A2(new_n602), .ZN(new_n609));
  INV_X1    g408(.A(new_n604), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n608), .A2(KEYINPUT18), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n593), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n599), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n452), .A2(new_n583), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n440), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT97), .B(G1gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(G1324gat));
  AOI21_X1  g418(.A(new_n467), .B1(new_n615), .B2(new_n351), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n620), .B(KEYINPUT99), .Z(new_n621));
  NAND2_X1  g420(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n463), .A2(new_n467), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n615), .A2(new_n351), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT42), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT42), .B1(new_n624), .B2(new_n625), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(G1325gat));
  NOR2_X1   g427(.A1(new_n431), .A2(new_n432), .ZN(new_n629));
  AOI21_X1  g428(.A(G15gat), .B1(new_n615), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n433), .A2(new_n437), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n634), .A2(G15gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n630), .B1(new_n615), .B2(new_n635), .ZN(G1326gat));
  NAND2_X1  g435(.A1(new_n615), .A2(new_n378), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT43), .B(G22gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(G1327gat));
  NAND2_X1  g438(.A1(new_n444), .A2(new_n451), .ZN(new_n640));
  INV_X1    g439(.A(new_n564), .ZN(new_n641));
  INV_X1    g440(.A(new_n614), .ZN(new_n642));
  INV_X1    g441(.A(new_n582), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n507), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n640), .A2(new_n641), .A3(new_n642), .A4(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n645), .A2(G29gat), .A3(new_n440), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT45), .Z(new_n647));
  OAI21_X1  g446(.A(KEYINPUT101), .B1(new_n607), .B2(new_n613), .ZN(new_n648));
  INV_X1    g447(.A(new_n606), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n649), .A2(new_n611), .A3(new_n599), .A4(new_n594), .ZN(new_n650));
  INV_X1    g449(.A(new_n599), .ZN(new_n651));
  INV_X1    g450(.A(new_n612), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n605), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT103), .B1(new_n562), .B2(new_n563), .ZN(new_n657));
  INV_X1    g456(.A(new_n563), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n658), .A2(new_n659), .A3(new_n561), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n443), .A2(KEYINPUT102), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n663), .B(new_n378), .C1(new_n441), .C2(new_n442), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n662), .A2(new_n397), .A3(new_n438), .A4(new_n664), .ZN(new_n665));
  AOI211_X1 g464(.A(KEYINPUT44), .B(new_n661), .C1(new_n665), .C2(new_n451), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n640), .B2(new_n641), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n656), .B(new_n644), .C1(new_n666), .C2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(G29gat), .B1(new_n669), .B2(new_n440), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n647), .A2(new_n670), .ZN(G1328gat));
  OAI21_X1  g470(.A(G36gat), .B1(new_n669), .B2(new_n350), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n645), .A2(G36gat), .A3(new_n350), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n673), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n675), .A2(KEYINPUT104), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(KEYINPUT104), .ZN(new_n677));
  OAI221_X1 g476(.A(new_n672), .B1(new_n673), .B2(new_n674), .C1(new_n676), .C2(new_n677), .ZN(G1329gat));
  INV_X1    g477(.A(new_n629), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n645), .A2(G43gat), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT47), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(KEYINPUT105), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G43gat), .B1(new_n669), .B2(new_n438), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  INV_X1    g483(.A(new_n669), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n533), .B1(new_n685), .B2(new_n634), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(KEYINPUT105), .B2(new_n680), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n684), .B1(new_n687), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g487(.A(G50gat), .B1(new_n669), .B2(new_n379), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n645), .A2(G50gat), .A3(new_n379), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n690), .B1(new_n689), .B2(new_n692), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT48), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n689), .A2(new_n692), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT106), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT48), .B1(new_n699), .B2(new_n693), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n697), .A2(new_n700), .ZN(G1331gat));
  INV_X1    g500(.A(new_n507), .ZN(new_n702));
  AOI211_X1 g501(.A(new_n702), .B(new_n641), .C1(new_n665), .C2(new_n451), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n656), .A2(new_n582), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n616), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g507(.A1(new_n705), .A2(new_n350), .ZN(new_n709));
  NOR2_X1   g508(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n710));
  AND2_X1   g509(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n709), .B2(new_n710), .ZN(G1333gat));
  NAND3_X1  g512(.A1(new_n706), .A2(new_n424), .A3(new_n629), .ZN(new_n714));
  OAI21_X1  g513(.A(G71gat), .B1(new_n705), .B2(new_n633), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g516(.A1(new_n705), .A2(new_n379), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n475), .ZN(G1335gat));
  OAI211_X1 g518(.A(new_n702), .B(new_n704), .C1(new_n666), .C2(new_n668), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(new_n262), .A3(new_n440), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n665), .A2(new_n451), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n656), .A2(new_n507), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(new_n641), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n722), .A2(KEYINPUT51), .A3(new_n641), .A4(new_n723), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n728), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT107), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n729), .A2(new_n731), .A3(new_n616), .A4(new_n643), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n721), .B1(new_n732), .B2(new_n262), .ZN(G1336gat));
  NOR2_X1   g532(.A1(new_n350), .A2(G92gat), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n729), .A2(new_n731), .A3(new_n643), .A4(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736));
  OAI21_X1  g535(.A(G92gat), .B1(new_n720), .B2(new_n350), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n726), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n643), .B(new_n734), .C1(new_n740), .C2(new_n730), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n736), .B1(new_n741), .B2(new_n737), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n741), .A2(new_n737), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n738), .B(new_n744), .C1(new_n745), .C2(new_n736), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1337gat));
  OR3_X1    g546(.A1(new_n720), .A2(KEYINPUT109), .A3(new_n633), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT109), .B1(new_n720), .B2(new_n633), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(G99gat), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n679), .A2(G99gat), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n729), .A2(new_n731), .A3(new_n643), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1338gat));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT110), .B(G106gat), .Z(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n720), .B2(new_n379), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n379), .A2(new_n582), .A3(G106gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n729), .A2(new_n731), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n754), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AND4_X1   g560(.A1(new_n754), .A2(new_n760), .A3(new_n756), .A4(new_n757), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n740), .B2(new_n730), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n756), .A2(new_n763), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n761), .A2(new_n762), .B1(new_n757), .B2(new_n764), .ZN(G1339gat));
  NOR2_X1   g564(.A1(new_n583), .A2(new_n656), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n657), .A2(new_n660), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n570), .A2(new_n571), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n567), .A2(new_n569), .A3(G230gat), .A4(G233gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(KEYINPUT54), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n577), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n768), .A2(KEYINPUT54), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n768), .A2(KEYINPUT112), .A3(KEYINPUT54), .A4(new_n769), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n772), .A2(KEYINPUT55), .A3(new_n773), .A4(new_n774), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n579), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n603), .B2(new_n604), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n781), .A2(new_n598), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n650), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n783), .A2(new_n582), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n777), .A2(new_n579), .A3(new_n778), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n656), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n788), .B2(new_n767), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n766), .B1(new_n789), .B2(new_n702), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT113), .B1(new_n790), .B2(new_n378), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n779), .B1(new_n648), .B2(new_n655), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n661), .B1(new_n793), .B2(new_n786), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n507), .B1(new_n794), .B2(new_n785), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n792), .B(new_n379), .C1(new_n795), .C2(new_n766), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n351), .A2(new_n440), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n791), .A2(new_n629), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n207), .B1(new_n800), .B2(new_n642), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n790), .A2(new_n449), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n797), .ZN(new_n803));
  INV_X1    g602(.A(new_n656), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n803), .A2(new_n209), .A3(new_n804), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n801), .A2(new_n805), .ZN(G1340gat));
  AOI21_X1  g605(.A(new_n210), .B1(new_n800), .B2(new_n643), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n803), .A2(new_n208), .A3(new_n582), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n807), .A2(new_n808), .ZN(G1341gat));
  NAND3_X1  g608(.A1(new_n800), .A2(G127gat), .A3(new_n507), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n800), .A2(KEYINPUT115), .A3(G127gat), .A4(new_n507), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n802), .A2(new_n507), .A3(new_n797), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(KEYINPUT116), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(KEYINPUT116), .ZN(new_n816));
  OR3_X1    g615(.A1(new_n815), .A2(new_n816), .A3(G127gat), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n812), .A2(new_n813), .A3(new_n817), .ZN(G1342gat));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819));
  INV_X1    g618(.A(G134gat), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n800), .B2(new_n641), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n802), .A2(new_n820), .A3(new_n641), .A4(new_n797), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT56), .Z(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n819), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n791), .A2(new_n629), .A3(new_n796), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n799), .A3(new_n797), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n798), .A2(KEYINPUT114), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n641), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G134gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(KEYINPUT117), .A3(new_n823), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n825), .A2(new_n831), .ZN(G1343gat));
  NAND2_X1  g631(.A1(new_n438), .A2(new_n797), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT118), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n779), .A2(new_n614), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n564), .B1(new_n835), .B2(new_n786), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n507), .B1(new_n836), .B2(new_n785), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n378), .B1(new_n837), .B2(new_n766), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n834), .B1(KEYINPUT57), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n790), .A2(new_n379), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G141gat), .B1(new_n843), .B2(new_n614), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n840), .A2(new_n633), .A3(new_n797), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n217), .A3(new_n642), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G141gat), .B1(new_n843), .B2(new_n804), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(new_n846), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n850), .B2(new_n847), .ZN(G1344gat));
  NAND3_X1  g650(.A1(new_n845), .A2(new_n220), .A3(new_n643), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(G148gat), .C1(new_n843), .C2(new_n582), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT119), .ZN(new_n855));
  XNOR2_X1  g654(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT57), .B1(new_n790), .B2(new_n379), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n784), .A2(new_n641), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n507), .B1(new_n836), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n583), .A2(new_n642), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n841), .B(new_n378), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n643), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(new_n834), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n856), .B1(new_n865), .B2(G148gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n852), .B1(new_n855), .B2(new_n866), .ZN(G1345gat));
  NOR3_X1   g666(.A1(new_n843), .A2(new_n224), .A3(new_n702), .ZN(new_n868));
  AOI21_X1  g667(.A(G155gat), .B1(new_n845), .B2(new_n507), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(G1346gat));
  OAI21_X1  g669(.A(G162gat), .B1(new_n843), .B2(new_n661), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n845), .A2(new_n225), .A3(new_n641), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1347gat));
  NOR2_X1   g672(.A1(new_n616), .A2(new_n350), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n802), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(G169gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n656), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT121), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n791), .A2(new_n629), .A3(new_n796), .A4(new_n874), .ZN(new_n879));
  OAI21_X1  g678(.A(G169gat), .B1(new_n879), .B2(new_n614), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT122), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n878), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1348gat));
  AOI21_X1  g684(.A(G176gat), .B1(new_n875), .B2(new_n643), .ZN(new_n886));
  INV_X1    g685(.A(new_n879), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n643), .A2(G176gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(G1349gat));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(KEYINPUT60), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(KEYINPUT60), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n826), .A2(KEYINPUT123), .A3(new_n507), .A4(new_n874), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n894), .B1(new_n879), .B2(new_n702), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(G183gat), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n875), .A2(new_n507), .A3(new_n319), .ZN(new_n897));
  AOI211_X1 g696(.A(new_n891), .B(new_n892), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  AND4_X1   g697(.A1(new_n890), .A2(new_n896), .A3(KEYINPUT60), .A4(new_n897), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n875), .A2(new_n315), .A3(new_n767), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n826), .A2(new_n641), .A3(new_n874), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(G190gat), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n902), .B(G190gat), .C1(new_n879), .C2(new_n564), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n901), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n909), .B(new_n901), .C1(new_n904), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1351gat));
  AND2_X1   g710(.A1(new_n633), .A2(new_n874), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT127), .Z(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n862), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n642), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G197gat), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n840), .A2(new_n912), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(G197gat), .A3(new_n804), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT126), .Z(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1352gat));
  NOR3_X1   g719(.A1(new_n917), .A2(G204gat), .A3(new_n582), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT62), .ZN(new_n922));
  OAI21_X1  g721(.A(G204gat), .B1(new_n864), .B2(new_n913), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1353gat));
  NOR2_X1   g723(.A1(new_n862), .A2(new_n702), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n279), .B1(new_n925), .B2(new_n912), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(KEYINPUT63), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(KEYINPUT63), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n507), .A2(new_n279), .ZN(new_n929));
  OAI22_X1  g728(.A1(new_n927), .A2(new_n928), .B1(new_n917), .B2(new_n929), .ZN(G1354gat));
  NAND3_X1  g729(.A1(new_n914), .A2(G218gat), .A3(new_n641), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n280), .B1(new_n917), .B2(new_n661), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(G1355gat));
endmodule


