//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003;
  XNOR2_X1  g000(.A(G134gat), .B(G162gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  AND2_X1   g003(.A1(G232gat), .A2(G233gat), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n205), .A2(KEYINPUT41), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT92), .B(G50gat), .Z(new_n208));
  INV_X1    g007(.A(KEYINPUT93), .ZN(new_n209));
  INV_X1    g008(.A(G43gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n210), .A2(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(new_n208), .B2(new_n210), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n207), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n210), .A2(G50gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT14), .ZN(new_n221));
  NAND2_X1  g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n215), .A2(new_n217), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n217), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(KEYINPUT91), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n222), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n221), .A2(KEYINPUT91), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n224), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT7), .ZN(new_n231));
  INV_X1    g030(.A(G99gat), .ZN(new_n232));
  INV_X1    g031(.A(G106gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT8), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n231), .B(new_n234), .C1(G85gat), .C2(G92gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(G99gat), .B(G106gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n206), .B1(new_n229), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT101), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n237), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(new_n223), .B2(new_n228), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT101), .B1(new_n242), .B2(new_n206), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n223), .A2(new_n245), .A3(new_n228), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n223), .B2(new_n228), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n241), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT100), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT100), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n251), .B(new_n241), .C1(new_n247), .C2(new_n248), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n205), .A2(KEYINPUT41), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n254), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n244), .A2(new_n250), .A3(new_n256), .A4(new_n252), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n204), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(new_n204), .A3(new_n257), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n202), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n260), .ZN(new_n262));
  INV_X1    g061(.A(new_n202), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n262), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G15gat), .B(G22gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT16), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n266), .B1(new_n267), .B2(G1gat), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n268), .A2(KEYINPUT94), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n266), .A2(G1gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n268), .A3(KEYINPUT94), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n271), .A3(G8gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT95), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n269), .A2(new_n271), .A3(KEYINPUT95), .A4(G8gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G8gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n268), .A3(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G57gat), .B(G64gat), .Z(new_n279));
  NAND2_X1  g078(.A1(G71gat), .A2(G78gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT9), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G71gat), .B(G78gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT21), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(new_n278), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT99), .ZN(new_n288));
  AND2_X1   g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G127gat), .B(G155gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT20), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n285), .A2(KEYINPUT21), .ZN(new_n294));
  XNOR2_X1  g093(.A(G183gat), .B(G211gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT98), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT19), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n294), .B(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n292), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n293), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n293), .B2(new_n299), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G230gat), .ZN(new_n303));
  INV_X1    g102(.A(G233gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n236), .A2(KEYINPUT102), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n285), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n236), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n235), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n235), .A2(new_n308), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n237), .A2(new_n285), .A3(new_n306), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT10), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n237), .A2(KEYINPUT10), .A3(new_n285), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n305), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n311), .A2(new_n312), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n305), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G120gat), .B(G148gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G176gat), .B(G204gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n323), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n317), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n265), .A2(new_n302), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT76), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT66), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(KEYINPUT67), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(new_n335), .B2(new_n336), .ZN(new_n343));
  INV_X1    g142(.A(new_n339), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT65), .B(KEYINPUT23), .Z(new_n346));
  INV_X1    g145(.A(new_n333), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n340), .A2(new_n345), .A3(KEYINPUT25), .A4(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G183gat), .ZN(new_n350));
  INV_X1    g149(.A(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(KEYINPUT24), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(KEYINPUT24), .B2(new_n353), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT64), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n333), .A2(KEYINPUT23), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(KEYINPUT64), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n355), .A2(new_n344), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT25), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT27), .B(G183gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(KEYINPUT28), .A3(new_n351), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT70), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n365), .A2(KEYINPUT70), .A3(KEYINPUT28), .A4(new_n351), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT28), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT68), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n350), .A2(KEYINPUT27), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G183gat), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n371), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n371), .B1(new_n373), .B2(G183gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n351), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n370), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT69), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(KEYINPUT69), .B(new_n370), .C1(new_n375), .C2(new_n377), .ZN(new_n381));
  AOI221_X4 g180(.A(KEYINPUT71), .B1(new_n368), .B2(new_n369), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT71), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n381), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT26), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n337), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n344), .B1(new_n347), .B2(KEYINPUT26), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n389), .A2(new_n390), .B1(G183gat), .B2(G190gat), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n364), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n332), .B1(new_n392), .B2(KEYINPUT29), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(new_n392), .B2(new_n332), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n351), .B(new_n376), .C1(new_n365), .C2(new_n371), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT69), .B1(new_n396), .B2(new_n370), .ZN(new_n397));
  INV_X1    g196(.A(new_n381), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n385), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT71), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n383), .A3(new_n385), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n391), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n360), .A2(new_n362), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n403), .A2(KEYINPUT25), .B1(new_n355), .B2(new_n349), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n332), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT77), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n393), .A2(new_n395), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G197gat), .B(G204gat), .ZN(new_n408));
  INV_X1    g207(.A(G211gat), .ZN(new_n409));
  INV_X1    g208(.A(G218gat), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n408), .A2(KEYINPUT22), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n409), .B2(new_n410), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT22), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n409), .A2(new_n410), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n408), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n407), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n404), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n331), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n420), .A2(new_n416), .A3(new_n405), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n417), .A2(KEYINPUT30), .A3(new_n422), .A4(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n416), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT77), .B1(new_n418), .B2(new_n331), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n394), .B(new_n332), .C1(new_n402), .C2(new_n404), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n431), .B2(new_n393), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n425), .B1(new_n432), .B2(new_n421), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT78), .ZN(new_n435));
  INV_X1    g234(.A(G120gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G113gat), .ZN(new_n437));
  INV_X1    g236(.A(G113gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G120gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT1), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(G127gat), .B(G134gat), .Z(new_n443));
  AND2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n443), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT72), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n438), .B2(G120gat), .ZN(new_n448));
  MUX2_X1   g247(.A(new_n447), .B(new_n448), .S(new_n437), .Z(new_n449));
  INV_X1    g248(.A(KEYINPUT73), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n437), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT72), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n448), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n441), .B1(new_n454), .B2(KEYINPUT73), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n445), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(G141gat), .B(G148gat), .Z(new_n457));
  INV_X1    g256(.A(KEYINPUT2), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460));
  NAND2_X1  g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461));
  OR2_X1    g260(.A1(G155gat), .A2(G162gat), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(KEYINPUT2), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n457), .ZN(new_n465));
  XNOR2_X1  g264(.A(G141gat), .B(G148gat), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n461), .B(new_n462), .C1(new_n466), .C2(KEYINPUT2), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT80), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT82), .B1(new_n456), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT1), .B1(new_n449), .B2(new_n450), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n443), .B1(new_n454), .B2(KEYINPUT73), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n444), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT82), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n470), .B(new_n476), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT81), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT3), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n475), .B2(new_n483), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n469), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n456), .B(new_n481), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n473), .A2(new_n475), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n480), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT5), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n456), .A2(new_n469), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n476), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n493), .B2(new_n479), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n477), .B1(new_n470), .B2(new_n476), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n487), .A2(new_n477), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n479), .A2(KEYINPUT5), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n497), .A2(new_n486), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G57gat), .B(G85gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G1gat), .B(G29gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n504), .B(new_n505), .Z(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n495), .A2(new_n500), .A3(new_n506), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(KEYINPUT6), .A3(new_n507), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n417), .A2(new_n422), .A3(new_n426), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT78), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n427), .A2(new_n433), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n435), .A2(new_n513), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT32), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n418), .B(new_n456), .ZN(new_n522));
  INV_X1    g321(.A(G227gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(new_n304), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n522), .A2(KEYINPUT34), .A3(new_n524), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT34), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n418), .B(new_n473), .ZN(new_n528));
  INV_X1    g327(.A(new_n524), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n525), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT32), .B1(new_n528), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT34), .B1(new_n522), .B2(new_n524), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n527), .A3(new_n529), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT74), .B(G71gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(new_n232), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G43gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n538), .B(new_n539), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n524), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT33), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n536), .A2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n415), .A2(KEYINPUT84), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n415), .A2(KEYINPUT84), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n412), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n419), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n475), .B1(new_n550), .B2(new_n483), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n419), .B1(new_n484), .B2(new_n485), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(new_n416), .ZN(new_n553));
  AND2_X1   g352(.A1(G228gat), .A2(G233gat), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT85), .B(G22gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n483), .B1(new_n416), .B2(KEYINPUT29), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n469), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n475), .A2(new_n482), .A3(new_n483), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT81), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT29), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n554), .B(new_n559), .C1(new_n562), .C2(new_n428), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(new_n557), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT87), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n563), .B1(new_n553), .B2(new_n554), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT86), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT86), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n563), .B(new_n569), .C1(new_n553), .C2(new_n554), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(G22gat), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n555), .A2(KEYINPUT87), .A3(new_n557), .A4(new_n563), .ZN(new_n572));
  XNOR2_X1  g371(.A(G78gat), .B(G106gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT31), .B(G50gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n566), .A2(new_n571), .A3(new_n572), .A4(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  INV_X1    g376(.A(new_n564), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n567), .A2(new_n556), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n531), .A2(new_n535), .A3(new_n544), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n546), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT35), .B1(new_n520), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n582), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n544), .B1(new_n531), .B2(new_n535), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n421), .B1(new_n407), .B2(new_n416), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n515), .B1(new_n588), .B2(new_n426), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n434), .A2(new_n589), .A3(KEYINPUT35), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n587), .A2(new_n590), .A3(new_n513), .A4(new_n581), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT37), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(new_n432), .B2(new_n421), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n417), .A2(KEYINPUT37), .A3(new_n422), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n425), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT89), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT38), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n511), .A2(new_n514), .A3(new_n512), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n416), .B1(new_n420), .B2(new_n405), .ZN(new_n601));
  OAI211_X1 g400(.A(KEYINPUT37), .B(new_n601), .C1(new_n407), .C2(new_n416), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT38), .B1(new_n594), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n600), .B1(new_n603), .B2(new_n425), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n426), .B1(new_n594), .B2(new_n595), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT38), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT89), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n493), .A2(new_n479), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n456), .A2(new_n481), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n561), .B2(new_n560), .ZN(new_n611));
  INV_X1    g410(.A(new_n498), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n496), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(KEYINPUT39), .B(new_n609), .C1(new_n613), .C2(new_n478), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n497), .A2(new_n486), .A3(new_n498), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n616), .A3(new_n479), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n506), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT88), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(KEYINPUT40), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n618), .A2(new_n620), .B1(new_n507), .B2(new_n501), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n621), .B(new_n622), .C1(new_n434), .C2(new_n589), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n623), .A2(new_n581), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n608), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(KEYINPUT75), .B(KEYINPUT36), .C1(new_n585), .C2(new_n586), .ZN(new_n626));
  NAND2_X1  g425(.A1(KEYINPUT75), .A2(KEYINPUT36), .ZN(new_n627));
  OR2_X1    g426(.A1(KEYINPUT75), .A2(KEYINPUT36), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n546), .A2(new_n627), .A3(new_n628), .A4(new_n582), .ZN(new_n629));
  INV_X1    g428(.A(new_n519), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n513), .A2(new_n517), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n518), .B1(new_n427), .B2(new_n433), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n626), .B(new_n629), .C1(new_n633), .C2(new_n581), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n592), .B1(new_n625), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT90), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n608), .A2(new_n624), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n626), .A2(new_n629), .ZN(new_n639));
  INV_X1    g438(.A(new_n581), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n520), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(KEYINPUT90), .A3(new_n592), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT18), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n229), .A2(KEYINPUT17), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n276), .A2(new_n278), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n645), .A2(new_n246), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n276), .A2(KEYINPUT96), .A3(new_n278), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n229), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G229gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n644), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n651), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n646), .A2(new_n229), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n653), .B(KEYINPUT13), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n656), .B1(new_n648), .B2(new_n649), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(KEYINPUT18), .A3(new_n653), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n655), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G113gat), .B(G141gat), .ZN(new_n664));
  INV_X1    g463(.A(G197gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT11), .B(G169gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT12), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n669), .A3(new_n660), .A4(new_n662), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n637), .A2(new_n643), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT97), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT97), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n637), .A2(new_n676), .A3(new_n643), .A4(new_n673), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n329), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n513), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g480(.A1(new_n675), .A2(new_n677), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n434), .A2(new_n589), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n329), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G8gat), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n682), .A2(new_n684), .A3(new_n685), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n678), .A2(new_n684), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G8gat), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(KEYINPUT103), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(G1325gat));
  AOI21_X1  g494(.A(G15gat), .B1(new_n678), .B2(new_n587), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n626), .A2(new_n629), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n697), .A2(G15gat), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n678), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n678), .A2(new_n640), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  INV_X1    g501(.A(new_n302), .ZN(new_n703));
  INV_X1    g502(.A(new_n265), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n328), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT105), .Z(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n675), .B2(new_n677), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n218), .A3(new_n679), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(KEYINPUT45), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710));
  INV_X1    g509(.A(new_n643), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT90), .B1(new_n642), .B2(new_n592), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n265), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n584), .A2(KEYINPUT107), .A3(new_n591), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT107), .B1(new_n584), .B2(new_n591), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n630), .A2(new_n632), .ZN(new_n719));
  INV_X1    g518(.A(new_n631), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n581), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n639), .B1(new_n721), .B2(KEYINPUT106), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n520), .A2(KEYINPUT106), .A3(new_n640), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n638), .A2(new_n723), .ZN(new_n724));
  OAI22_X1  g523(.A1(new_n717), .A2(new_n718), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n704), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n713), .A2(new_n715), .B1(new_n726), .B2(new_n714), .ZN(new_n727));
  INV_X1    g526(.A(new_n673), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n302), .A2(new_n728), .A3(new_n327), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n727), .A2(new_n679), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n710), .B1(new_n730), .B2(G29gat), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n709), .B1(new_n708), .B2(new_n731), .ZN(G1328gat));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n707), .A2(new_n733), .A3(new_n219), .A4(new_n684), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n592), .A2(new_n735), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n721), .A2(KEYINPUT106), .B1(new_n608), .B2(new_n624), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n697), .B1(new_n641), .B2(new_n738), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n736), .A2(new_n716), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n714), .B1(new_n740), .B2(new_n265), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n637), .A2(new_n643), .A3(new_n715), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n741), .A2(new_n742), .A3(new_n684), .A4(new_n729), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G36gat), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n706), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n682), .A2(new_n219), .A3(new_n684), .A4(new_n746), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n747), .A2(KEYINPUT108), .A3(KEYINPUT46), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT108), .B1(new_n747), .B2(KEYINPUT46), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  INV_X1    g550(.A(new_n587), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(G43gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n707), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n741), .A2(new_n742), .A3(new_n697), .A4(new_n729), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G43gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n751), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  AND4_X1   g556(.A1(KEYINPUT110), .A2(new_n682), .A3(new_n746), .A4(new_n753), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n751), .A2(KEYINPUT110), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n707), .B2(new_n753), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n755), .A2(new_n762), .A3(G43gat), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n755), .B2(G43gat), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n757), .B1(new_n761), .B2(new_n765), .ZN(G1330gat));
  INV_X1    g565(.A(new_n208), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n707), .A2(new_n640), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT48), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n741), .A2(new_n742), .A3(new_n640), .A4(new_n729), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n208), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n769), .B1(new_n768), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1331gat));
  NOR2_X1   g573(.A1(new_n740), .A2(new_n328), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n704), .A2(new_n703), .A3(new_n673), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n679), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g579(.A1(new_n777), .A2(new_n683), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(G1333gat));
  OR3_X1    g584(.A1(new_n777), .A2(G71gat), .A3(new_n752), .ZN(new_n786));
  OAI21_X1  g585(.A(G71gat), .B1(new_n777), .B2(new_n639), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1334gat));
  NAND2_X1  g589(.A1(new_n778), .A2(new_n640), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g591(.A1(new_n302), .A2(new_n673), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n328), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n727), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n679), .A2(G85gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n725), .A2(new_n704), .A3(new_n793), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n736), .A2(new_n716), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n737), .A2(new_n739), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n265), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n513), .B(new_n328), .C1(new_n800), .C2(new_n804), .ZN(new_n805));
  OAI221_X1 g604(.A(KEYINPUT111), .B1(new_n796), .B2(new_n797), .C1(new_n805), .C2(G85gat), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n328), .B1(new_n800), .B2(new_n804), .ZN(new_n808));
  AOI21_X1  g607(.A(G85gat), .B1(new_n808), .B2(new_n679), .ZN(new_n809));
  INV_X1    g608(.A(new_n797), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n727), .A2(new_n795), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n812), .ZN(G1336gat));
  NOR2_X1   g612(.A1(new_n683), .A2(G92gat), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n741), .A2(new_n742), .A3(new_n684), .A4(new_n795), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(new_n818), .B2(G92gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n808), .A2(KEYINPUT113), .A3(new_n814), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(G92gat), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n814), .A2(new_n327), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT112), .Z(new_n824));
  AOI21_X1  g623(.A(KEYINPUT51), .B1(new_n803), .B2(new_n793), .ZN(new_n825));
  NOR4_X1   g624(.A1(new_n740), .A2(new_n799), .A3(new_n265), .A4(new_n794), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT52), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n821), .A2(new_n829), .ZN(G1337gat));
  NOR3_X1   g629(.A1(new_n796), .A2(new_n232), .A3(new_n639), .ZN(new_n831));
  AOI21_X1  g630(.A(G99gat), .B1(new_n808), .B2(new_n587), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(G1338gat));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n727), .A2(new_n834), .A3(new_n640), .A4(new_n795), .ZN(new_n835));
  XNOR2_X1  g634(.A(KEYINPUT114), .B(G106gat), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n741), .A2(new_n742), .A3(new_n640), .A4(new_n795), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT115), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n808), .A2(new_n233), .A3(new_n640), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n837), .A2(new_n836), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n233), .B(new_n327), .C1(new_n825), .C2(new_n826), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n581), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(new_n846), .ZN(G1339gat));
  NAND3_X1  g646(.A1(new_n259), .A2(new_n202), .A3(new_n260), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n263), .B1(new_n262), .B2(new_n258), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n652), .A2(new_n850), .A3(new_n654), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n658), .A2(new_n659), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n661), .B2(new_n653), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n668), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n855), .A2(new_n672), .A3(new_n327), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n316), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n314), .A2(new_n305), .A3(new_n315), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT54), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n859), .B(new_n323), .C1(new_n861), .C2(new_n316), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n317), .A2(KEYINPUT54), .A3(new_n860), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n325), .B1(new_n316), .B2(new_n858), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n864), .A2(new_n326), .A3(new_n865), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n671), .B2(new_n672), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n848), .B(new_n849), .C1(new_n856), .C2(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n855), .A2(new_n672), .ZN(new_n872));
  INV_X1    g671(.A(new_n869), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n872), .B(new_n873), .C1(new_n261), .C2(new_n264), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n703), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n329), .A2(new_n673), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n583), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n679), .A3(new_n683), .ZN(new_n883));
  OAI21_X1  g682(.A(G113gat), .B1(new_n883), .B2(new_n728), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n878), .A2(new_n703), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n877), .B1(new_n871), .B2(new_n874), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n881), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n583), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n679), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT119), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n887), .A2(new_n891), .A3(new_n679), .A4(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n683), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n673), .A2(new_n438), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n884), .B1(new_n894), .B2(new_n895), .ZN(G1340gat));
  OAI21_X1  g695(.A(G120gat), .B1(new_n883), .B2(new_n328), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n327), .A2(new_n436), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n894), .B2(new_n898), .ZN(G1341gat));
  AOI21_X1  g698(.A(new_n891), .B1(new_n882), .B2(new_n679), .ZN(new_n900));
  AND4_X1   g699(.A1(new_n891), .A2(new_n887), .A3(new_n679), .A4(new_n888), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n683), .B(new_n302), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(G127gat), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n893), .A2(KEYINPUT120), .A3(new_n683), .A4(new_n302), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n883), .A2(new_n905), .A3(new_n703), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(G1342gat));
  NOR2_X1   g708(.A1(new_n265), .A2(new_n684), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G134gat), .B1(new_n889), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n911), .B(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(G134gat), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n913), .B1(new_n893), .B2(new_n917), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT122), .B(new_n916), .C1(new_n890), .C2(new_n892), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT56), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n900), .B2(new_n901), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT122), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n893), .A2(new_n913), .A3(new_n917), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n912), .B1(new_n920), .B2(new_n925), .ZN(G1343gat));
  AOI21_X1  g725(.A(new_n581), .B1(new_n879), .B2(new_n881), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n697), .A2(new_n513), .A3(new_n684), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n302), .B1(new_n871), .B2(new_n874), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n640), .B1(new_n880), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n933), .B2(KEYINPUT57), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G141gat), .B1(new_n935), .B2(new_n728), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n927), .A2(new_n930), .ZN(new_n937));
  OR3_X1    g736(.A1(new_n937), .A2(G141gat), .A3(new_n728), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g739(.A(G148gat), .ZN(new_n941));
  INV_X1    g740(.A(new_n935), .ZN(new_n942));
  AOI211_X1 g741(.A(KEYINPUT59), .B(new_n941), .C1(new_n942), .C2(new_n327), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n927), .A2(new_n928), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n703), .B1(new_n875), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT123), .B1(new_n871), .B2(new_n874), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n881), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n928), .A3(new_n640), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n945), .A2(new_n327), .A3(new_n930), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n944), .B1(new_n951), .B2(G148gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n327), .A2(new_n941), .ZN(new_n953));
  OAI22_X1  g752(.A1(new_n943), .A2(new_n952), .B1(new_n937), .B2(new_n953), .ZN(G1345gat));
  NAND3_X1  g753(.A1(new_n927), .A2(new_n302), .A3(new_n930), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT124), .ZN(new_n956));
  INV_X1    g755(.A(G155gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n302), .A2(G155gat), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT125), .Z(new_n959));
  AOI22_X1  g758(.A1(new_n956), .A2(new_n957), .B1(new_n942), .B2(new_n959), .ZN(G1346gat));
  OAI21_X1  g759(.A(G162gat), .B1(new_n935), .B2(new_n265), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n915), .A2(G162gat), .A3(new_n513), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n639), .A3(new_n927), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n964), .B(new_n965), .ZN(G1347gat));
  NOR2_X1   g765(.A1(new_n683), .A2(new_n679), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n887), .A2(new_n888), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(new_n673), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n327), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g771(.A1(new_n968), .A2(new_n302), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n350), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n974), .B1(new_n365), .B2(new_n973), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT60), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n975), .B(new_n976), .ZN(G1350gat));
  NAND2_X1  g776(.A1(new_n968), .A2(new_n704), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n978), .A2(new_n979), .A3(new_n351), .ZN(new_n980));
  XOR2_X1   g779(.A(KEYINPUT61), .B(G190gat), .Z(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n978), .B2(new_n981), .ZN(G1351gat));
  NOR3_X1   g781(.A1(new_n697), .A2(new_n679), .A3(new_n683), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n927), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(G197gat), .B1(new_n985), .B2(new_n673), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n945), .A2(new_n950), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n983), .B(KEYINPUT127), .Z(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n728), .A2(new_n665), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(G1352gat));
  NOR3_X1   g790(.A1(new_n984), .A2(G204gat), .A3(new_n328), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT62), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n945), .A2(new_n327), .A3(new_n950), .ZN(new_n994));
  OAI21_X1  g793(.A(G204gat), .B1(new_n994), .B2(new_n988), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(new_n995), .ZN(G1353gat));
  NAND3_X1  g795(.A1(new_n985), .A2(new_n409), .A3(new_n302), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n945), .A2(new_n302), .A3(new_n950), .A4(new_n983), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n998), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n999));
  AOI21_X1  g798(.A(KEYINPUT63), .B1(new_n998), .B2(G211gat), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(G1354gat));
  AOI21_X1  g800(.A(G218gat), .B1(new_n985), .B2(new_n704), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n265), .A2(new_n410), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1002), .B1(new_n989), .B2(new_n1003), .ZN(G1355gat));
endmodule


