//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n626,
    new_n627, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT66), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT66), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  INV_X1    g014(.A(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G120), .Z(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR3_X1   g028(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n454));
  NAND3_X1  g029(.A1(new_n437), .A2(new_n454), .A3(new_n438), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT70), .Z(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT72), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n468), .A2(G137), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT73), .A3(G101), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(KEYINPUT73), .B1(new_n473), .B2(G101), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n471), .A2(new_n478), .A3(KEYINPUT71), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT71), .B1(new_n471), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g055(.A(G125), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n469), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n468), .A2(new_n471), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n469), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND4_X1  g068(.A1(new_n468), .A2(G126), .A3(G2105), .A4(new_n471), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n468), .A2(new_n471), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n470), .A2(G2104), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n471), .A2(new_n478), .A3(KEYINPUT71), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n497), .B1(new_n501), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n518), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n519), .A2(G51), .A3(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT74), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n515), .A2(new_n519), .A3(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT74), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n529), .A2(new_n533), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n513), .A2(new_n514), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI211_X1 g114(.A(KEYINPUT75), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n539), .B1(new_n513), .B2(new_n514), .ZN(new_n542));
  INV_X1    g117(.A(new_n537), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n540), .A2(G651), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n540), .A2(KEYINPUT76), .A3(new_n544), .A4(G651), .ZN(new_n548));
  INV_X1    g123(.A(new_n522), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n515), .A2(new_n519), .ZN(new_n550));
  AOI22_X1  g125(.A1(G52), .A2(new_n549), .B1(new_n550), .B2(G90), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AOI22_X1  g128(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n517), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n515), .A2(new_n519), .A3(G81), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n519), .A2(G43), .A3(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT77), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n555), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT78), .Z(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  XNOR2_X1  g144(.A(KEYINPUT79), .B(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n538), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(new_n550), .B2(G91), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n519), .A2(G53), .A3(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n519), .A2(new_n576), .A3(G53), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n572), .A2(new_n573), .A3(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n573), .B1(new_n572), .B2(new_n578), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n515), .A2(new_n519), .A3(G87), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n519), .A2(G49), .A3(G543), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT81), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G288));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n513), .B2(new_n514), .ZN(new_n594));
  AND2_X1   g169(.A1(G73), .A2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n515), .A2(new_n519), .A3(G86), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n519), .A2(G48), .A3(G543), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n517), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  XOR2_X1   g177(.A(KEYINPUT82), .B(G47), .Z(new_n603));
  OAI22_X1  g178(.A1(new_n520), .A2(new_n602), .B1(new_n522), .B2(new_n603), .ZN(new_n604));
  OR3_X1    g179(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT83), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT83), .B1(new_n601), .B2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  AOI22_X1  g182(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G54), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n608), .A2(new_n517), .B1(new_n609), .B2(new_n522), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n520), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n550), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G171), .B2(new_n617), .ZN(G284));
  XNOR2_X1  g194(.A(G284), .B(KEYINPUT84), .ZN(G321));
  NAND2_X1  g195(.A1(G299), .A2(new_n617), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n617), .B2(G168), .ZN(G297));
  OAI21_X1  g197(.A(new_n621), .B1(new_n617), .B2(G168), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n615), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n615), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n562), .ZN(G323));
  XOR2_X1   g203(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n629));
  XNOR2_X1  g204(.A(G323), .B(new_n629), .ZN(G282));
  NAND2_X1  g205(.A1(new_n507), .A2(new_n473), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT12), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT12), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n507), .A2(new_n633), .A3(new_n473), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n486), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n488), .A2(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(KEYINPUT87), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(KEYINPUT87), .ZN(new_n644));
  OR3_X1    g219(.A1(new_n469), .A2(KEYINPUT86), .A3(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(KEYINPUT86), .B1(new_n469), .B2(G111), .ZN(new_n646));
  NAND4_X1  g221(.A1(new_n643), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n640), .A2(new_n641), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n638), .A2(new_n639), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT88), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2430), .Z(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(G14), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n663), .ZN(G401));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT89), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n669), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n674), .ZN(new_n676));
  OAI21_X1  g251(.A(KEYINPUT17), .B1(new_n672), .B2(new_n673), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n670), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(new_n692), .B(new_n691), .S(new_n684), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  NAND2_X1  g276(.A1(G299), .A2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G20), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT23), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G1956), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G1961), .ZN(new_n709));
  NOR2_X1   g284(.A1(G171), .A2(new_n703), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G5), .B2(new_n703), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G35), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT100), .Z(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G162), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT29), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n708), .B1(new_n709), .B2(new_n711), .C1(G2090), .C2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT99), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n468), .A2(new_n471), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n719), .A2(G141), .A3(new_n469), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n719), .A2(G129), .A3(G2105), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT26), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  AOI22_X1  g300(.A1(G105), .A2(new_n473), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n720), .A2(new_n721), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(new_n712), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n712), .B2(G32), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G160), .A2(G29), .ZN(new_n732));
  AND2_X1   g307(.A1(KEYINPUT24), .A2(G34), .ZN(new_n733));
  NOR2_X1   g308(.A1(KEYINPUT24), .A2(G34), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n712), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT96), .Z(new_n736));
  AOI21_X1  g311(.A(G2084), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n731), .B(new_n737), .C1(new_n709), .C2(new_n711), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n717), .B1(new_n718), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n703), .A2(G4), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n615), .B2(new_n703), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1348), .ZN(new_n742));
  INV_X1    g317(.A(G1341), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n562), .A2(G16), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G16), .B2(G19), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n742), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n712), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n468), .A2(G140), .A3(new_n469), .A4(new_n471), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n468), .A2(G128), .A3(G2105), .A4(new_n471), .ZN(new_n750));
  OR2_X1    g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n751), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(new_n712), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n746), .B(new_n757), .C1(new_n743), .C2(new_n745), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT94), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n738), .A2(new_n718), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n712), .A2(G33), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n507), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(new_n469), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n719), .A2(G139), .A3(new_n469), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT25), .Z(new_n766));
  AND3_X1   g341(.A1(new_n764), .A2(KEYINPUT95), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(KEYINPUT95), .B1(new_n764), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n763), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n761), .B1(new_n769), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2072), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT97), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n716), .A2(G2090), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n770), .A2(new_n771), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n703), .A2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G168), .B2(new_n703), .ZN(new_n778));
  INV_X1    g353(.A(G1966), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G27), .A2(G29), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G164), .B2(G29), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n780), .B1(G2078), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT31), .B(G11), .Z(new_n784));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n712), .B1(new_n785), .B2(G28), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT98), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n787), .A2(KEYINPUT98), .B1(new_n785), .B2(G28), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n648), .B2(new_n712), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n729), .B2(new_n730), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n782), .A2(G2078), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n732), .A2(G2084), .A3(new_n736), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR4_X1   g370(.A1(new_n773), .A2(new_n776), .A3(new_n783), .A4(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n739), .A2(new_n759), .A3(new_n760), .A4(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G24), .B(G290), .S(G16), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1986), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n712), .A2(G25), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n486), .A2(G131), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n488), .A2(G119), .ZN(new_n802));
  OR2_X1    g377(.A1(G95), .A2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n803), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(new_n712), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n807), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n799), .A2(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G6), .B(G305), .S(G16), .Z(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT32), .B(G1981), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT91), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n812), .B(new_n814), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n703), .A2(G22), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G166), .B2(new_n703), .ZN(new_n817));
  INV_X1    g392(.A(G1971), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n703), .A2(G23), .ZN(new_n820));
  INV_X1    g395(.A(new_n587), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n703), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT33), .B(G1976), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n815), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT34), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n811), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n825), .A2(KEYINPUT34), .B1(new_n830), .B2(KEYINPUT36), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n829), .A2(new_n831), .A3(new_n833), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n797), .B1(new_n835), .B2(new_n836), .ZN(G311));
  INV_X1    g412(.A(new_n797), .ZN(new_n838));
  INV_X1    g413(.A(new_n836), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n833), .B1(new_n829), .B2(new_n831), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(G150));
  AOI22_X1  g416(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n517), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  INV_X1    g419(.A(G55), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n520), .A2(new_n844), .B1(new_n522), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n562), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n562), .A2(new_n852), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n848), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n562), .A2(new_n852), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n857), .A2(new_n847), .A3(new_n853), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT38), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n616), .A2(new_n624), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n856), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n861), .B1(new_n860), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n851), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT102), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  AOI21_X1  g443(.A(G860), .B1(new_n868), .B2(KEYINPUT39), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n867), .A2(KEYINPUT103), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT103), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n850), .B1(new_n870), .B2(new_n871), .ZN(G145));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n769), .A2(KEYINPUT105), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n763), .B(new_n875), .C1(new_n767), .C2(new_n768), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(G164), .A2(KEYINPUT104), .ZN(new_n878));
  NAND2_X1  g453(.A1(G164), .A2(KEYINPUT104), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n720), .A2(new_n721), .A3(new_n726), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n754), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n754), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n878), .B(new_n879), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n727), .A2(new_n753), .ZN(new_n885));
  AND2_X1   g460(.A1(G164), .A2(KEYINPUT104), .ZN(new_n886));
  NOR2_X1   g461(.A1(G164), .A2(KEYINPUT104), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n881), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n877), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n874), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n884), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n486), .A2(G142), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n488), .A2(G130), .ZN(new_n895));
  OR2_X1    g470(.A1(G106), .A2(G2105), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n896), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n635), .A2(new_n894), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(new_n632), .A3(new_n634), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n898), .A2(new_n900), .A3(new_n806), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n806), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT106), .B1(new_n893), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  AOI211_X1 g481(.A(new_n906), .B(new_n903), .C1(new_n890), .C2(new_n892), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n873), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n874), .A2(new_n876), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n884), .B2(new_n888), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n891), .A2(new_n884), .A3(new_n888), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n906), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n893), .A2(KEYINPUT106), .A3(new_n904), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(KEYINPUT107), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n893), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n903), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n908), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n492), .B(new_n648), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(G160), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n913), .A2(new_n914), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n916), .B2(new_n903), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n921), .A2(KEYINPUT40), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT40), .B1(new_n921), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(G395));
  XNOR2_X1  g502(.A(new_n626), .B(KEYINPUT108), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n859), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n616), .B1(new_n580), .B2(new_n581), .ZN(new_n930));
  INV_X1    g505(.A(new_n581), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n579), .A3(new_n615), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n935), .A2(KEYINPUT109), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n938));
  NOR2_X1   g513(.A1(G166), .A2(KEYINPUT112), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n518), .A2(new_n524), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(G290), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(G305), .B(new_n587), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n606), .B(new_n605), .C1(new_n939), .C2(new_n942), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n938), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(new_n946), .ZN(new_n950));
  INV_X1    g525(.A(new_n945), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(KEYINPUT113), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n937), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT42), .ZN(new_n956));
  OR3_X1    g531(.A1(new_n955), .A2(KEYINPUT114), .A3(new_n956), .ZN(new_n957));
  XOR2_X1   g532(.A(KEYINPUT111), .B(KEYINPUT41), .Z(new_n958));
  OR2_X1    g533(.A1(new_n933), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n930), .A2(new_n932), .A3(KEYINPUT110), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n616), .B(new_n962), .C1(new_n580), .C2(new_n581), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n935), .A2(KEYINPUT109), .B1(new_n929), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT114), .B1(new_n955), .B2(new_n956), .ZN(new_n967));
  AND4_X1   g542(.A1(new_n936), .A2(new_n957), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n967), .A2(new_n957), .B1(new_n936), .B2(new_n966), .ZN(new_n969));
  OAI21_X1  g544(.A(G868), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n848), .A2(new_n617), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(G295));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n971), .ZN(G331));
  AND2_X1   g548(.A1(new_n949), .A2(new_n954), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n960), .A2(new_n963), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT41), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n533), .A2(new_n534), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n977), .B1(new_n978), .B2(new_n528), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n529), .A2(new_n533), .A3(KEYINPUT115), .A4(new_n534), .ZN(new_n980));
  NAND3_X1  g555(.A1(G301), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  NAND2_X1  g557(.A1(G171), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n856), .A2(new_n858), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n981), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n854), .A2(new_n855), .A3(new_n848), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n847), .B1(new_n857), .B2(new_n853), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n976), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n933), .A3(new_n984), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n933), .A2(new_n958), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n974), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  INV_X1    g569(.A(G37), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n988), .A2(new_n984), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n965), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n949), .A2(new_n954), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n990), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT116), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n964), .A2(new_n959), .B1(new_n988), .B2(new_n984), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n988), .A2(new_n933), .A3(new_n984), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G37), .B1(new_n1004), .B2(new_n998), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n994), .A4(new_n993), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n999), .A2(new_n995), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1004), .A2(new_n998), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT43), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1001), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n994), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1005), .A2(KEYINPUT43), .A3(new_n993), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT44), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(G397));
  INV_X1    g593(.A(G40), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n477), .A2(new_n483), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  INV_X1    g596(.A(G1384), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n507), .A2(new_n508), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(new_n497), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1996), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n727), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT117), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1025), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n754), .A2(new_n756), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n753), .A2(G2067), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n880), .A2(G1996), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1029), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1028), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n805), .A2(new_n809), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n806), .A2(new_n808), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1029), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(G290), .B(G1986), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1029), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT57), .B1(new_n578), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n572), .A2(new_n1045), .A3(new_n578), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n572), .B2(new_n578), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n572), .A2(new_n578), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT122), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n572), .A2(new_n1045), .A3(new_n578), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1043), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1055), .B(new_n1022), .C1(new_n1023), .C2(new_n497), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1020), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n707), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1024), .A2(new_n1021), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT45), .B(new_n1022), .C1(new_n1023), .C2(new_n497), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(new_n1020), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1053), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1058), .A2(new_n1053), .A3(new_n1062), .ZN(new_n1064));
  INV_X1    g639(.A(G1348), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1057), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G125), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n505), .B2(new_n506), .ZN(new_n1068));
  INV_X1    g643(.A(new_n482), .ZN(new_n1069));
  OAI21_X1  g644(.A(G2105), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n473), .A2(G101), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT73), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n474), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1070), .A2(G40), .A3(new_n1074), .A4(new_n472), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n1024), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n756), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n616), .B1(new_n1066), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1063), .B1(new_n1064), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1058), .A2(new_n1053), .A3(new_n1062), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1063), .ZN(new_n1082));
  AOI221_X4 g657(.A(new_n615), .B1(new_n1076), .B2(new_n756), .C1(new_n1057), .C2(new_n1065), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1078), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1053), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1075), .B1(KEYINPUT50), .B2(new_n1024), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1956), .B1(new_n1086), .B2(new_n1056), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1062), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(new_n1064), .A3(KEYINPUT61), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1082), .A2(new_n1084), .A3(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n616), .A2(KEYINPUT60), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1066), .A2(new_n1077), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1059), .A2(new_n1060), .A3(new_n1020), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT123), .B(G1996), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT58), .B(G1341), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n1094), .A2(new_n1095), .B1(new_n1076), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(KEYINPUT59), .A4(new_n562), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1097), .A2(new_n562), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n1101));
  OAI211_X1 g676(.A(new_n1093), .B(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1079), .B1(new_n1091), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1976), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT52), .B1(G288), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1024), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1020), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n821), .A2(G1976), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1105), .A2(new_n1107), .A3(G8), .A4(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(G8), .B(new_n1108), .C1(new_n1075), .C2(new_n1024), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT52), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n1112));
  NAND2_X1  g687(.A1(G305), .A2(G1981), .ZN(new_n1113));
  INV_X1    g688(.A(G1981), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n596), .A2(new_n1114), .A3(new_n597), .A4(new_n598), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT49), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1112), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g693(.A(KEYINPUT118), .B(KEYINPUT49), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1118), .A2(new_n1119), .B1(new_n1117), .B2(new_n1116), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1107), .A2(G8), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1109), .B(new_n1111), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(G303), .A2(G8), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT55), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1054), .A2(new_n1020), .A3(new_n1056), .ZN(new_n1126));
  INV_X1    g701(.A(G2090), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1126), .A2(new_n1127), .B1(new_n1094), .B2(new_n818), .ZN(new_n1128));
  INV_X1    g703(.A(G8), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1125), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1124), .B(KEYINPUT55), .Z(new_n1131));
  AND3_X1   g706(.A1(new_n1059), .A2(new_n1060), .A3(new_n1020), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(G1971), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1057), .A2(G2090), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1131), .B(G8), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1123), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1094), .A2(new_n779), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1137), .B(G168), .C1(G2084), .C2(new_n1057), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(G8), .ZN(new_n1139));
  INV_X1    g714(.A(G2084), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1126), .A2(new_n1140), .B1(new_n1094), .B2(new_n779), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(G168), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT51), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT51), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1138), .A2(new_n1144), .A3(G8), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1136), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G2078), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1132), .A2(KEYINPUT53), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1094), .B2(G2078), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1057), .A2(new_n709), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  OR2_X1    g728(.A1(KEYINPUT125), .A2(G2078), .ZN(new_n1154));
  NAND2_X1  g729(.A1(KEYINPUT125), .A2(G2078), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1149), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1132), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(new_n1150), .A3(G301), .A4(new_n1151), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1152), .A2(G171), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1160), .B1(new_n1162), .B2(G171), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1159), .A2(new_n1160), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1103), .A2(new_n1146), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1135), .A2(new_n1122), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1104), .B(new_n591), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1115), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1168), .A2(KEYINPUT119), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1121), .B1(new_n1168), .B2(KEYINPUT119), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1166), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1141), .A2(new_n1129), .A3(G286), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1172), .A2(new_n1123), .A3(new_n1130), .A4(new_n1135), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1177));
  OAI21_X1  g752(.A(G8), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1122), .B1(new_n1178), .B2(new_n1125), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1179), .A2(KEYINPUT63), .A3(new_n1135), .A4(new_n1172), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1180), .A3(KEYINPUT120), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1165), .A2(new_n1171), .A3(new_n1176), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1184), .B2(KEYINPUT62), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n1186));
  AOI211_X1 g761(.A(KEYINPUT126), .B(new_n1186), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1143), .A2(new_n1186), .A3(new_n1145), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1136), .A2(new_n1153), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1185), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1041), .B1(new_n1182), .B2(new_n1191), .ZN(new_n1192));
  OR3_X1    g767(.A1(new_n1025), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT46), .B1(new_n1025), .B2(G1996), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n727), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1193), .A2(new_n1194), .B1(new_n1029), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1025), .B1(new_n1199), .B2(new_n1030), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1039), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1025), .A2(G1986), .A3(G290), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT48), .Z(new_n1203));
  AOI211_X1 g778(.A(new_n1198), .B(new_n1200), .C1(new_n1201), .C2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1192), .A2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g780(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n700), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g782(.A(new_n1208), .B1(new_n921), .B2(new_n924), .ZN(new_n1209));
  AND2_X1   g783(.A1(new_n1209), .A2(new_n1011), .ZN(G308));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n1011), .ZN(G225));
endmodule


