//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n546,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI211_X1 g035(.A(G137), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n464), .B2(G101), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n458), .A2(G101), .A3(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(KEYINPUT67), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n458), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(new_n460), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT68), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n458), .B1(new_n473), .B2(new_n474), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G124), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n477), .A2(new_n482), .ZN(G162));
  OAI211_X1 g058(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n484));
  OR2_X1    g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n487), .A3(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n459), .B2(new_n460), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n494), .C1(new_n460), .C2(new_n459), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(G164));
  XNOR2_X1  g071(.A(KEYINPUT6), .B(G651), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G50), .ZN(new_n499));
  XNOR2_X1  g074(.A(new_n499), .B(KEYINPUT69), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n497), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n500), .A2(new_n508), .ZN(G303));
  INV_X1    g084(.A(G303), .ZN(G166));
  NAND2_X1  g085(.A1(new_n497), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n497), .A2(KEYINPUT70), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G51), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n503), .A2(new_n497), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT72), .B(G89), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n516), .A2(new_n519), .A3(new_n522), .A4(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  NAND2_X1  g100(.A1(G77), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n502), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n505), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n533), .B1(new_n532), .B2(new_n531), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n515), .A2(G52), .B1(G90), .B2(new_n517), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  NAND2_X1  g112(.A1(new_n515), .A2(G43), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n505), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n538), .B(new_n540), .C1(new_n541), .C2(new_n507), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT74), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND3_X1  g124(.A1(new_n517), .A2(KEYINPUT75), .A3(G91), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n551));
  INV_X1    g126(.A(G91), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n507), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n511), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n497), .A2(new_n557), .A3(G53), .A4(G543), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n529), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n554), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT76), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n550), .A2(new_n553), .B1(G651), .B2(new_n562), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(new_n567), .A3(new_n559), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n517), .A2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n498), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n501), .B2(new_n502), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(KEYINPUT77), .A2(G73), .A3(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n503), .A2(new_n497), .A3(G86), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n497), .A2(G48), .A3(G543), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n515), .A2(G47), .ZN(new_n586));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n529), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(G651), .A2(new_n589), .B1(new_n517), .B2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n515), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n513), .A2(KEYINPUT78), .A3(new_n514), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n594), .A2(G54), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n503), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n505), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n507), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n599), .A2(new_n600), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n592), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n592), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n569), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n569), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n607), .B1(new_n613), .B2(G860), .ZN(G148));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n542), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n606), .A2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g194(.A(KEYINPUT3), .B(G2104), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n464), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT80), .B(G2100), .Z(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n475), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n481), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n458), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND3_X1  g207(.A1(new_n625), .A2(new_n626), .A3(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(KEYINPUT15), .B(G2435), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(new_n637), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n653), .A2(new_n654), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(G2096), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n658), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT84), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G19), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n543), .B2(new_n683), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G1341), .Z(new_n686));
  OR2_X1    g261(.A1(G4), .A2(G16), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n606), .B2(new_n683), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT87), .B(G1348), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n688), .A2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n475), .A2(G140), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n481), .A2(G128), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n458), .A2(G116), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n693), .B(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G29), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G26), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G2067), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n686), .A2(new_n691), .A3(new_n692), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT88), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT91), .B(KEYINPUT23), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n683), .A2(G20), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n569), .B2(new_n683), .ZN(new_n711));
  INV_X1    g286(.A(G1956), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n699), .A2(G35), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G162), .B2(new_n699), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G2090), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT93), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT26), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G129), .B2(new_n481), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n475), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n699), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n699), .B2(G32), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT30), .B(G28), .ZN(new_n731));
  OR2_X1    g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(KEYINPUT31), .A2(G11), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n731), .A2(new_n699), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n631), .B2(new_n699), .ZN(new_n735));
  NAND2_X1  g310(.A1(G164), .A2(G29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G27), .B2(G29), .ZN(new_n737));
  INV_X1    g312(.A(G2078), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR4_X1   g314(.A1(new_n729), .A2(new_n730), .A3(new_n735), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(G160), .A2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n742), .B2(KEYINPUT24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(KEYINPUT24), .B2(new_n742), .ZN(new_n744));
  AOI21_X1  g319(.A(G2084), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n741), .A2(G2084), .A3(new_n744), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n745), .B(new_n746), .C1(new_n738), .C2(new_n737), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n683), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n683), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n740), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n683), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n683), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G1966), .ZN(new_n755));
  NOR2_X1   g330(.A1(G29), .A2(G33), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT89), .Z(new_n757));
  NAND3_X1  g332(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT90), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT25), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n475), .A2(G139), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n620), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n760), .B(new_n761), .C1(new_n458), .C2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n757), .B1(new_n763), .B2(new_n699), .ZN(new_n764));
  INV_X1    g339(.A(G2072), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  AOI22_X1  g342(.A1(G1966), .A2(new_n754), .B1(new_n764), .B2(new_n765), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(new_n716), .C2(G2090), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n752), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n706), .A2(new_n719), .A3(new_n770), .ZN(new_n771));
  MUX2_X1   g346(.A(G6), .B(G305), .S(G16), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  INV_X1    g348(.A(G1981), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n683), .A2(G22), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G166), .B2(new_n683), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(G1971), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n683), .A2(G23), .ZN(new_n779));
  INV_X1    g354(.A(G288), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n683), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT33), .B(G1976), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n777), .B2(G1971), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n775), .A2(new_n778), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n786));
  NOR2_X1   g361(.A1(G16), .A2(G24), .ZN(new_n787));
  XNOR2_X1  g362(.A(G290), .B(KEYINPUT85), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1986), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n475), .A2(G131), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n481), .A2(G119), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n458), .A2(G107), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G25), .B(new_n795), .S(G29), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT35), .B(G1991), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n790), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n786), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT86), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n785), .A2(new_n801), .A3(KEYINPUT34), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n785), .B2(KEYINPUT34), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT36), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n800), .B(new_n806), .C1(new_n803), .C2(new_n802), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n771), .B1(new_n805), .B2(new_n807), .ZN(G311));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n809));
  NOR2_X1   g384(.A1(G311), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g385(.A(KEYINPUT94), .B(new_n771), .C1(new_n805), .C2(new_n807), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(G150));
  AND2_X1   g387(.A1(new_n515), .A2(G55), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n517), .A2(G93), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT95), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n515), .A2(G55), .B1(G93), .B2(new_n517), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n505), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n543), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n819), .A2(new_n543), .A3(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n606), .A2(new_n613), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT96), .B(G860), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n819), .B2(new_n822), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(G145));
  XNOR2_X1  g411(.A(new_n697), .B(KEYINPUT97), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n763), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n795), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n622), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n838), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n724), .B(G164), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n481), .A2(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n458), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G142), .B2(new_n475), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n843), .B(new_n848), .Z(new_n849));
  OR2_X1    g424(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n631), .B(G160), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G162), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n842), .A2(new_n849), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT99), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n852), .B1(new_n850), .B2(new_n853), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(G37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g434(.A(G303), .B(G290), .Z(new_n860));
  XNOR2_X1  g435(.A(G288), .B(G305), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G303), .B(G290), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT42), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n863), .A2(KEYINPUT102), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n867), .A3(KEYINPUT42), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT103), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT103), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n826), .B(new_n617), .Z(new_n876));
  NAND2_X1  g451(.A1(G299), .A2(new_n607), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n569), .A2(new_n606), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n878), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n569), .A2(new_n606), .ZN(new_n882));
  XOR2_X1   g457(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n883));
  NOR3_X1   g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n877), .B2(new_n878), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n876), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n873), .B1(new_n875), .B2(new_n888), .ZN(new_n889));
  NOR4_X1   g464(.A1(new_n874), .A2(KEYINPUT103), .A3(new_n880), .A4(new_n887), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n819), .A2(new_n822), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n615), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(G295));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n893), .ZN(G331));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n897));
  XNOR2_X1  g472(.A(G301), .B(G286), .ZN(new_n898));
  AOI211_X1 g473(.A(new_n821), .B(new_n542), .C1(new_n815), .C2(new_n818), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n823), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT104), .ZN(new_n901));
  INV_X1    g476(.A(new_n898), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n824), .A2(new_n825), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n904), .B(new_n898), .C1(new_n899), .C2(new_n823), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n879), .B2(new_n883), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n907), .B(new_n883), .C1(new_n881), .C2(new_n882), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(new_n879), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n906), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n903), .A2(new_n900), .A3(new_n879), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n866), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n901), .A2(new_n879), .A3(new_n903), .A4(new_n905), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n902), .B1(new_n824), .B2(new_n825), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n899), .A2(new_n823), .A3(new_n898), .ZN(new_n919));
  OAI22_X1  g494(.A1(new_n918), .A2(new_n919), .B1(new_n884), .B2(new_n885), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n920), .A3(new_n866), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n916), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n922), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n866), .B1(new_n917), .B2(new_n920), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n897), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n926), .B1(new_n915), .B2(new_n914), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT106), .B1(new_n930), .B2(new_n924), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n896), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(new_n927), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT43), .B1(new_n923), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT44), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(G397));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G164), .B2(G1384), .ZN(new_n939));
  INV_X1    g514(.A(new_n471), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n464), .A2(new_n462), .A3(G101), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n466), .A2(KEYINPUT67), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(KEYINPUT107), .B(G40), .Z(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n940), .A2(new_n461), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n939), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(KEYINPUT46), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT125), .Z(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(KEYINPUT46), .ZN(new_n953));
  INV_X1    g528(.A(new_n947), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n697), .B(new_n703), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n725), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT126), .Z(new_n957));
  NAND3_X1  g532(.A1(new_n952), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT127), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n724), .B(new_n948), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n963), .A2(new_n955), .ZN(new_n964));
  INV_X1    g539(.A(new_n797), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n795), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n697), .A2(G2067), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n954), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(G290), .A2(G1986), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT48), .B1(new_n970), .B2(new_n947), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n795), .B(new_n797), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n973), .B2(new_n947), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n947), .A3(KEYINPUT48), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n961), .A2(new_n962), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT63), .ZN(new_n978));
  INV_X1    g553(.A(G8), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  INV_X1    g555(.A(new_n495), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n494), .B1(new_n620), .B2(new_n491), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n983), .B2(new_n489), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n946), .B1(new_n984), .B2(KEYINPUT50), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n493), .A2(new_n495), .ZN(new_n986));
  INV_X1    g561(.A(new_n489), .ZN(new_n987));
  AOI21_X1  g562(.A(G1384), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(G2090), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n468), .A2(new_n471), .A3(new_n944), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT45), .B(new_n980), .C1(new_n983), .C2(new_n489), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n939), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1971), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n939), .A2(new_n994), .A3(KEYINPUT109), .A4(new_n993), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n992), .B1(new_n1000), .B2(KEYINPUT110), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n997), .A2(new_n1002), .A3(new_n998), .A4(new_n999), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n979), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT55), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n993), .B1(new_n988), .B2(new_n989), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT116), .B(new_n993), .C1(new_n988), .C2(new_n989), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n990), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1000), .B1(G2090), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT111), .B(G8), .Z(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1006), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n780), .A2(G1976), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n988), .A2(new_n993), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(new_n1016), .ZN(new_n1024));
  AOI211_X1 g599(.A(KEYINPUT112), .B(new_n1015), .C1(new_n988), .C2(new_n993), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1019), .B(new_n1021), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT113), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1016), .B1(new_n984), .B2(new_n946), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT112), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(new_n1022), .A3(new_n1016), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  INV_X1    g610(.A(new_n581), .ZN(new_n1036));
  OAI21_X1  g611(.A(G61), .B1(new_n527), .B2(new_n528), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n505), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n583), .A2(new_n584), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n582), .A2(new_n774), .A3(new_n583), .A4(new_n584), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1040), .A2(new_n1043), .A3(new_n1041), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1048), .A2(KEYINPUT115), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1049), .B2(KEYINPUT49), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1019), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1050), .A2(new_n1031), .B1(new_n1051), .B2(KEYINPUT52), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1034), .A2(new_n1035), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1035), .B1(new_n1034), .B2(new_n1052), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1008), .B(new_n1018), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n985), .A2(new_n1056), .A3(new_n990), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n995), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(G168), .A3(new_n1016), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n978), .B1(new_n1055), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1034), .A2(new_n1052), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1065), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(KEYINPUT118), .C1(new_n1007), .C2(new_n1004), .ZN(new_n1068));
  AOI211_X1 g643(.A(new_n978), .B(new_n1061), .C1(new_n1004), .C2(new_n1007), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1012), .A2(new_n990), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT116), .B1(new_n1074), .B2(new_n993), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n712), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT56), .B(G2072), .Z(new_n1077));
  NOR2_X1   g652(.A1(new_n995), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n564), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n1080));
  OR2_X1    g655(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1081));
  NAND2_X1  g656(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n566), .A2(new_n559), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1076), .A2(new_n1079), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1072), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT122), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1078), .B1(new_n1013), .B2(new_n712), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1072), .B1(new_n1089), .B2(new_n1084), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1080), .A2(new_n1091), .A3(new_n1083), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1089), .B2(KEYINPUT120), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1076), .A2(new_n1079), .A3(KEYINPUT120), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1090), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n988), .A2(new_n993), .A3(new_n703), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n990), .A2(new_n1074), .A3(new_n993), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(G1348), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n607), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n606), .B(new_n1099), .C1(new_n1100), .C2(G1348), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1098), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n939), .A2(new_n994), .A3(new_n948), .A4(new_n993), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT58), .B(G1341), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1023), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1105), .B1(new_n1109), .B2(new_n543), .ZN(new_n1110));
  AOI211_X1 g685(.A(KEYINPUT59), .B(new_n542), .C1(new_n1106), .C2(new_n1108), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n607), .A2(new_n1098), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1110), .A2(new_n1111), .B1(new_n1101), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1104), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(new_n1072), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1088), .A2(new_n1097), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1102), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1085), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n997), .A2(new_n999), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n738), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1961), .B1(new_n985), .B2(new_n990), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1125), .A2(G2078), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n939), .A2(new_n994), .A3(new_n993), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1127), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(KEYINPUT123), .B(new_n1130), .C1(new_n1100), .C2(G1961), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G301), .B1(new_n1126), .B2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n939), .A2(new_n994), .ZN(new_n1136));
  AND3_X1   g711(.A1(G160), .A2(G40), .A3(new_n1129), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n991), .A2(new_n750), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(G2078), .B1(new_n997), .B2(new_n999), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1138), .B(G301), .C1(new_n1139), .C2(KEYINPUT53), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1122), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1126), .A2(new_n1134), .A3(G301), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1138), .B1(new_n1139), .B2(KEYINPUT53), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(G171), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(KEYINPUT54), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1060), .A2(G286), .A3(new_n1016), .ZN(new_n1147));
  NOR2_X1   g722(.A1(G168), .A2(new_n1015), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n979), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1147), .B(KEYINPUT51), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1060), .A2(new_n1016), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(KEYINPUT51), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1142), .A2(new_n1146), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1055), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1121), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1050), .A2(G1976), .A3(G288), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1041), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1031), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1008), .B2(new_n1065), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1150), .A2(KEYINPUT62), .A3(new_n1153), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n1135), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT62), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1161), .B1(new_n1156), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1071), .A2(new_n1157), .A3(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(G290), .B(G1986), .Z(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(new_n954), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(new_n947), .B2(new_n973), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT108), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1167), .A2(KEYINPUT124), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT124), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n977), .B1(new_n1172), .B2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g749(.A(G319), .ZN(new_n1176));
  NOR4_X1   g750(.A1(G229), .A2(new_n1176), .A3(G401), .A4(G227), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n858), .B(new_n1177), .C1(new_n929), .C2(new_n931), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


