//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n461), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n467), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NAND3_X1  g049(.A1(new_n465), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n462), .A2(new_n464), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(new_n467), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT69), .Z(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n461), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n477), .A2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n482), .A2(new_n484), .B1(new_n485), .B2(G136), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n480), .A2(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n467), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(new_n467), .A3(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n477), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n491), .A2(new_n467), .A3(G138), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n494), .A2(KEYINPUT70), .A3(new_n462), .A4(new_n464), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n489), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n477), .A2(new_n467), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G126), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n496), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n497), .B1(new_n496), .B2(new_n502), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n506), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  INV_X1    g096(.A(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n513), .A2(KEYINPUT73), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n513), .A2(G89), .A3(new_n522), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n511), .A2(new_n512), .A3(new_n527), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n520), .A2(G51), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n528), .A2(new_n529), .A3(new_n532), .A4(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND2_X1  g113(.A1(new_n520), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n523), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n513), .A2(G64), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n515), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT74), .B1(new_n541), .B2(new_n544), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n515), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n520), .A2(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n523), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT75), .ZN(G188));
  AOI22_X1  g137(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n515), .ZN(new_n564));
  OAI211_X1 g139(.A(G53), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n523), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G166), .ZN(G303));
  NAND4_X1  g149(.A1(new_n522), .A2(new_n511), .A3(G87), .A4(new_n512), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n511), .A2(new_n512), .ZN(new_n577));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n515), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(G49), .B2(new_n520), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n515), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n520), .A2(G48), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n523), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n520), .A2(G47), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n523), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n513), .A2(G60), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n515), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OR3_X1    g169(.A1(new_n591), .A2(new_n594), .A3(KEYINPUT77), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT77), .B1(new_n591), .B2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  AND3_X1   g172(.A1(new_n513), .A2(G92), .A3(new_n522), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n577), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n520), .A2(G54), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g183(.A(new_n607), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n571), .B2(G868), .ZN(G280));
  XOR2_X1   g186(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g187(.A(new_n606), .ZN(new_n613));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n485), .A2(G2104), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT13), .Z(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(G2100), .ZN(new_n624));
  INV_X1    g199(.A(G111), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n625), .A2(KEYINPUT79), .A3(G2105), .ZN(new_n626));
  AOI21_X1  g201(.A(KEYINPUT79), .B1(new_n625), .B2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n485), .A2(G135), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n479), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n623), .A2(new_n624), .A3(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  AOI21_X1  g231(.A(KEYINPUT18), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT81), .B(KEYINPUT20), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  AND2_X1   g245(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n664), .A2(new_n671), .A3(new_n667), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT83), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1981), .B(G1986), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  XNOR2_X1  g257(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(G29), .B1(new_n684), .B2(G34), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G34), .B2(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(G160), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT89), .Z(new_n689));
  INV_X1    g264(.A(G2084), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT91), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n479), .A2(G129), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n485), .A2(G141), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT26), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n469), .A2(G105), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n693), .A2(new_n694), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G32), .B(new_n698), .S(G29), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT27), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1996), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G4), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n613), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G1348), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(G5), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G171), .B2(new_n702), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(G1961), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n692), .A2(new_n701), .A3(new_n706), .A4(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n687), .A2(G33), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT87), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  NAND2_X1  g289(.A1(G115), .A2(G2104), .ZN(new_n715));
  INV_X1    g290(.A(G127), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n477), .B2(new_n716), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n717), .A2(G2105), .B1(new_n485), .B2(G139), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n711), .B1(new_n719), .B2(G29), .ZN(new_n720));
  INV_X1    g295(.A(G2072), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT31), .B(G11), .Z(new_n724));
  INV_X1    g299(.A(G28), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n726));
  AOI21_X1  g301(.A(G29), .B1(new_n725), .B2(KEYINPUT30), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n723), .B(new_n728), .C1(new_n687), .C2(new_n633), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n687), .A2(G35), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G162), .B2(new_n687), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT29), .Z(new_n732));
  INV_X1    g307(.A(G2090), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n722), .B(new_n729), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n689), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n702), .A2(G19), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n555), .B2(new_n702), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n735), .A2(G2084), .B1(G1341), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n734), .B(new_n738), .C1(G1341), .C2(new_n737), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n702), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n702), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT90), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n687), .A2(G26), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n479), .A2(G128), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n467), .A2(G116), .ZN(new_n748));
  OAI21_X1  g323(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n485), .A2(G140), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(KEYINPUT86), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(KEYINPUT86), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n746), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n708), .A2(G1961), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n744), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n702), .A2(G20), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT23), .Z(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G299), .B2(G16), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1956), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n687), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n687), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G2078), .Z(new_n767));
  OAI211_X1 g342(.A(new_n764), .B(new_n767), .C1(new_n732), .C2(new_n733), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n710), .A2(new_n739), .A3(new_n760), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G23), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n771));
  NAND2_X1  g346(.A1(G288), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n576), .A2(new_n580), .A3(KEYINPUT85), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n770), .B1(new_n775), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT33), .B(G1976), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n776), .B(new_n777), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n702), .A2(G22), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G166), .B2(new_n702), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1971), .ZN(new_n781));
  NOR2_X1   g356(.A1(G6), .A2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G305), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT32), .B(G1981), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OR3_X1    g361(.A1(new_n778), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT34), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n687), .A2(G25), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n479), .A2(G119), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n485), .A2(G131), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n467), .A2(G107), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT84), .Z(new_n797));
  OAI21_X1  g372(.A(new_n791), .B1(new_n797), .B2(new_n687), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G1991), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G16), .A2(G24), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n595), .A2(new_n596), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1986), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n800), .B(new_n805), .C1(new_n787), .C2(KEYINPUT34), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT36), .B1(new_n790), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n790), .A2(new_n806), .A3(KEYINPUT36), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n769), .B1(new_n808), .B2(new_n809), .ZN(G150));
  INV_X1    g385(.A(G150), .ZN(G311));
  NAND2_X1  g386(.A1(new_n613), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n520), .A2(G55), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n814), .B1(new_n523), .B2(new_n815), .C1(new_n816), .C2(new_n515), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n555), .B2(KEYINPUT92), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT93), .B1(new_n555), .B2(KEYINPUT92), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT93), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n820), .B(new_n821), .C1(new_n551), .C2(new_n554), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n818), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n818), .B1(new_n819), .B2(new_n822), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n813), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n828));
  AOI21_X1  g403(.A(G860), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT94), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n817), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(G145));
  XNOR2_X1  g409(.A(new_n633), .B(G160), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G162), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n698), .B(new_n719), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n752), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n496), .A2(new_n502), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT95), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n496), .A2(new_n502), .A3(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n838), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n485), .A2(G142), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(KEYINPUT96), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT96), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G118), .B2(new_n467), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n845), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G130), .B2(new_n479), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n621), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n796), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n844), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n844), .A2(new_n853), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n836), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n836), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(G37), .B1(new_n861), .B2(new_n857), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g439(.A(G868), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n817), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G166), .B(KEYINPUT100), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n775), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n869));
  XNOR2_X1  g444(.A(G166), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n774), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n802), .A2(G305), .ZN(new_n873));
  NAND2_X1  g448(.A1(G290), .A2(new_n783), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n872), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(KEYINPUT101), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(KEYINPUT101), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n606), .A2(KEYINPUT98), .A3(G299), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n571), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(KEYINPUT98), .B1(new_n564), .B2(new_n570), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n883), .A2(new_n599), .A3(new_n605), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n885), .A3(KEYINPUT41), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n885), .A2(new_n881), .A3(KEYINPUT99), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT99), .B1(new_n885), .B2(new_n881), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n826), .B(new_n616), .ZN(new_n895));
  MUX2_X1   g470(.A(new_n891), .B(new_n894), .S(new_n895), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n880), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n866), .B1(new_n897), .B2(new_n865), .ZN(G295));
  OAI21_X1  g473(.A(new_n866), .B1(new_n897), .B2(new_n865), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n819), .A2(new_n822), .ZN(new_n901));
  INV_X1    g476(.A(new_n817), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n551), .A2(new_n554), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n820), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n547), .A2(G168), .A3(new_n548), .ZN(new_n906));
  NAND2_X1  g481(.A1(G171), .A2(G286), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n905), .A2(new_n823), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n906), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n824), .B2(new_n825), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n890), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n872), .A2(new_n875), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n868), .A2(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n908), .A3(KEYINPUT103), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n917));
  INV_X1    g492(.A(new_n909), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n826), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n912), .B(new_n915), .C1(new_n920), .C2(new_n886), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n886), .B1(new_n916), .B2(new_n919), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n876), .B1(new_n922), .B2(new_n911), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n921), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n922), .A2(new_n911), .A3(new_n876), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n916), .A2(new_n891), .A3(new_n919), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n894), .A2(new_n908), .A3(new_n910), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n915), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n927), .A2(new_n930), .A3(G37), .ZN(new_n931));
  OAI211_X1 g506(.A(KEYINPUT44), .B(new_n926), .C1(new_n931), .C2(new_n924), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n921), .A2(new_n925), .A3(new_n923), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n922), .A2(new_n911), .ZN(new_n938));
  AOI21_X1  g513(.A(G37), .B1(new_n938), .B2(new_n915), .ZN(new_n939));
  INV_X1    g514(.A(new_n930), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n924), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n935), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n900), .B1(new_n933), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n924), .B1(new_n939), .B2(new_n923), .ZN(new_n944));
  NOR4_X1   g519(.A1(new_n927), .A2(new_n930), .A3(KEYINPUT43), .A4(G37), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n934), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(KEYINPUT104), .A3(new_n932), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(G397));
  XOR2_X1   g523(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n843), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G40), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n468), .A2(new_n473), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n752), .A2(G2067), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n747), .A2(new_n757), .A3(new_n751), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n698), .B(G1996), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n961), .A2(KEYINPUT107), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(KEYINPUT107), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n962), .A2(new_n797), .A3(new_n799), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n955), .B1(new_n964), .B2(new_n958), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n796), .B(new_n799), .Z(new_n966));
  NAND2_X1  g541(.A1(new_n956), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT125), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n962), .A2(KEYINPUT125), .A3(new_n963), .A4(new_n967), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n956), .A2(new_n804), .A3(new_n802), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT48), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n965), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n977));
  OR3_X1    g552(.A1(new_n955), .A2(new_n977), .A3(G1996), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n956), .B1(new_n698), .B2(new_n959), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n955), .B2(G1996), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT124), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(KEYINPUT124), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n982), .A2(new_n976), .A3(new_n983), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n975), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT126), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n975), .B(KEYINPUT126), .C1(new_n984), .C2(new_n985), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT110), .B(G8), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(G286), .A2(KEYINPUT119), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT119), .B1(G286), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n839), .A2(new_n951), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n954), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n951), .B1(new_n503), .B2(new_n504), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(KEYINPUT50), .B2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n485), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(G40), .C1(new_n467), .C2(new_n466), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n1001), .B2(new_n949), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1002), .A2(new_n690), .B1(new_n1007), .B2(new_n743), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n998), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n743), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n496), .B2(new_n502), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1004), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n839), .A2(KEYINPUT71), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n496), .A2(new_n502), .A3(new_n497), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n690), .B(new_n1014), .C1(new_n1017), .C2(new_n1012), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n996), .B1(new_n1019), .B2(new_n992), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1010), .B1(new_n1020), .B2(KEYINPUT51), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT120), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n1019), .B2(new_n996), .ZN(new_n1023));
  AOI211_X1 g598(.A(KEYINPUT120), .B(new_n995), .C1(new_n1011), .C2(new_n1018), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1014), .B1(new_n1017), .B2(new_n1012), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT116), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(new_n1014), .C1(new_n1017), .C2(new_n1012), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n705), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n999), .A2(new_n1004), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n757), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT115), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1031), .A2(new_n606), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n606), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT60), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1001), .A2(new_n949), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n840), .A2(KEYINPUT45), .A3(new_n951), .A4(new_n842), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT56), .B(G2072), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n954), .A4(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1012), .B(new_n951), .C1(new_n503), .C2(new_n504), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1004), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1956), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n571), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1048), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n564), .B2(new_n570), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1041), .A2(new_n1046), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT61), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1031), .A2(new_n1034), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT58), .B(G1341), .Z(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n999), .B2(new_n1004), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1039), .B(new_n954), .C1(new_n1017), .C2(new_n950), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(G1996), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n555), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1062), .B(new_n555), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT61), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1051), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n564), .A2(new_n570), .A3(new_n1050), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT117), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1049), .A2(new_n1073), .A3(new_n1051), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1069), .B1(new_n1047), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1067), .A2(new_n1068), .B1(new_n1076), .B2(new_n1054), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1037), .A2(new_n1058), .A3(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1047), .A2(new_n1075), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1054), .B1(new_n1036), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1026), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT108), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1061), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1971), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1038), .A2(KEYINPUT108), .A3(new_n1039), .A4(new_n954), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT109), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1083), .A2(KEYINPUT109), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1002), .A2(new_n733), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(G303), .A2(G8), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT55), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(G8), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1086), .B1(G2090), .B2(new_n1044), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n992), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1093), .ZN(new_n1098));
  INV_X1    g673(.A(G1981), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n583), .A2(new_n587), .A3(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n582), .A2(new_n515), .ZN(new_n1101));
  OAI21_X1  g676(.A(G1981), .B1(new_n1101), .B2(new_n586), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(KEYINPUT111), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT111), .ZN(new_n1105));
  NAND3_X1  g680(.A1(G305), .A2(new_n1105), .A3(G1981), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1103), .A2(new_n1106), .A3(KEYINPUT112), .A4(new_n1104), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1032), .A2(new_n991), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(KEYINPUT49), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n772), .A2(G1976), .A3(new_n773), .ZN(new_n1117));
  INV_X1    g692(.A(G1976), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(G288), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1117), .A2(new_n1112), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1112), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(KEYINPUT52), .B2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1095), .A2(new_n1098), .A3(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1125));
  INV_X1    g700(.A(G1961), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1028), .A2(new_n1126), .A3(new_n1030), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n1128));
  OR3_X1    g703(.A1(new_n1007), .A2(new_n1128), .A3(G2078), .ZN(new_n1129));
  AOI21_X1  g704(.A(G2078), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1127), .B(new_n1129), .C1(new_n1130), .C2(KEYINPUT53), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n952), .A2(new_n1128), .A3(G2078), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1039), .A2(new_n954), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1127), .B(new_n1135), .C1(new_n1130), .C2(KEYINPUT53), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1125), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(G301), .B1(new_n1136), .B2(KEYINPUT122), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1128), .B1(new_n1140), .B2(G2078), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(new_n1142), .A3(new_n1127), .A4(new_n1135), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1131), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(G301), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1081), .A2(new_n1124), .A3(new_n1138), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1090), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1009), .B1(new_n1152), .B2(new_n1089), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1150), .B1(new_n1153), .B2(new_n1094), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1008), .A2(G286), .A3(new_n991), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1155), .A2(KEYINPUT63), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1093), .B1(new_n1153), .B2(KEYINPUT113), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1091), .A2(KEYINPUT113), .A3(G8), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1154), .B(new_n1156), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1095), .A2(new_n1098), .A3(new_n1123), .A4(new_n1155), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G288), .A2(G1976), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n1116), .A2(new_n1164), .B1(new_n1099), .B2(new_n783), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1095), .A2(new_n1150), .B1(new_n1165), .B2(new_n1113), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT62), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT120), .B1(new_n1008), .B2(new_n995), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1019), .A2(new_n1022), .A3(new_n996), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n995), .B1(new_n1008), .B2(new_n991), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n997), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1170), .A2(new_n1172), .A3(new_n1173), .A4(new_n1010), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1167), .A2(new_n1132), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1166), .B1(new_n1175), .B2(new_n1124), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1149), .A2(new_n1163), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n956), .A2(G1986), .A3(G290), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n972), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT106), .Z(new_n1180));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n968), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1177), .A2(KEYINPUT123), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT123), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n990), .B1(new_n1182), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g759(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1186));
  OAI211_X1 g760(.A(new_n863), .B(new_n1186), .C1(new_n944), .C2(new_n945), .ZN(G225));
  INV_X1    g761(.A(G225), .ZN(G308));
endmodule


