

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579;

  XOR2_X1 U317 ( .A(n335), .B(n334), .Z(n285) );
  INV_X1 U318 ( .A(KEYINPUT121), .ZN(n408) );
  XNOR2_X1 U319 ( .A(n408), .B(KEYINPUT54), .ZN(n409) );
  XNOR2_X1 U320 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U321 ( .A(n336), .B(n285), .ZN(n337) );
  XNOR2_X1 U322 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U323 ( .A(KEYINPUT91), .B(n461), .Z(n507) );
  XNOR2_X1 U324 ( .A(n449), .B(G176GAT), .ZN(n450) );
  XNOR2_X1 U325 ( .A(n451), .B(n450), .ZN(G1349GAT) );
  XNOR2_X1 U326 ( .A(G120GAT), .B(G148GAT), .ZN(n286) );
  XOR2_X1 U327 ( .A(n286), .B(G57GAT), .Z(n343) );
  XNOR2_X1 U328 ( .A(KEYINPUT90), .B(n343), .ZN(n288) );
  XNOR2_X1 U329 ( .A(G29GAT), .B(G134GAT), .ZN(n309) );
  INV_X1 U330 ( .A(n309), .ZN(n310) );
  XNOR2_X1 U331 ( .A(G85GAT), .B(n310), .ZN(n287) );
  XNOR2_X1 U332 ( .A(n288), .B(n287), .ZN(n294) );
  XOR2_X1 U333 ( .A(G127GAT), .B(KEYINPUT0), .Z(n290) );
  XNOR2_X1 U334 ( .A(G113GAT), .B(KEYINPUT80), .ZN(n289) );
  XNOR2_X1 U335 ( .A(n290), .B(n289), .ZN(n435) );
  XOR2_X1 U336 ( .A(n435), .B(KEYINPUT6), .Z(n292) );
  NAND2_X1 U337 ( .A1(G225GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U339 ( .A(n294), .B(n293), .Z(n303) );
  XOR2_X1 U340 ( .A(KEYINPUT2), .B(G162GAT), .Z(n296) );
  XNOR2_X1 U341 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U343 ( .A(G141GAT), .B(n297), .ZN(n425) );
  INV_X1 U344 ( .A(n425), .ZN(n301) );
  XOR2_X1 U345 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n299) );
  XNOR2_X1 U346 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n461) );
  XOR2_X1 U350 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n305) );
  XNOR2_X1 U351 ( .A(G50GAT), .B(G43GAT), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U353 ( .A(KEYINPUT67), .B(n306), .ZN(n339) );
  INV_X1 U354 ( .A(n339), .ZN(n326) );
  XOR2_X1 U355 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n308) );
  XNOR2_X1 U356 ( .A(G106GAT), .B(G92GAT), .ZN(n307) );
  XOR2_X1 U357 ( .A(n308), .B(n307), .Z(n317) );
  XOR2_X1 U358 ( .A(G36GAT), .B(G190GAT), .Z(n399) );
  NAND2_X1 U359 ( .A1(n399), .A2(n309), .ZN(n313) );
  INV_X1 U360 ( .A(n399), .ZN(n311) );
  NAND2_X1 U361 ( .A1(n311), .A2(n310), .ZN(n312) );
  NAND2_X1 U362 ( .A1(n313), .A2(n312), .ZN(n315) );
  XNOR2_X1 U363 ( .A(G162GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n319) );
  NAND2_X1 U366 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n321) );
  INV_X1 U368 ( .A(KEYINPUT75), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n324) );
  XNOR2_X1 U370 ( .A(G99GAT), .B(G85GAT), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n322), .B(KEYINPUT74), .ZN(n344) );
  XNOR2_X1 U372 ( .A(n344), .B(KEYINPUT11), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n379) );
  BUF_X1 U375 ( .A(n379), .Z(n557) );
  XOR2_X1 U376 ( .A(KEYINPUT68), .B(G1GAT), .Z(n328) );
  XNOR2_X1 U377 ( .A(G22GAT), .B(G15GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n367) );
  XOR2_X1 U379 ( .A(G169GAT), .B(G8GAT), .Z(n403) );
  XOR2_X1 U380 ( .A(n367), .B(n403), .Z(n330) );
  XNOR2_X1 U381 ( .A(G29GAT), .B(G36GAT), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n338) );
  XOR2_X1 U383 ( .A(KEYINPUT29), .B(G113GAT), .Z(n332) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(G197GAT), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n333), .B(KEYINPUT30), .ZN(n336) );
  XOR2_X1 U387 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n335) );
  NAND2_X1 U388 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XOR2_X1 U389 ( .A(n340), .B(n339), .Z(n563) );
  INV_X1 U390 ( .A(n563), .ZN(n553) );
  XOR2_X1 U391 ( .A(G78GAT), .B(G204GAT), .Z(n342) );
  XNOR2_X1 U392 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n342), .B(n341), .ZN(n418) );
  XNOR2_X1 U394 ( .A(n418), .B(n343), .ZN(n356) );
  XOR2_X1 U395 ( .A(n344), .B(KEYINPUT32), .Z(n346) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U398 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n348) );
  XNOR2_X1 U399 ( .A(KEYINPUT72), .B(KEYINPUT31), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U401 ( .A(n350), .B(n349), .Z(n354) );
  XNOR2_X1 U402 ( .A(G176GAT), .B(G92GAT), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n351), .B(G64GAT), .ZN(n398) );
  XNOR2_X1 U404 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n352), .B(KEYINPUT70), .ZN(n366) );
  XNOR2_X1 U406 ( .A(n398), .B(n366), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n383) );
  XNOR2_X1 U409 ( .A(KEYINPUT41), .B(n383), .ZN(n545) );
  NAND2_X1 U410 ( .A1(n553), .A2(n545), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n357), .B(KEYINPUT46), .ZN(n376) );
  XOR2_X1 U412 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n359) );
  XNOR2_X1 U413 ( .A(G8GAT), .B(G64GAT), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n375) );
  XOR2_X1 U415 ( .A(G57GAT), .B(G78GAT), .Z(n361) );
  XNOR2_X1 U416 ( .A(G183GAT), .B(G127GAT), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n363) );
  XOR2_X1 U418 ( .A(G155GAT), .B(G211GAT), .Z(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n371) );
  XNOR2_X1 U420 ( .A(KEYINPUT76), .B(KEYINPUT12), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n364), .B(KEYINPUT14), .ZN(n365) );
  XOR2_X1 U422 ( .A(n365), .B(KEYINPUT15), .Z(n369) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n371), .B(n370), .ZN(n373) );
  NAND2_X1 U426 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U428 ( .A(n375), .B(n374), .Z(n555) );
  INV_X1 U429 ( .A(n555), .ZN(n572) );
  NAND2_X1 U430 ( .A1(n376), .A2(n572), .ZN(n377) );
  NOR2_X1 U431 ( .A1(n557), .A2(n377), .ZN(n378) );
  XNOR2_X1 U432 ( .A(KEYINPUT47), .B(n378), .ZN(n389) );
  XNOR2_X1 U433 ( .A(KEYINPUT36), .B(n379), .ZN(n575) );
  NAND2_X1 U434 ( .A1(n575), .A2(n555), .ZN(n382) );
  XNOR2_X1 U435 ( .A(KEYINPUT110), .B(KEYINPUT45), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n380), .B(KEYINPUT65), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n386) );
  INV_X1 U438 ( .A(n383), .ZN(n384) );
  NOR2_X1 U439 ( .A1(n553), .A2(n384), .ZN(n385) );
  AND2_X1 U440 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n387), .B(KEYINPUT111), .ZN(n388) );
  NAND2_X1 U442 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n390), .B(KEYINPUT48), .ZN(n540) );
  XOR2_X1 U444 ( .A(KEYINPUT18), .B(KEYINPUT84), .Z(n392) );
  XNOR2_X1 U445 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U447 ( .A(KEYINPUT19), .B(n393), .Z(n442) );
  XNOR2_X1 U448 ( .A(G211GAT), .B(KEYINPUT86), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n394), .B(KEYINPUT21), .ZN(n395) );
  XOR2_X1 U450 ( .A(n395), .B(KEYINPUT85), .Z(n397) );
  XNOR2_X1 U451 ( .A(G197GAT), .B(G218GAT), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n422) );
  XNOR2_X1 U453 ( .A(n442), .B(n422), .ZN(n407) );
  XOR2_X1 U454 ( .A(n399), .B(n398), .Z(n401) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U457 ( .A(n402), .B(KEYINPUT92), .Z(n405) );
  XNOR2_X1 U458 ( .A(n403), .B(G204GAT), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n509) );
  NAND2_X1 U461 ( .A1(n540), .A2(n509), .ZN(n410) );
  NOR2_X1 U462 ( .A1(n507), .A2(n411), .ZN(n561) );
  XOR2_X1 U463 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n413) );
  XNOR2_X1 U464 ( .A(G50GAT), .B(KEYINPUT88), .ZN(n412) );
  XNOR2_X1 U465 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U466 ( .A(KEYINPUT89), .B(G148GAT), .Z(n415) );
  XNOR2_X1 U467 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U469 ( .A(n417), .B(n416), .Z(n424) );
  XOR2_X1 U470 ( .A(G22GAT), .B(n418), .Z(n420) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U473 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U474 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U475 ( .A(n426), .B(n425), .ZN(n455) );
  AND2_X1 U476 ( .A1(n561), .A2(n455), .ZN(n428) );
  XNOR2_X1 U477 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n427) );
  XNOR2_X1 U478 ( .A(n428), .B(n427), .ZN(n447) );
  XOR2_X1 U479 ( .A(KEYINPUT64), .B(KEYINPUT81), .Z(n430) );
  XNOR2_X1 U480 ( .A(KEYINPUT20), .B(KEYINPUT82), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U482 ( .A(G190GAT), .B(G15GAT), .Z(n432) );
  XNOR2_X1 U483 ( .A(G169GAT), .B(G43GAT), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n446) );
  XOR2_X1 U486 ( .A(G134GAT), .B(n435), .Z(n437) );
  NAND2_X1 U487 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U489 ( .A(n438), .B(G99GAT), .Z(n444) );
  XOR2_X1 U490 ( .A(G71GAT), .B(G120GAT), .Z(n440) );
  XNOR2_X1 U491 ( .A(KEYINPUT83), .B(G176GAT), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U495 ( .A(n446), .B(n445), .ZN(n522) );
  NOR2_X2 U496 ( .A1(n447), .A2(n522), .ZN(n448) );
  XOR2_X1 U497 ( .A(KEYINPUT123), .B(n448), .Z(n558) );
  XNOR2_X1 U498 ( .A(n545), .B(KEYINPUT100), .ZN(n527) );
  NAND2_X1 U499 ( .A1(n558), .A2(n527), .ZN(n451) );
  XOR2_X1 U500 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n449) );
  XNOR2_X1 U501 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n470) );
  NAND2_X1 U502 ( .A1(n553), .A2(n383), .ZN(n483) );
  XOR2_X1 U503 ( .A(n455), .B(KEYINPUT28), .Z(n516) );
  XNOR2_X1 U504 ( .A(n509), .B(KEYINPUT27), .ZN(n457) );
  NAND2_X1 U505 ( .A1(n507), .A2(n457), .ZN(n542) );
  NOR2_X1 U506 ( .A1(n516), .A2(n542), .ZN(n521) );
  NAND2_X1 U507 ( .A1(n522), .A2(n521), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n452), .B(KEYINPUT93), .ZN(n464) );
  INV_X1 U509 ( .A(n522), .ZN(n513) );
  NAND2_X1 U510 ( .A1(n509), .A2(n513), .ZN(n453) );
  NAND2_X1 U511 ( .A1(n455), .A2(n453), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT25), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n455), .A2(n513), .ZN(n456) );
  XNOR2_X1 U514 ( .A(KEYINPUT26), .B(n456), .ZN(n562) );
  AND2_X1 U515 ( .A1(n562), .A2(n457), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U517 ( .A(KEYINPUT94), .B(n460), .ZN(n462) );
  NOR2_X1 U518 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n479) );
  NOR2_X1 U520 ( .A1(n557), .A2(n572), .ZN(n466) );
  XNOR2_X1 U521 ( .A(KEYINPUT79), .B(KEYINPUT16), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n467) );
  OR2_X1 U523 ( .A1(n479), .A2(n467), .ZN(n493) );
  NOR2_X1 U524 ( .A1(n483), .A2(n493), .ZN(n468) );
  XOR2_X1 U525 ( .A(KEYINPUT95), .B(n468), .Z(n475) );
  NAND2_X1 U526 ( .A1(n507), .A2(n475), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n470), .B(n469), .ZN(G1324GAT) );
  NAND2_X1 U528 ( .A1(n475), .A2(n509), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n473) );
  NAND2_X1 U531 ( .A1(n475), .A2(n513), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U533 ( .A(G15GAT), .B(n474), .ZN(G1326GAT) );
  NAND2_X1 U534 ( .A1(n475), .A2(n516), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n478) );
  XNOR2_X1 U537 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n486) );
  NOR2_X1 U539 ( .A1(n555), .A2(n479), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT97), .B(n480), .Z(n481) );
  NAND2_X1 U541 ( .A1(n481), .A2(n575), .ZN(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT37), .B(n482), .Z(n506) );
  NOR2_X1 U543 ( .A1(n483), .A2(n506), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT38), .ZN(n490) );
  NAND2_X1 U545 ( .A1(n490), .A2(n507), .ZN(n485) );
  XOR2_X1 U546 ( .A(n486), .B(n485), .Z(G1328GAT) );
  NAND2_X1 U547 ( .A1(n490), .A2(n509), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U549 ( .A1(n490), .A2(n513), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n489), .ZN(G1330GAT) );
  NAND2_X1 U552 ( .A1(n490), .A2(n516), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n496) );
  NAND2_X1 U555 ( .A1(n527), .A2(n563), .ZN(n492) );
  XOR2_X1 U556 ( .A(KEYINPUT101), .B(n492), .Z(n505) );
  NOR2_X1 U557 ( .A1(n493), .A2(n505), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(KEYINPUT102), .ZN(n501) );
  NAND2_X1 U559 ( .A1(n507), .A2(n501), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(n497), .ZN(G1332GAT) );
  NAND2_X1 U562 ( .A1(n501), .A2(n509), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(KEYINPUT104), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(n499), .ZN(G1333GAT) );
  NAND2_X1 U565 ( .A1(n501), .A2(n513), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n500), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n503) );
  NAND2_X1 U568 ( .A1(n516), .A2(n501), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U570 ( .A(G78GAT), .B(n504), .Z(G1335GAT) );
  NOR2_X1 U571 ( .A1(n506), .A2(n505), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n517), .A2(n507), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n511) );
  NAND2_X1 U575 ( .A1(n517), .A2(n509), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G92GAT), .B(n512), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n517), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(KEYINPUT108), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G99GAT), .B(n515), .ZN(G1338GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n519) );
  NAND2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  XOR2_X1 U585 ( .A(G113GAT), .B(KEYINPUT113), .Z(n526) );
  NAND2_X1 U586 ( .A1(n540), .A2(n521), .ZN(n523) );
  NOR2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(KEYINPUT112), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n553), .A2(n535), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n529) );
  NAND2_X1 U592 ( .A1(n535), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n531) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT114), .Z(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n533) );
  NAND2_X1 U597 ( .A1(n555), .A2(n535), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U601 ( .A1(n535), .A2(n557), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n539) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT118), .Z(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  XOR2_X1 U605 ( .A(G141GAT), .B(KEYINPUT119), .Z(n544) );
  NAND2_X1 U606 ( .A1(n540), .A2(n562), .ZN(n541) );
  NOR2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n550), .A2(n553), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n547) );
  NAND2_X1 U611 ( .A1(n550), .A2(n545), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n550), .A2(n555), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n557), .A2(n550), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(KEYINPUT120), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G162GAT), .B(n552), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n553), .A2(n558), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  NAND2_X1 U621 ( .A1(n558), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n562), .ZN(n574) );
  NOR2_X1 U627 ( .A1(n563), .A2(n574), .ZN(n568) );
  XOR2_X1 U628 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n565) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(n566), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  NOR2_X1 U633 ( .A1(n383), .A2(n574), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G204GAT), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n574), .ZN(n573) );
  XOR2_X1 U638 ( .A(G211GAT), .B(n573), .Z(G1354GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n578) );
  INV_X1 U640 ( .A(n574), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

