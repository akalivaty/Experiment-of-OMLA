//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT83), .ZN(new_n203));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT26), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT27), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT28), .A4(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT27), .B(G183gat), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n223), .A2(KEYINPUT67), .A3(KEYINPUT28), .A4(new_n219), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT65), .A4(new_n219), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n214), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n233), .A2(new_n212), .B1(new_n234), .B2(KEYINPUT64), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT23), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(G169gat), .B2(G176gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(new_n210), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n233), .A2(new_n212), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n234), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n243), .A2(new_n244), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n205), .B1(new_n232), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G211gat), .A2(G218gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT22), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(G197gat), .A2(G204gat), .ZN(new_n253));
  AND2_X1   g052(.A1(G197gat), .A2(G204gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G211gat), .B(G218gat), .Z(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G211gat), .B(G218gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n252), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n257), .A2(KEYINPUT71), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n214), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n222), .A2(new_n224), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n245), .A2(new_n247), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n241), .B1(new_n236), .B2(new_n235), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n272), .B2(KEYINPUT25), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT29), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n249), .B(new_n266), .C1(new_n274), .C2(new_n205), .ZN(new_n275));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT73), .ZN(new_n277));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n204), .B1(new_n270), .B2(new_n273), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(new_n232), .B2(new_n248), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n204), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n275), .B(new_n279), .C1(new_n283), .C2(new_n266), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT74), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n273), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n205), .B1(new_n287), .B2(new_n281), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n265), .B1(new_n288), .B2(new_n280), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n289), .A2(new_n290), .A3(new_n275), .A4(new_n279), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n285), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n279), .B1(new_n289), .B2(new_n275), .ZN(new_n293));
  INV_X1    g092(.A(new_n284), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(KEYINPUT30), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT40), .ZN(new_n297));
  INV_X1    g096(.A(G141gat), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G162gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G155gat), .ZN(new_n305));
  INV_X1    g104(.A(G155gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G162gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(KEYINPUT75), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G155gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n301), .B1(new_n313), .B2(G162gat), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n300), .A2(new_n305), .A3(new_n307), .A4(new_n302), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317));
  INV_X1    g116(.A(G127gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(G134gat), .ZN(new_n319));
  INV_X1    g118(.A(G134gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(G127gat), .ZN(new_n321));
  OAI22_X1  g120(.A1(new_n317), .A2(KEYINPUT1), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G113gat), .ZN(new_n324));
  INV_X1    g123(.A(G113gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G120gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G127gat), .B(G134gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT4), .B1(new_n316), .B2(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n322), .A2(new_n330), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT75), .B(G155gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT2), .B1(new_n334), .B2(new_n304), .ZN(new_n335));
  AND4_X1   g134(.A1(new_n300), .A2(new_n305), .A3(new_n307), .A4(new_n302), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n335), .A2(new_n336), .B1(new_n303), .B2(new_n308), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n333), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n330), .A3(KEYINPUT76), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n331), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n309), .B(new_n345), .C1(new_n314), .C2(new_n315), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n341), .A2(new_n342), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT39), .ZN(new_n349));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n353));
  XOR2_X1   g152(.A(G1gat), .B(G29gat), .Z(new_n354));
  XNOR2_X1  g153(.A(G57gat), .B(G85gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G57gat), .B(G85gat), .Z(new_n357));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n353), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(new_n359), .A3(new_n353), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(KEYINPUT82), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n364));
  INV_X1    g163(.A(new_n362), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n364), .B1(new_n365), .B2(new_n360), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n344), .A2(new_n342), .A3(new_n316), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n333), .A2(new_n337), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT39), .B1(new_n372), .B2(new_n351), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n350), .B1(new_n340), .B2(new_n347), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n297), .B1(new_n369), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n367), .B1(new_n374), .B2(new_n349), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(KEYINPUT40), .C1(new_n374), .C2(new_n373), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n340), .A2(new_n347), .A3(new_n350), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(new_n351), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT5), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT5), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n340), .A2(new_n347), .A3(new_n382), .A4(new_n350), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n367), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n376), .A2(new_n378), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n203), .B1(new_n296), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n292), .A2(new_n295), .ZN(new_n388));
  INV_X1    g187(.A(new_n386), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(KEYINPUT83), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n391));
  INV_X1    g190(.A(G228gat), .ZN(new_n392));
  INV_X1    g191(.A(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n281), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n257), .B2(new_n260), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n255), .A2(new_n256), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n258), .B1(new_n252), .B2(new_n259), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n281), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT79), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n316), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n346), .A2(new_n281), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n265), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n394), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT29), .B1(new_n257), .B2(new_n260), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n316), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n341), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT80), .B(new_n316), .C1(new_n408), .C2(KEYINPUT3), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n406), .A2(new_n411), .A3(new_n394), .A4(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n391), .B1(new_n407), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G22gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT31), .B(G50gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND3_X1  g218(.A1(new_n415), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n337), .B1(new_n398), .B2(new_n402), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n263), .A2(new_n264), .B1(new_n346), .B2(new_n281), .ZN(new_n422));
  OAI22_X1  g221(.A1(new_n421), .A2(new_n422), .B1(new_n392), .B2(new_n393), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT81), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  INV_X1    g223(.A(new_n419), .ZN(new_n425));
  OAI21_X1  g224(.A(G22gat), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n407), .A2(new_n414), .A3(new_n391), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n420), .B2(new_n426), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n361), .A2(new_n362), .ZN(new_n432));
  AOI211_X1 g231(.A(new_n431), .B(new_n432), .C1(new_n381), .C2(new_n383), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n381), .A2(new_n432), .A3(new_n383), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n434), .A2(new_n431), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n435), .B2(new_n385), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT37), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n279), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n275), .B1(new_n283), .B2(new_n266), .ZN(new_n439));
  INV_X1    g238(.A(new_n279), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n437), .B1(new_n289), .B2(new_n275), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT38), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n285), .A2(new_n291), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT38), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n249), .B(new_n265), .C1(new_n274), .C2(new_n205), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT37), .B(new_n446), .C1(new_n283), .C2(new_n265), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n445), .B(new_n447), .C1(new_n293), .C2(new_n438), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n436), .A2(new_n443), .A3(new_n444), .A4(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n387), .A2(new_n390), .A3(new_n430), .A4(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT78), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n431), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n432), .B1(new_n381), .B2(new_n383), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n433), .ZN(new_n455));
  INV_X1    g254(.A(new_n432), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n384), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(KEYINPUT78), .A3(new_n431), .A4(new_n434), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n420), .A2(new_n426), .ZN(new_n461));
  INV_X1    g260(.A(new_n427), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n296), .A2(new_n459), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G15gat), .B(G43gat), .Z(new_n465));
  XOR2_X1   g264(.A(new_n465), .B(KEYINPUT68), .Z(new_n466));
  XOR2_X1   g265(.A(G71gat), .B(G99gat), .Z(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT69), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n466), .B(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(G227gat), .A2(G233gat), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n331), .B1(new_n232), .B2(new_n248), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n270), .A2(new_n333), .A3(new_n273), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n469), .B1(new_n473), .B2(KEYINPUT33), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT32), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(new_n472), .ZN(new_n478));
  INV_X1    g277(.A(new_n470), .ZN(new_n479));
  AOI221_X4 g278(.A(new_n475), .B1(new_n469), .B2(KEYINPUT33), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n471), .A2(new_n470), .A3(new_n472), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT70), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n482), .A2(new_n483), .A3(new_n481), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n477), .A2(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n478), .A2(new_n479), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(new_n469), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n485), .A2(new_n484), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n476), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n486), .A2(new_n494), .A3(KEYINPUT36), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n464), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n450), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n430), .A2(new_n495), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n296), .A2(new_n459), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT35), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT84), .B(KEYINPUT35), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n388), .A2(new_n436), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(new_n430), .A3(new_n495), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT18), .ZN(new_n510));
  INV_X1    g309(.A(G1gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT16), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n416), .A2(G15gat), .ZN(new_n516));
  INV_X1    g315(.A(G15gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G22gat), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n516), .A2(new_n518), .A3(new_n514), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n512), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n518), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT90), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n513), .A2(new_n514), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n511), .ZN(new_n524));
  NAND2_X1  g323(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT91), .ZN(new_n527));
  INV_X1    g326(.A(G8gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530));
  OR2_X1    g329(.A1(G43gat), .A2(G50gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(G43gat), .A2(G50gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT14), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT14), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(G29gat), .B2(G36gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G36gat), .ZN(new_n540));
  OR2_X1    g339(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n534), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT89), .B(G50gat), .ZN(new_n545));
  INV_X1    g344(.A(G43gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n533), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n536), .A2(new_n538), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n541), .A2(new_n542), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G36gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n544), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n527), .A2(new_n528), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n520), .A2(new_n524), .A3(new_n556), .A4(new_n525), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n529), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI211_X1 g357(.A(KEYINPUT91), .B(G8gat), .C1(new_n520), .C2(new_n524), .ZN(new_n559));
  INV_X1    g358(.A(new_n557), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(KEYINPUT17), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n544), .B(new_n563), .C1(new_n549), .C2(new_n553), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n558), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n510), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n529), .A2(new_n557), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n562), .A3(new_n564), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n571), .A2(KEYINPUT18), .A3(new_n567), .A4(new_n558), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n558), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n567), .B(KEYINPUT13), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n569), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G169gat), .B(G197gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT86), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G113gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT87), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G141gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n579), .B(new_n325), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n582), .B(new_n298), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT12), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n587), .A3(KEYINPUT12), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n592), .A2(new_n569), .A3(new_n572), .A4(new_n576), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n202), .B1(new_n509), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n501), .A2(new_n508), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(KEYINPUT92), .A3(new_n596), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n602));
  INV_X1    g401(.A(G57gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(G64gat), .ZN(new_n604));
  INV_X1    g403(.A(G64gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(G57gat), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n602), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n608), .A2(KEYINPUT93), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(KEYINPUT93), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G71gat), .B(G78gat), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n608), .B(KEYINPUT93), .ZN(new_n614));
  INV_X1    g413(.A(new_n612), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n615), .A3(new_n607), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G127gat), .B(G155gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT20), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n621), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n617), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n570), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n627), .A2(KEYINPUT96), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(KEYINPUT96), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n621), .B(new_n623), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n628), .B2(new_n629), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n631), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n634), .B1(new_n631), .B2(new_n636), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G190gat), .B(G218gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G85gat), .A2(G92gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT7), .ZN(new_n644));
  NAND2_X1  g443(.A1(G99gat), .A2(G106gat), .ZN(new_n645));
  INV_X1    g444(.A(G85gat), .ZN(new_n646));
  INV_X1    g445(.A(G92gat), .ZN(new_n647));
  AOI22_X1  g446(.A1(KEYINPUT8), .A2(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G99gat), .B(G106gat), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n644), .A3(new_n648), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(G232gat), .A2(G233gat), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n555), .A2(new_n655), .B1(KEYINPUT41), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n562), .A2(new_n564), .A3(new_n654), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n642), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n656), .A2(KEYINPUT41), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G134gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n304), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n657), .A2(new_n658), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n641), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n667), .A2(KEYINPUT97), .A3(new_n659), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT97), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n666), .A2(new_n669), .A3(new_n641), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n665), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n659), .A2(KEYINPUT97), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n641), .B2(new_n666), .ZN(new_n673));
  INV_X1    g472(.A(new_n670), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n673), .A2(new_n661), .A3(new_n664), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n617), .A2(new_n654), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT10), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n613), .A2(new_n651), .A3(new_n616), .A4(new_n653), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n625), .A2(new_n655), .A3(KEYINPUT10), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(G230gat), .A2(G233gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n677), .A2(new_n679), .ZN(new_n685));
  INV_X1    g484(.A(new_n683), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G176gat), .B(G204gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n684), .A2(new_n687), .A3(new_n691), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n640), .A2(new_n676), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n601), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n459), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT99), .B(G1gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1324gat));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n697), .A2(new_n296), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n528), .ZN(new_n703));
  OAI211_X1 g502(.A(KEYINPUT100), .B(G8gat), .C1(new_n697), .C2(new_n296), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT16), .B(G8gat), .Z(new_n706));
  AND3_X1   g505(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n702), .B2(new_n706), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n703), .B(new_n704), .C1(new_n707), .C2(new_n708), .ZN(G1325gat));
  INV_X1    g508(.A(new_n498), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT36), .B1(new_n486), .B2(new_n494), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n517), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n495), .A2(new_n517), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n697), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT101), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n718));
  OAI221_X1 g517(.A(new_n718), .B1(new_n697), .B2(new_n715), .C1(new_n713), .C2(new_n517), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1326gat));
  NOR2_X1   g519(.A1(new_n697), .A2(new_n430), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT43), .B(G22gat), .Z(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1327gat));
  INV_X1    g522(.A(new_n695), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n640), .A2(new_n676), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n598), .B2(new_n600), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n454), .A2(new_n455), .A3(new_n458), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n541), .A4(new_n542), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT45), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n449), .A2(new_n430), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n203), .B(new_n386), .C1(new_n292), .C2(new_n295), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT83), .B1(new_n388), .B2(new_n389), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n463), .A2(new_n460), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n727), .B2(new_n388), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n712), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n734), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT102), .B1(new_n450), .B2(new_n500), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n508), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(new_n742), .A3(new_n676), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n599), .B2(new_n676), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n639), .A2(new_n597), .A3(new_n695), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n730), .B1(new_n749), .B2(new_n727), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n746), .A2(new_n730), .A3(new_n727), .A4(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n551), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n729), .B1(new_n750), .B2(new_n752), .ZN(G1328gat));
  NOR2_X1   g552(.A1(new_n296), .A2(G36gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n726), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT104), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n726), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n748), .B2(new_n296), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n746), .A2(KEYINPUT105), .A3(new_n388), .A4(new_n747), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(G36gat), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n758), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n765), .A3(new_n766), .ZN(G1329gat));
  NAND3_X1  g566(.A1(new_n746), .A2(new_n499), .A3(new_n747), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G43gat), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770));
  INV_X1    g569(.A(new_n495), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(G43gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n726), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n769), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n770), .B1(new_n769), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1330gat));
  INV_X1    g575(.A(new_n545), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n749), .A2(new_n735), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n726), .B2(new_n735), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n748), .A2(new_n430), .A3(new_n545), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT48), .B1(new_n783), .B2(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1331gat));
  NOR4_X1   g584(.A1(new_n640), .A2(new_n596), .A3(new_n676), .A4(new_n724), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n741), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n459), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT106), .B(G57gat), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1332gat));
  INV_X1    g589(.A(new_n787), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n296), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT107), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(new_n795), .A3(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1333gat));
  INV_X1    g598(.A(G71gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n787), .B2(new_n771), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n712), .A2(new_n800), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n791), .A2(KEYINPUT108), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT108), .B1(new_n791), .B2(new_n802), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n735), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g607(.A1(new_n640), .A2(new_n597), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n724), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n743), .B2(new_n745), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(new_n727), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n738), .B1(new_n734), .B2(new_n737), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n450), .A2(new_n500), .A3(KEYINPUT102), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n815), .A2(new_n816), .B1(new_n504), .B2(new_n507), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n671), .A2(new_n675), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n809), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n814), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n741), .A2(KEYINPUT51), .A3(new_n819), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n727), .A2(new_n646), .A3(new_n695), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n813), .A2(new_n646), .B1(new_n824), .B2(new_n825), .ZN(G1336gat));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(KEYINPUT109), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n724), .B1(new_n821), .B2(new_n822), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n388), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n647), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n296), .A2(new_n647), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n676), .A2(new_n742), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n815), .A2(new_n816), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n835), .B2(new_n508), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n810), .B(new_n833), .C1(new_n836), .C2(new_n744), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(KEYINPUT52), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n829), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(G92gat), .B1(new_n830), .B2(new_n388), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(new_n828), .A3(new_n839), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n841), .A2(new_n843), .ZN(G1337gat));
  INV_X1    g643(.A(G99gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n812), .A2(new_n499), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(KEYINPUT110), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(KEYINPUT110), .B2(new_n846), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n845), .A3(new_n495), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1338gat));
  OAI211_X1 g649(.A(new_n735), .B(new_n810), .C1(new_n836), .C2(new_n744), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n851), .A2(KEYINPUT111), .A3(G106gat), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT111), .B1(new_n851), .B2(G106gat), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n430), .A2(G106gat), .A3(new_n724), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(KEYINPUT112), .Z(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n821), .B2(new_n822), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT53), .B1(new_n823), .B2(new_n854), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n851), .A2(G106gat), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n859), .A2(KEYINPUT113), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT113), .B1(new_n859), .B2(new_n860), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n857), .A2(new_n858), .B1(new_n861), .B2(new_n862), .ZN(G1339gat));
  AOI21_X1  g662(.A(new_n686), .B1(new_n680), .B2(new_n681), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n691), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n684), .A2(KEYINPUT54), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n682), .A2(new_n683), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT55), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n596), .A2(new_n694), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n574), .B2(new_n575), .ZN(new_n875));
  INV_X1    g674(.A(new_n575), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n573), .A2(new_n558), .A3(KEYINPUT115), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n566), .A2(KEYINPUT114), .A3(new_n568), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT114), .B1(new_n566), .B2(new_n568), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n595), .B(new_n695), .C1(new_n881), .C2(new_n588), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n676), .B1(new_n873), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n595), .B1(new_n881), .B2(new_n588), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n871), .A2(new_n694), .A3(new_n872), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n818), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n640), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n639), .A2(new_n597), .A3(new_n818), .A4(new_n724), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n459), .B(new_n502), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(new_n296), .ZN(new_n890));
  AOI21_X1  g689(.A(G113gat), .B1(new_n890), .B2(new_n596), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n888), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n502), .A2(new_n459), .A3(new_n388), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(new_n325), .A3(new_n597), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n891), .A2(new_n896), .ZN(G1340gat));
  NAND2_X1  g696(.A1(new_n695), .A2(new_n323), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT116), .Z(new_n899));
  NAND2_X1  g698(.A1(new_n890), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G120gat), .B1(new_n895), .B2(new_n724), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1341gat));
  NAND3_X1  g701(.A1(new_n890), .A2(new_n318), .A3(new_n639), .ZN(new_n903));
  OAI21_X1  g702(.A(G127gat), .B1(new_n895), .B2(new_n640), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1342gat));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n320), .A3(new_n296), .A4(new_n676), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n907));
  OAI21_X1  g706(.A(G134gat), .B1(new_n895), .B2(new_n818), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT117), .ZN(G1343gat));
  NAND3_X1  g710(.A1(new_n712), .A2(new_n727), .A3(new_n296), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n430), .B1(new_n887), .B2(new_n888), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT57), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n882), .A2(KEYINPUT118), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n872), .A2(new_n694), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n864), .A2(new_n865), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n918), .B1(new_n682), .B2(new_n683), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT55), .B1(new_n919), .B2(new_n866), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n882), .A2(KEYINPUT118), .B1(new_n921), .B2(new_n596), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n676), .B1(new_n916), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n640), .B1(new_n923), .B2(new_n886), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n430), .B1(new_n924), .B2(new_n888), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n915), .B(new_n596), .C1(new_n925), .C2(new_n914), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G141gat), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n499), .A2(new_n430), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n892), .A2(new_n727), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n596), .A2(new_n298), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n929), .A2(new_n388), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT120), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n935), .B1(new_n926), .B2(G141gat), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n927), .A2(new_n939), .A3(new_n932), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n927), .B2(new_n932), .ZN(new_n942));
  AOI211_X1 g741(.A(KEYINPUT120), .B(new_n931), .C1(new_n926), .C2(G141gat), .ZN(new_n943));
  OAI22_X1  g742(.A1(new_n942), .A2(new_n943), .B1(new_n937), .B2(new_n936), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n941), .A2(new_n944), .ZN(G1344gat));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n388), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(new_n299), .A3(new_n695), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n925), .A2(new_n914), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n913), .A2(new_n914), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n912), .A2(new_n724), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n949), .A2(KEYINPUT121), .A3(new_n950), .A4(new_n952), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n956), .A2(G148gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n948), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n915), .B1(new_n925), .B2(new_n914), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(new_n724), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n960), .A2(KEYINPUT59), .A3(new_n299), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n947), .B1(new_n958), .B2(new_n961), .ZN(G1345gat));
  OAI21_X1  g761(.A(new_n313), .B1(new_n959), .B2(new_n640), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n334), .A3(new_n639), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1346gat));
  OAI21_X1  g764(.A(G162gat), .B1(new_n959), .B2(new_n818), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n296), .A2(new_n304), .A3(new_n676), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n929), .B2(new_n967), .ZN(G1347gat));
  NOR2_X1   g767(.A1(new_n727), .A2(new_n296), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI211_X1 g769(.A(new_n502), .B(new_n970), .C1(new_n887), .C2(new_n888), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(new_n596), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n695), .ZN(new_n974));
  XNOR2_X1  g773(.A(KEYINPUT122), .B(G176gat), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n974), .B(new_n975), .ZN(G1349gat));
  INV_X1    g775(.A(KEYINPUT60), .ZN(new_n977));
  INV_X1    g776(.A(new_n223), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n971), .A2(new_n978), .A3(new_n639), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n971), .A2(new_n639), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(G183gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n977), .B1(new_n981), .B2(KEYINPUT123), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT123), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n983), .B(new_n979), .C1(new_n980), .C2(G183gat), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n982), .A2(KEYINPUT124), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n982), .A2(new_n984), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT124), .B1(new_n981), .B2(new_n977), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(G1350gat));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n676), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n989), .A2(G190gat), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(G190gat), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT125), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n994), .B1(new_n993), .B2(new_n992), .ZN(G1351gat));
  NOR2_X1   g794(.A1(new_n970), .A2(new_n499), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n913), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(G197gat), .B1(new_n997), .B2(new_n596), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n996), .B(KEYINPUT126), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n951), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n596), .A2(G197gat), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(G1352gat));
  INV_X1    g801(.A(G204gat), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n997), .A2(new_n1003), .A3(new_n695), .ZN(new_n1004));
  XOR2_X1   g803(.A(new_n1004), .B(KEYINPUT62), .Z(new_n1005));
  AND2_X1   g804(.A1(new_n1000), .A2(new_n695), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1005), .B1(new_n1006), .B2(new_n1003), .ZN(G1353gat));
  INV_X1    g806(.A(G211gat), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n997), .A2(new_n1008), .A3(new_n639), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n951), .A2(new_n639), .A3(new_n999), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n1010), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1011));
  AOI21_X1  g810(.A(KEYINPUT63), .B1(new_n1010), .B2(G211gat), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(G1354gat));
  INV_X1    g812(.A(G218gat), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n997), .A2(new_n1014), .A3(new_n676), .ZN(new_n1015));
  AND2_X1   g814(.A1(new_n1000), .A2(new_n676), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1015), .B1(new_n1016), .B2(new_n1014), .ZN(G1355gat));
endmodule


