//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(G137), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(new_n197), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n201), .A3(new_n202), .A4(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n190), .A2(new_n193), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n202), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  AND4_X1   g023(.A1(new_n194), .A2(new_n206), .A3(new_n207), .A4(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n189), .A2(new_n192), .A3(KEYINPUT0), .A4(G128), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n189), .A2(new_n192), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT0), .B(G128), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n205), .A2(new_n202), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n204), .B1(new_n217), .B2(new_n197), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n215), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n215), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n200), .A2(new_n220), .A3(new_n202), .A4(new_n205), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n214), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G116), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT2), .B(G113), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n228), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n210), .A2(new_n222), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(G237), .A2(G953), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G210), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT27), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT26), .B(G101), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT30), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n239), .A2(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(KEYINPUT66), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n240), .B(new_n241), .C1(new_n210), .C2(new_n222), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n219), .A2(new_n221), .ZN(new_n243));
  INV_X1    g057(.A(new_n214), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n194), .A2(new_n206), .A3(new_n207), .A4(new_n209), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n245), .A2(KEYINPUT66), .A3(new_n239), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  AOI211_X1 g062(.A(new_n232), .B(new_n238), .C1(new_n248), .C2(new_n231), .ZN(new_n249));
  AOI21_X1  g063(.A(G902), .B1(new_n249), .B2(KEYINPUT31), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT31), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n231), .B1(new_n210), .B2(new_n222), .ZN(new_n253));
  INV_X1    g067(.A(new_n231), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n245), .A2(new_n254), .A3(new_n246), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n232), .A2(KEYINPUT28), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n238), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n248), .A2(new_n231), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n255), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n251), .B(new_n258), .C1(new_n260), .C2(new_n238), .ZN(new_n261));
  INV_X1    g075(.A(G472), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n250), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT32), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n250), .A2(new_n261), .A3(new_n265), .A4(new_n262), .ZN(new_n266));
  INV_X1    g080(.A(G902), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n255), .A2(new_n252), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n253), .A2(new_n255), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n237), .B(new_n268), .C1(new_n269), .C2(new_n252), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n273));
  INV_X1    g087(.A(new_n260), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n271), .B(new_n270), .C1(new_n274), .C2(new_n237), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n264), .A2(new_n266), .B1(new_n278), .B2(G472), .ZN(new_n279));
  INV_X1    g093(.A(G234), .ZN(new_n280));
  OAI21_X1  g094(.A(G217), .B1(new_n280), .B2(G902), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT68), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT16), .ZN(new_n284));
  INV_X1    g098(.A(G140), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(G125), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(G125), .ZN(new_n287));
  INV_X1    g101(.A(G125), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G140), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n286), .B1(new_n290), .B2(new_n284), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(new_n188), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT23), .B1(new_n187), .B2(G119), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT69), .B1(new_n187), .B2(G119), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G119), .B(G128), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT24), .B(G110), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n295), .A2(G110), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  OAI22_X1  g114(.A1(new_n295), .A2(G110), .B1(new_n296), .B2(new_n298), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n291), .A2(new_n188), .ZN(new_n302));
  OR3_X1    g116(.A1(new_n290), .A2(KEYINPUT70), .A3(G146), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT70), .B1(new_n290), .B2(G146), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT22), .B(G137), .ZN(new_n308));
  INV_X1    g122(.A(G221), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n309), .A2(new_n280), .A3(G953), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n308), .B(new_n310), .Z(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n300), .A2(new_n306), .A3(new_n311), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n283), .B1(new_n315), .B2(G902), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n313), .A2(KEYINPUT25), .A3(new_n267), .A4(new_n314), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n282), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n281), .A2(new_n267), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n279), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n264), .A2(new_n266), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n278), .A2(G472), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n321), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT71), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT9), .B(G234), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n309), .B1(new_n333), .B2(new_n267), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT12), .ZN(new_n335));
  INV_X1    g149(.A(new_n243), .ZN(new_n336));
  INV_X1    g150(.A(G107), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT73), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G107), .ZN(new_n340));
  AOI21_X1  g154(.A(G104), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(G104), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G101), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n337), .B2(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n342), .ZN(new_n347));
  INV_X1    g161(.A(G104), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n338), .A3(new_n340), .ZN(new_n350));
  INV_X1    g164(.A(G101), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n344), .A2(KEYINPUT74), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n354), .B(G101), .C1(new_n341), .C2(new_n343), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT75), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n194), .A2(new_n207), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n359), .A3(new_n355), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n358), .B1(new_n353), .B2(new_n355), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n336), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n358), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT10), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(new_n357), .B2(new_n360), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n351), .B1(new_n347), .B2(new_n350), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(new_n368), .ZN(new_n372));
  OAI22_X1  g186(.A1(new_n362), .A2(KEYINPUT10), .B1(new_n372), .B2(new_n214), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n335), .A2(new_n364), .B1(new_n374), .B2(new_n336), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G140), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT72), .ZN(new_n378));
  INV_X1    g192(.A(G953), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n379), .A2(G227), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n378), .B(new_n380), .Z(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n361), .A2(new_n363), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n243), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT12), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n375), .A2(new_n376), .A3(new_n382), .A4(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n353), .A2(new_n359), .A3(new_n355), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n359), .B1(new_n353), .B2(new_n355), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n387), .A2(new_n388), .A3(new_n365), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n335), .B(new_n243), .C1(new_n389), .C2(new_n362), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT10), .B(new_n365), .C1(new_n387), .C2(new_n388), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n362), .A2(KEYINPUT10), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n372), .A2(new_n214), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n336), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n335), .B1(new_n383), .B2(new_n243), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n395), .A2(new_n381), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n243), .B1(new_n367), .B2(new_n373), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT76), .B1(new_n399), .B2(new_n381), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n386), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G469), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(new_n267), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n267), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n399), .A2(new_n381), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n375), .A2(new_n385), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n381), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n404), .B1(new_n407), .B2(G469), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n334), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G237), .ZN(new_n411));
  OAI211_X1 g225(.A(G952), .B(new_n379), .C1(new_n280), .C2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT95), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(G902), .B(G953), .C1(new_n280), .C2(new_n411), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n415), .B(KEYINPUT96), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(G898), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G214), .B1(G237), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT5), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(G113), .C1(KEYINPUT5), .C2(new_n224), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n229), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(new_n387), .B2(new_n388), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n370), .B(new_n231), .C1(new_n371), .C2(new_n368), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G122), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n430), .B(KEYINPUT77), .Z(new_n431));
  AOI21_X1  g245(.A(new_n422), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n433));
  INV_X1    g247(.A(new_n428), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n357), .A2(new_n360), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n426), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n433), .B1(new_n436), .B2(new_n430), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n427), .A2(new_n433), .A3(new_n430), .A4(new_n428), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n432), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n244), .A2(new_n288), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n288), .B2(new_n358), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n379), .A2(G224), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n425), .B1(new_n357), .B2(new_n360), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n422), .B(new_n431), .C1(new_n445), .C2(new_n434), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT79), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT79), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n429), .A2(new_n448), .A3(new_n422), .A4(new_n431), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n443), .A2(KEYINPUT7), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n442), .B(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n427), .A2(new_n430), .A3(new_n428), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT78), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n455), .B2(new_n438), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n430), .B(KEYINPUT8), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n356), .A2(new_n426), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n445), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT80), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n461), .B(new_n457), .C1(new_n445), .C2(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(G902), .B1(new_n456), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n451), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n451), .B2(new_n464), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n420), .B(new_n421), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n233), .A2(G143), .A3(G214), .ZN(new_n471));
  AOI21_X1  g285(.A(G143), .B1(new_n233), .B2(G214), .ZN(new_n472));
  OAI21_X1  g286(.A(G131), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n233), .A2(G214), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n191), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n233), .A2(G143), .A3(G214), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n201), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT86), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n291), .B(G146), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n473), .A2(new_n477), .A3(new_n482), .A4(new_n478), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n476), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT17), .A3(G131), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n480), .A2(new_n481), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT81), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n290), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT81), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(G146), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n305), .ZN(new_n491));
  NAND2_X1  g305(.A1(KEYINPUT18), .A2(G131), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n484), .B(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G113), .B(G122), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT85), .B(G104), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n496), .B(new_n497), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n473), .A2(new_n477), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n488), .A2(KEYINPUT19), .A3(new_n489), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT82), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n504), .A2(KEYINPUT19), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(KEYINPUT19), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n505), .A2(new_n287), .A3(new_n289), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n188), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT83), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT83), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n503), .A2(new_n510), .A3(new_n188), .A4(new_n507), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n302), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n502), .B1(new_n512), .B2(KEYINPUT84), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT84), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n509), .A2(new_n514), .A3(new_n302), .A4(new_n511), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n513), .A2(new_n515), .B1(new_n491), .B2(new_n493), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n501), .B1(new_n516), .B2(new_n498), .ZN(new_n517));
  NOR2_X1   g331(.A1(G475), .A2(G902), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n470), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n495), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n486), .A2(new_n494), .A3(KEYINPUT88), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(KEYINPUT89), .A3(new_n499), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n501), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n498), .B1(new_n495), .B2(new_n520), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT89), .B1(new_n525), .B2(new_n522), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n267), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n469), .A2(new_n519), .B1(new_n527), .B2(G475), .ZN(new_n528));
  XNOR2_X1  g342(.A(G128), .B(G143), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n529), .B(KEYINPUT93), .Z(new_n530));
  OAI21_X1  g344(.A(KEYINPUT13), .B1(new_n191), .B2(G128), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n187), .B2(G143), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n532), .A2(KEYINPUT92), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n187), .A2(G143), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(KEYINPUT13), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n195), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n530), .A2(new_n195), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n225), .A2(G122), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT90), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n225), .A2(G122), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n540), .A2(KEYINPUT91), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT91), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n338), .A2(new_n340), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n540), .A2(new_n541), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n540), .A2(KEYINPUT91), .A3(new_n541), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n538), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n530), .A2(new_n195), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n529), .B(KEYINPUT93), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G134), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n545), .B1(new_n542), .B2(new_n543), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n541), .A2(KEYINPUT14), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n541), .A2(KEYINPUT14), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n540), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n560), .A2(new_n561), .A3(G107), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n560), .B2(G107), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n556), .B(new_n557), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n552), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n333), .A2(G217), .A3(new_n379), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n566), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n552), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G478), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n570), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n512), .A2(KEYINPUT84), .ZN(new_n575));
  INV_X1    g389(.A(new_n502), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n515), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n494), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n500), .B1(new_n578), .B2(new_n499), .ZN(new_n579));
  INV_X1    g393(.A(new_n518), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT87), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n517), .A2(new_n470), .A3(new_n518), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(KEYINPUT20), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n528), .A2(new_n574), .A3(new_n583), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n410), .A2(new_n468), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n331), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  OAI21_X1  g401(.A(new_n421), .B1(new_n466), .B2(new_n467), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(KEYINPUT97), .B(new_n421), .C1(new_n466), .C2(new_n467), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n419), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n250), .A2(new_n261), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n263), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n409), .A2(new_n321), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n528), .A2(new_n583), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n567), .A2(new_n569), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n569), .B2(KEYINPUT98), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n567), .B(new_n569), .C1(KEYINPUT98), .C2(new_n600), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(G478), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n571), .A2(new_n267), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n570), .B2(new_n571), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n598), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n592), .A2(new_n597), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NAND3_X1  g427(.A1(new_n528), .A2(new_n573), .A3(new_n583), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n592), .A2(new_n597), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NOR2_X1   g432(.A1(new_n312), .A2(KEYINPUT36), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n307), .B(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n620), .A2(new_n267), .A3(new_n281), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n318), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n585), .A2(new_n596), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT99), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT37), .B(G110), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  NAND2_X1  g441(.A1(new_n590), .A2(new_n591), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n622), .B1(new_n326), .B2(new_n327), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n409), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT100), .B(G900), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n413), .B1(new_n416), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n633), .A2(KEYINPUT101), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(KEYINPUT101), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n614), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n628), .A2(new_n630), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  NAND2_X1  g454(.A1(new_n519), .A2(new_n469), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n527), .A2(G475), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n583), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n574), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n421), .A3(new_n622), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n645), .A2(KEYINPUT103), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(KEYINPUT103), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n260), .A2(new_n237), .ZN(new_n648));
  AOI21_X1  g462(.A(G902), .B1(new_n269), .B2(new_n238), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n326), .B1(new_n262), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n451), .A2(new_n464), .ZN(new_n654));
  INV_X1    g468(.A(new_n465), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n451), .A2(new_n464), .A3(new_n465), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT38), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n646), .A2(new_n647), .A3(new_n653), .A4(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n636), .B(KEYINPUT39), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n409), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT40), .ZN(new_n664));
  OR3_X1    g478(.A1(new_n660), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n661), .B1(new_n660), .B2(new_n664), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G143), .ZN(G45));
  AOI211_X1 g482(.A(new_n637), .B(new_n607), .C1(new_n528), .C2(new_n583), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n628), .A2(new_n630), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT105), .B(G146), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G48));
  NAND2_X1  g486(.A1(new_n401), .A2(new_n267), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G469), .ZN(new_n674));
  INV_X1    g488(.A(new_n334), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n675), .A3(new_n403), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n329), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n592), .A2(new_n610), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT41), .B(G113), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT106), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n678), .B(new_n680), .ZN(G15));
  NAND3_X1  g495(.A1(new_n592), .A2(new_n615), .A3(new_n677), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  NAND4_X1  g497(.A1(new_n629), .A2(new_n420), .A3(new_n643), .A4(new_n574), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n674), .A2(new_n675), .A3(new_n403), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT97), .B1(new_n658), .B2(new_n421), .ZN(new_n686));
  INV_X1    g500(.A(new_n591), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT107), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n628), .A2(new_n690), .A3(new_n685), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n684), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n223), .ZN(G21));
  XNOR2_X1  g507(.A(KEYINPUT108), .B(G472), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n593), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT109), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n696), .A2(new_n263), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n321), .A2(KEYINPUT110), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n321), .A2(KEYINPUT110), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n695), .A2(KEYINPUT109), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n697), .A2(new_n420), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n676), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n644), .A3(new_n628), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  INV_X1    g520(.A(new_n669), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n697), .A2(new_n623), .A3(new_n702), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI211_X1 g523(.A(KEYINPUT107), .B(new_n676), .C1(new_n590), .C2(new_n591), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n690), .B1(new_n628), .B2(new_n685), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  INV_X1    g527(.A(new_n421), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n466), .A2(new_n467), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n409), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n700), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n279), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n717), .A2(new_n719), .A3(KEYINPUT42), .A4(new_n669), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n323), .A2(new_n669), .A3(new_n409), .A4(new_n715), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n721), .B2(new_n722), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n720), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT112), .B(G131), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G33));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n638), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n716), .A2(new_n329), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND2_X1  g548(.A1(new_n643), .A2(new_n608), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT43), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n643), .A2(new_n737), .A3(new_n608), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n595), .A3(new_n623), .A4(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n715), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n740), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n739), .A2(KEYINPUT116), .A3(new_n740), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(G469), .B1(new_n407), .B2(KEYINPUT45), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n751), .B(new_n405), .C1(new_n406), .C2(new_n381), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n404), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT46), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT114), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n403), .B1(new_n754), .B2(KEYINPUT46), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n334), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n741), .A2(new_n742), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n662), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n749), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n203), .ZN(G39));
  NOR2_X1   g577(.A1(new_n328), .A2(new_n321), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n669), .A3(new_n715), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n759), .A2(KEYINPUT47), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n755), .A2(KEYINPUT114), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n755), .A2(KEYINPUT114), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n757), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n767), .B1(new_n770), .B2(new_n334), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n765), .B1(new_n766), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT117), .B(G140), .Z(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G42));
  NAND2_X1  g588(.A1(new_n674), .A2(new_n403), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n659), .B1(KEYINPUT49), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n653), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n735), .A2(new_n718), .A3(new_n714), .A4(new_n334), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n775), .A2(KEYINPUT49), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT118), .Z(new_n781));
  AND3_X1   g595(.A1(new_n736), .A2(new_n414), .A3(new_n738), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n676), .A2(new_n714), .A3(new_n658), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n719), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT48), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n689), .A2(new_n691), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n696), .A2(new_n263), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n718), .A2(new_n701), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n788), .A3(new_n782), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n379), .A2(G952), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n321), .A2(new_n777), .A3(new_n414), .A4(new_n783), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n791), .B2(new_n610), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n785), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n782), .A2(new_n788), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n659), .A2(new_n421), .A3(new_n676), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n796));
  OR3_X1    g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n796), .B1(new_n794), .B2(new_n795), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n598), .A2(new_n608), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n782), .A2(new_n783), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n787), .A2(new_n622), .A3(new_n701), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n791), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n799), .A2(new_n803), .A3(KEYINPUT51), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n674), .A2(new_n334), .A3(new_n403), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n766), .A2(new_n771), .A3(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n794), .A2(new_n714), .A3(new_n658), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n793), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n799), .A2(new_n803), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n756), .A2(new_n758), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT47), .B1(new_n811), .B2(new_n675), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n770), .A2(new_n767), .A3(new_n334), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT121), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n766), .A2(new_n815), .A3(new_n771), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n816), .A3(new_n805), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n810), .B1(new_n817), .B2(new_n807), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n809), .B1(new_n818), .B2(KEYINPUT51), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n639), .A2(new_n670), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n628), .A2(new_n644), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n636), .B(KEYINPUT119), .Z(new_n823));
  NAND4_X1  g637(.A1(new_n409), .A2(new_n651), .A3(new_n622), .A4(new_n823), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n712), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n468), .B1(new_n609), .B2(new_n614), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n331), .A2(new_n585), .B1(new_n828), .B2(new_n597), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n592), .B(new_n677), .C1(new_n610), .C2(new_n615), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n830), .A3(new_n624), .A4(new_n705), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n692), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n638), .B(KEYINPUT113), .ZN(new_n833));
  INV_X1    g647(.A(new_n732), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n584), .A2(new_n637), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n802), .A2(new_n669), .B1(new_n835), .B2(new_n629), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n833), .A2(new_n834), .B1(new_n716), .B2(new_n836), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n721), .A2(new_n722), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n723), .A3(new_n725), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n839), .B2(new_n720), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n712), .A2(new_n821), .A3(new_n841), .A4(new_n825), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n827), .A2(new_n832), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n835), .A2(new_n629), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n707), .B2(new_n708), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n731), .A2(new_n732), .B1(new_n847), .B2(new_n717), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n727), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n849), .A2(new_n692), .A3(new_n831), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(KEYINPUT53), .A3(new_n827), .A4(new_n842), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n845), .A2(new_n851), .A3(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT54), .B1(new_n845), .B2(new_n851), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n820), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n639), .A2(new_n670), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n786), .B2(new_n709), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n841), .B1(new_n857), .B2(new_n825), .ZN(new_n858));
  INV_X1    g672(.A(new_n842), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT53), .B1(new_n860), .B2(new_n850), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n843), .A2(new_n844), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n855), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n845), .A2(new_n851), .A3(KEYINPUT54), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(KEYINPUT120), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n819), .B1(new_n854), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(G952), .A2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n781), .B1(new_n866), .B2(new_n867), .ZN(G75));
  AOI21_X1  g682(.A(new_n267), .B1(new_n845), .B2(new_n851), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(G210), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n440), .A2(new_n450), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(new_n444), .Z(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(KEYINPUT123), .A2(KEYINPUT56), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n870), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n379), .A2(G952), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G51));
  AND3_X1   g693(.A1(new_n869), .A2(KEYINPUT124), .A3(new_n753), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT124), .B1(new_n869), .B2(new_n753), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n404), .B(KEYINPUT57), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n863), .A2(new_n864), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n401), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n878), .B1(new_n882), .B2(new_n885), .ZN(G54));
  AND2_X1   g700(.A1(KEYINPUT58), .A2(G475), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n869), .A2(new_n517), .A3(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(KEYINPUT125), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(KEYINPUT125), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n869), .A2(new_n887), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n878), .B1(new_n891), .B2(new_n579), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(G60));
  AND2_X1   g707(.A1(new_n602), .A2(new_n603), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n605), .B(KEYINPUT59), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n863), .A2(new_n864), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(G952), .B2(new_n379), .ZN(new_n898));
  INV_X1    g712(.A(new_n895), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n854), .A2(new_n865), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n898), .B1(new_n900), .B2(new_n894), .ZN(G63));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT60), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n845), .B2(new_n851), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT126), .B1(new_n904), .B2(new_n620), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n878), .B1(new_n904), .B2(new_n620), .ZN(new_n907));
  INV_X1    g721(.A(new_n903), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n861), .B2(new_n862), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n315), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n910), .B(new_n907), .C1(new_n905), .C2(KEYINPUT61), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(G66));
  INV_X1    g728(.A(G224), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n418), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n832), .B2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n871), .B1(G898), .B2(new_n379), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G69));
  INV_X1    g733(.A(new_n749), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n759), .A2(new_n662), .A3(new_n760), .ZN(new_n921));
  AOI22_X1  g735(.A1(new_n920), .A2(new_n921), .B1(new_n839), .B2(new_n720), .ZN(new_n922));
  INV_X1    g736(.A(new_n772), .ZN(new_n923));
  INV_X1    g737(.A(new_n822), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n759), .A2(new_n662), .A3(new_n924), .A4(new_n719), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n925), .A2(new_n733), .A3(new_n857), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n379), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n503), .A2(new_n507), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n248), .B(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(G900), .B2(G953), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n379), .B1(G227), .B2(G900), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n331), .B(new_n662), .C1(new_n610), .C2(new_n615), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n716), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n762), .A2(new_n772), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n667), .A2(new_n939), .A3(new_n857), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n665), .A2(new_n666), .A3(new_n857), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n938), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n943), .A2(new_n379), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n933), .B(new_n935), .C1(new_n944), .C2(new_n930), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n930), .B1(new_n943), .B2(new_n379), .ZN(new_n946));
  INV_X1    g760(.A(new_n932), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n927), .B2(new_n379), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n934), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n949), .ZN(G72));
  NAND4_X1  g764(.A1(new_n938), .A2(new_n940), .A3(new_n942), .A4(new_n832), .ZN(new_n951));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  AOI21_X1  g767(.A(new_n648), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n922), .A2(new_n926), .A3(new_n923), .A4(new_n832), .ZN(new_n955));
  AOI211_X1 g769(.A(new_n260), .B(new_n237), .C1(new_n955), .C2(new_n953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n274), .A2(new_n237), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n953), .B1(new_n957), .B2(new_n249), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT127), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n845), .B2(new_n851), .ZN(new_n960));
  NOR4_X1   g774(.A1(new_n954), .A2(new_n956), .A3(new_n878), .A4(new_n960), .ZN(G57));
endmodule


