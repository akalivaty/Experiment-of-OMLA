

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U555 ( .A1(G164), .A2(G1384), .ZN(n775) );
  INV_X1 U556 ( .A(n525), .ZN(n859) );
  BUF_X1 U557 ( .A(n577), .Z(n551) );
  NOR2_X1 U558 ( .A1(n520), .A2(n940), .ZN(n761) );
  NOR2_X2 U559 ( .A1(G2104), .A2(n528), .ZN(n862) );
  INV_X1 U560 ( .A(KEYINPUT97), .ZN(n809) );
  NOR2_X1 U561 ( .A1(n808), .A2(n807), .ZN(n810) );
  AND2_X1 U562 ( .A1(n581), .A2(n580), .ZN(n582) );
  OR2_X1 U563 ( .A1(n770), .A2(n769), .ZN(n519) );
  AND2_X1 U564 ( .A1(KEYINPUT33), .A2(n760), .ZN(n520) );
  AND2_X1 U565 ( .A1(n771), .A2(n519), .ZN(n521) );
  OR2_X1 U566 ( .A1(KEYINPUT33), .A2(n758), .ZN(n522) );
  INV_X1 U567 ( .A(n742), .ZN(n720) );
  INV_X1 U568 ( .A(KEYINPUT29), .ZN(n717) );
  NOR2_X1 U569 ( .A1(n690), .A2(n773), .ZN(n691) );
  NAND2_X1 U570 ( .A1(n691), .A2(n775), .ZN(n742) );
  AND2_X1 U571 ( .A1(n772), .A2(n521), .ZN(n808) );
  NOR2_X2 U572 ( .A1(G651), .A2(G543), .ZN(n647) );
  XNOR2_X1 U573 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n524) );
  NOR2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XNOR2_X1 U575 ( .A(n524), .B(n523), .ZN(n623) );
  NAND2_X1 U576 ( .A1(G138), .A2(n623), .ZN(n527) );
  INV_X1 U577 ( .A(G2105), .ZN(n528) );
  AND2_X1 U578 ( .A1(n528), .A2(G2104), .ZN(n547) );
  INV_X1 U579 ( .A(n547), .ZN(n525) );
  NAND2_X1 U580 ( .A1(G102), .A2(n859), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n527), .A2(n526), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G126), .A2(n862), .ZN(n530) );
  AND2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n863) );
  NAND2_X1 U584 ( .A1(G114), .A2(n863), .ZN(n529) );
  NAND2_X1 U585 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U586 ( .A1(n532), .A2(n531), .ZN(G164) );
  XNOR2_X1 U587 ( .A(G2446), .B(KEYINPUT98), .ZN(n542) );
  XOR2_X1 U588 ( .A(KEYINPUT99), .B(G2427), .Z(n534) );
  XNOR2_X1 U589 ( .A(G2435), .B(G2438), .ZN(n533) );
  XNOR2_X1 U590 ( .A(n534), .B(n533), .ZN(n538) );
  XOR2_X1 U591 ( .A(G2454), .B(G2430), .Z(n536) );
  XNOR2_X1 U592 ( .A(G1348), .B(G1341), .ZN(n535) );
  XNOR2_X1 U593 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U594 ( .A(n538), .B(n537), .Z(n540) );
  XNOR2_X1 U595 ( .A(G2443), .B(G2451), .ZN(n539) );
  XNOR2_X1 U596 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U597 ( .A(n542), .B(n541), .ZN(n543) );
  AND2_X1 U598 ( .A1(n543), .A2(G14), .ZN(G401) );
  NAND2_X1 U599 ( .A1(G137), .A2(n623), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G113), .A2(n863), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U602 ( .A(KEYINPUT66), .B(n546), .ZN(n690) );
  AND2_X1 U603 ( .A1(n862), .A2(G125), .ZN(n687) );
  NOR2_X1 U604 ( .A1(n690), .A2(n687), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G101), .A2(n547), .ZN(n548) );
  XOR2_X1 U606 ( .A(KEYINPUT23), .B(n548), .Z(n686) );
  AND2_X1 U607 ( .A1(n549), .A2(n686), .ZN(G160) );
  INV_X1 U608 ( .A(G651), .ZN(n553) );
  NOR2_X1 U609 ( .A1(G543), .A2(n553), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT1), .B(n550), .Z(n577) );
  NAND2_X1 U611 ( .A1(G64), .A2(n551), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT69), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G90), .A2(n647), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT0), .B(G543), .Z(n557) );
  NOR2_X2 U615 ( .A1(n557), .A2(n553), .ZN(n650) );
  NAND2_X1 U616 ( .A1(G77), .A2(n650), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n556), .B(KEYINPUT9), .ZN(n559) );
  NOR2_X2 U619 ( .A1(G651), .A2(n557), .ZN(n656) );
  NAND2_X1 U620 ( .A1(G52), .A2(n656), .ZN(n558) );
  NAND2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U622 ( .A1(n561), .A2(n560), .ZN(G171) );
  AND2_X1 U623 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  INV_X1 U625 ( .A(G132), .ZN(G219) );
  NAND2_X1 U626 ( .A1(n650), .A2(G75), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G88), .A2(n647), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT77), .B(n562), .Z(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G50), .A2(n656), .ZN(n566) );
  NAND2_X1 U631 ( .A1(G62), .A2(n551), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(G166) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U636 ( .A(G223), .ZN(n827) );
  NAND2_X1 U637 ( .A1(n827), .A2(G567), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U639 ( .A1(G68), .A2(n650), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n647), .A2(G81), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n571), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n574), .B(KEYINPUT13), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G43), .A2(n656), .ZN(n575) );
  AND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n581) );
  INV_X1 U646 ( .A(KEYINPUT14), .ZN(n579) );
  AND2_X1 U647 ( .A1(n577), .A2(G56), .ZN(n578) );
  XNOR2_X1 U648 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X2 U649 ( .A(n582), .B(KEYINPUT72), .ZN(n960) );
  NAND2_X1 U650 ( .A1(G860), .A2(n960), .ZN(G153) );
  XNOR2_X1 U651 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G54), .A2(n656), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G66), .A2(n551), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G92), .A2(n647), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G79), .A2(n650), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n589), .B(KEYINPUT15), .ZN(n703) );
  INV_X1 U661 ( .A(G868), .ZN(n617) );
  NAND2_X1 U662 ( .A1(n703), .A2(n617), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G53), .A2(n656), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G78), .A2(n650), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n647), .A2(G91), .ZN(n594) );
  XOR2_X1 U668 ( .A(KEYINPUT70), .B(n594), .Z(n595) );
  NOR2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n551), .A2(G65), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(G299) );
  NAND2_X1 U672 ( .A1(G51), .A2(n656), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G63), .A2(n551), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U675 ( .A(KEYINPUT6), .B(n601), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n647), .A2(G89), .ZN(n602) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT4), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G76), .A2(n650), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U680 ( .A(n605), .B(KEYINPUT5), .Z(n606) );
  NOR2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U682 ( .A(KEYINPUT7), .B(n608), .Z(n609) );
  XNOR2_X1 U683 ( .A(KEYINPUT74), .B(n609), .ZN(G168) );
  XOR2_X1 U684 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U685 ( .A1(G299), .A2(n617), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G868), .A2(G286), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U688 ( .A(KEYINPUT75), .B(n612), .Z(G297) );
  INV_X1 U689 ( .A(G860), .ZN(n631) );
  NAND2_X1 U690 ( .A1(n631), .A2(G559), .ZN(n613) );
  INV_X1 U691 ( .A(n703), .ZN(n942) );
  NAND2_X1 U692 ( .A1(n613), .A2(n942), .ZN(n614) );
  XNOR2_X1 U693 ( .A(n614), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U694 ( .A1(n942), .A2(G868), .ZN(n615) );
  NOR2_X1 U695 ( .A1(G559), .A2(n615), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n616), .B(KEYINPUT76), .ZN(n619) );
  AND2_X1 U697 ( .A1(n960), .A2(n617), .ZN(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U699 ( .A1(n862), .A2(G123), .ZN(n620) );
  XNOR2_X1 U700 ( .A(n620), .B(KEYINPUT18), .ZN(n622) );
  NAND2_X1 U701 ( .A1(G111), .A2(n863), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n627) );
  BUF_X1 U703 ( .A(n623), .Z(n858) );
  NAND2_X1 U704 ( .A1(G135), .A2(n858), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G99), .A2(n859), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n1009) );
  XNOR2_X1 U708 ( .A(n1009), .B(G2096), .ZN(n629) );
  INV_X1 U709 ( .A(G2100), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(G156) );
  NAND2_X1 U711 ( .A1(G559), .A2(n942), .ZN(n630) );
  XNOR2_X1 U712 ( .A(n630), .B(n960), .ZN(n668) );
  NAND2_X1 U713 ( .A1(n631), .A2(n668), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G55), .A2(n656), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G67), .A2(n551), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G93), .A2(n647), .ZN(n635) );
  NAND2_X1 U718 ( .A1(G80), .A2(n650), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n670) );
  XOR2_X1 U721 ( .A(n638), .B(n670), .Z(G145) );
  NAND2_X1 U722 ( .A1(G47), .A2(n656), .ZN(n640) );
  NAND2_X1 U723 ( .A1(G60), .A2(n551), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U725 ( .A(KEYINPUT68), .B(n641), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G85), .A2(n647), .ZN(n642) );
  XNOR2_X1 U727 ( .A(KEYINPUT67), .B(n642), .ZN(n643) );
  NOR2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n650), .A2(G72), .ZN(n645) );
  NAND2_X1 U730 ( .A1(n646), .A2(n645), .ZN(G290) );
  NAND2_X1 U731 ( .A1(G48), .A2(n656), .ZN(n649) );
  NAND2_X1 U732 ( .A1(G86), .A2(n647), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n650), .A2(G73), .ZN(n651) );
  XOR2_X1 U735 ( .A(KEYINPUT2), .B(n651), .Z(n652) );
  NOR2_X1 U736 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n551), .A2(G61), .ZN(n654) );
  NAND2_X1 U738 ( .A1(n655), .A2(n654), .ZN(G305) );
  NAND2_X1 U739 ( .A1(G49), .A2(n656), .ZN(n658) );
  NAND2_X1 U740 ( .A1(G74), .A2(G651), .ZN(n657) );
  NAND2_X1 U741 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U742 ( .A1(n551), .A2(n659), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n557), .A2(G87), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n661), .A2(n660), .ZN(G288) );
  XNOR2_X1 U745 ( .A(n670), .B(G290), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n662), .B(G305), .ZN(n663) );
  XNOR2_X1 U747 ( .A(KEYINPUT78), .B(n663), .ZN(n665) );
  XNOR2_X1 U748 ( .A(G288), .B(KEYINPUT19), .ZN(n664) );
  XNOR2_X1 U749 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U750 ( .A(G166), .B(n666), .ZN(n667) );
  XNOR2_X1 U751 ( .A(n667), .B(G299), .ZN(n882) );
  XNOR2_X1 U752 ( .A(n668), .B(n882), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n669), .A2(G868), .ZN(n672) );
  OR2_X1 U754 ( .A1(n670), .A2(G868), .ZN(n671) );
  NAND2_X1 U755 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2084), .A2(G2078), .ZN(n673) );
  XNOR2_X1 U757 ( .A(n673), .B(KEYINPUT20), .ZN(n674) );
  XNOR2_X1 U758 ( .A(n674), .B(KEYINPUT79), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n675), .A2(G2090), .ZN(n676) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U763 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U764 ( .A1(G219), .A2(G220), .ZN(n678) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n678), .Z(n679) );
  NOR2_X1 U766 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U767 ( .A1(G96), .A2(n680), .ZN(n834) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n834), .ZN(n684) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n681) );
  NOR2_X1 U770 ( .A1(G237), .A2(n681), .ZN(n682) );
  NAND2_X1 U771 ( .A1(G108), .A2(n682), .ZN(n835) );
  NAND2_X1 U772 ( .A1(G567), .A2(n835), .ZN(n683) );
  NAND2_X1 U773 ( .A1(n684), .A2(n683), .ZN(n886) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n685) );
  NOR2_X1 U775 ( .A1(n886), .A2(n685), .ZN(n831) );
  NAND2_X1 U776 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  AND2_X1 U778 ( .A1(n686), .A2(G40), .ZN(n689) );
  INV_X1 U779 ( .A(n687), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n773) );
  NAND2_X1 U781 ( .A1(G8), .A2(n742), .ZN(n770) );
  NOR2_X1 U782 ( .A1(G1966), .A2(n770), .ZN(n738) );
  NOR2_X1 U783 ( .A1(G2084), .A2(n742), .ZN(n725) );
  NAND2_X1 U784 ( .A1(n725), .A2(G8), .ZN(n736) );
  NAND2_X1 U785 ( .A1(G1996), .A2(n720), .ZN(n692) );
  XNOR2_X1 U786 ( .A(n692), .B(KEYINPUT26), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n693), .A2(n960), .ZN(n696) );
  NAND2_X1 U788 ( .A1(G1341), .A2(n742), .ZN(n694) );
  XNOR2_X1 U789 ( .A(KEYINPUT89), .B(n694), .ZN(n695) );
  NOR2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n698) );
  INV_X1 U791 ( .A(KEYINPUT64), .ZN(n697) );
  XNOR2_X1 U792 ( .A(n698), .B(n697), .ZN(n704) );
  OR2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n702) );
  NOR2_X1 U794 ( .A1(n720), .A2(G1348), .ZN(n700) );
  NOR2_X1 U795 ( .A1(G2067), .A2(n742), .ZN(n699) );
  NOR2_X1 U796 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n720), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U801 ( .A(n707), .B(KEYINPUT27), .ZN(n709) );
  INV_X1 U802 ( .A(G1956), .ZN(n946) );
  NOR2_X1 U803 ( .A1(n946), .A2(n720), .ZN(n708) );
  NOR2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n712) );
  INV_X1 U805 ( .A(G299), .ZN(n947) );
  NAND2_X1 U806 ( .A1(n712), .A2(n947), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n716) );
  NOR2_X1 U808 ( .A1(n712), .A2(n947), .ZN(n714) );
  XOR2_X1 U809 ( .A(KEYINPUT88), .B(KEYINPUT28), .Z(n713) );
  XNOR2_X1 U810 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U812 ( .A(n718), .B(n717), .ZN(n724) );
  XOR2_X1 U813 ( .A(G2078), .B(KEYINPUT25), .Z(n719) );
  XNOR2_X1 U814 ( .A(KEYINPUT87), .B(n719), .ZN(n917) );
  NOR2_X1 U815 ( .A1(n742), .A2(n917), .ZN(n722) );
  INV_X1 U816 ( .A(G1961), .ZN(n967) );
  NOR2_X1 U817 ( .A1(n720), .A2(n967), .ZN(n721) );
  NOR2_X1 U818 ( .A1(n722), .A2(n721), .ZN(n729) );
  NAND2_X1 U819 ( .A1(G171), .A2(n729), .ZN(n723) );
  NAND2_X1 U820 ( .A1(n724), .A2(n723), .ZN(n734) );
  NOR2_X1 U821 ( .A1(n738), .A2(n725), .ZN(n726) );
  NAND2_X1 U822 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U824 ( .A1(G168), .A2(n728), .ZN(n731) );
  NOR2_X1 U825 ( .A1(G171), .A2(n729), .ZN(n730) );
  NOR2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U827 ( .A(KEYINPUT31), .B(n732), .Z(n733) );
  NAND2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n740) );
  XNOR2_X1 U829 ( .A(n740), .B(KEYINPUT90), .ZN(n735) );
  NAND2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U832 ( .A(n739), .B(KEYINPUT91), .ZN(n752) );
  NAND2_X1 U833 ( .A1(n740), .A2(G286), .ZN(n741) );
  XNOR2_X1 U834 ( .A(n741), .B(KEYINPUT92), .ZN(n748) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n742), .ZN(n743) );
  XNOR2_X1 U836 ( .A(KEYINPUT93), .B(n743), .ZN(n746) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n770), .ZN(n744) );
  NOR2_X1 U838 ( .A1(G166), .A2(n744), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U840 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U841 ( .A1(n749), .A2(G8), .ZN(n750) );
  XNOR2_X1 U842 ( .A(n750), .B(KEYINPUT32), .ZN(n751) );
  NAND2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n764) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n949) );
  XNOR2_X1 U845 ( .A(n949), .B(KEYINPUT95), .ZN(n754) );
  NOR2_X1 U846 ( .A1(G288), .A2(G1976), .ZN(n753) );
  XNOR2_X1 U847 ( .A(n753), .B(KEYINPUT94), .ZN(n953) );
  INV_X1 U848 ( .A(n953), .ZN(n759) );
  AND2_X1 U849 ( .A1(n754), .A2(n759), .ZN(n755) );
  NAND2_X1 U850 ( .A1(n764), .A2(n755), .ZN(n756) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n951) );
  NAND2_X1 U852 ( .A1(n756), .A2(n951), .ZN(n757) );
  NOR2_X1 U853 ( .A1(n770), .A2(n757), .ZN(n758) );
  NOR2_X1 U854 ( .A1(n770), .A2(n759), .ZN(n760) );
  XNOR2_X1 U855 ( .A(G1981), .B(G305), .ZN(n940) );
  NAND2_X1 U856 ( .A1(n522), .A2(n761), .ZN(n772) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U858 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U860 ( .A(n765), .B(KEYINPUT96), .ZN(n766) );
  NAND2_X1 U861 ( .A1(n766), .A2(n770), .ZN(n771) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U863 ( .A(n767), .B(KEYINPUT86), .Z(n768) );
  XNOR2_X1 U864 ( .A(KEYINPUT24), .B(n768), .ZN(n769) );
  OR2_X1 U865 ( .A1(n773), .A2(n690), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n822) );
  XNOR2_X1 U867 ( .A(G2067), .B(KEYINPUT37), .ZN(n776) );
  XNOR2_X1 U868 ( .A(n776), .B(KEYINPUT80), .ZN(n820) );
  NAND2_X1 U869 ( .A1(G140), .A2(n858), .ZN(n778) );
  NAND2_X1 U870 ( .A1(G104), .A2(n859), .ZN(n777) );
  NAND2_X1 U871 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U872 ( .A(KEYINPUT34), .B(n779), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G128), .A2(n862), .ZN(n781) );
  NAND2_X1 U874 ( .A1(G116), .A2(n863), .ZN(n780) );
  NAND2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U876 ( .A(KEYINPUT35), .B(n782), .ZN(n783) );
  XNOR2_X1 U877 ( .A(KEYINPUT81), .B(n783), .ZN(n784) );
  NOR2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U879 ( .A(KEYINPUT36), .B(n786), .ZN(n875) );
  NOR2_X1 U880 ( .A1(n820), .A2(n875), .ZN(n999) );
  NAND2_X1 U881 ( .A1(n822), .A2(n999), .ZN(n818) );
  XNOR2_X1 U882 ( .A(KEYINPUT84), .B(G1991), .ZN(n919) );
  NAND2_X1 U883 ( .A1(G119), .A2(n862), .ZN(n788) );
  NAND2_X1 U884 ( .A1(G107), .A2(n863), .ZN(n787) );
  NAND2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n858), .A2(G131), .ZN(n789) );
  XNOR2_X1 U887 ( .A(n789), .B(KEYINPUT82), .ZN(n791) );
  NAND2_X1 U888 ( .A1(G95), .A2(n859), .ZN(n790) );
  NAND2_X1 U889 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U890 ( .A(KEYINPUT83), .B(n792), .Z(n793) );
  OR2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n869) );
  AND2_X1 U892 ( .A1(n919), .A2(n869), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G105), .A2(n859), .ZN(n795) );
  XNOR2_X1 U894 ( .A(n795), .B(KEYINPUT38), .ZN(n802) );
  NAND2_X1 U895 ( .A1(G129), .A2(n862), .ZN(n797) );
  NAND2_X1 U896 ( .A1(G117), .A2(n863), .ZN(n796) );
  NAND2_X1 U897 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U898 ( .A1(G141), .A2(n858), .ZN(n798) );
  XNOR2_X1 U899 ( .A(KEYINPUT85), .B(n798), .ZN(n799) );
  NOR2_X1 U900 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U901 ( .A1(n802), .A2(n801), .ZN(n874) );
  AND2_X1 U902 ( .A1(n874), .A2(G1996), .ZN(n803) );
  NOR2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n1013) );
  INV_X1 U904 ( .A(n822), .ZN(n805) );
  NOR2_X1 U905 ( .A1(n1013), .A2(n805), .ZN(n815) );
  INV_X1 U906 ( .A(n815), .ZN(n806) );
  NAND2_X1 U907 ( .A1(n818), .A2(n806), .ZN(n807) );
  XNOR2_X1 U908 ( .A(n810), .B(n809), .ZN(n812) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n957) );
  NAND2_X1 U910 ( .A1(n957), .A2(n822), .ZN(n811) );
  NAND2_X1 U911 ( .A1(n812), .A2(n811), .ZN(n825) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n874), .ZN(n1001) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U914 ( .A1(n919), .A2(n869), .ZN(n1010) );
  NOR2_X1 U915 ( .A1(n813), .A2(n1010), .ZN(n814) );
  NOR2_X1 U916 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U917 ( .A1(n1001), .A2(n816), .ZN(n817) );
  XNOR2_X1 U918 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U919 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U920 ( .A1(n820), .A2(n875), .ZN(n1003) );
  NAND2_X1 U921 ( .A1(n821), .A2(n1003), .ZN(n823) );
  NAND2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U923 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n827), .ZN(G217) );
  NAND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n828) );
  XOR2_X1 U927 ( .A(KEYINPUT100), .B(n828), .Z(n829) );
  NAND2_X1 U928 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n830) );
  XOR2_X1 U930 ( .A(KEYINPUT101), .B(n830), .Z(n832) );
  NAND2_X1 U931 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n833), .B(KEYINPUT102), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  NAND2_X1 U939 ( .A1(G124), .A2(n862), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n836), .B(KEYINPUT44), .ZN(n839) );
  NAND2_X1 U941 ( .A1(G136), .A2(n858), .ZN(n837) );
  XOR2_X1 U942 ( .A(KEYINPUT105), .B(n837), .Z(n838) );
  NAND2_X1 U943 ( .A1(n839), .A2(n838), .ZN(n843) );
  NAND2_X1 U944 ( .A1(G100), .A2(n859), .ZN(n841) );
  NAND2_X1 U945 ( .A1(G112), .A2(n863), .ZN(n840) );
  NAND2_X1 U946 ( .A1(n841), .A2(n840), .ZN(n842) );
  NOR2_X1 U947 ( .A1(n843), .A2(n842), .ZN(G162) );
  XOR2_X1 U948 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n845) );
  XNOR2_X1 U949 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n844) );
  XNOR2_X1 U950 ( .A(n845), .B(n844), .ZN(n855) );
  NAND2_X1 U951 ( .A1(G130), .A2(n862), .ZN(n847) );
  NAND2_X1 U952 ( .A1(G118), .A2(n863), .ZN(n846) );
  NAND2_X1 U953 ( .A1(n847), .A2(n846), .ZN(n853) );
  NAND2_X1 U954 ( .A1(G142), .A2(n858), .ZN(n849) );
  NAND2_X1 U955 ( .A1(G106), .A2(n859), .ZN(n848) );
  NAND2_X1 U956 ( .A1(n849), .A2(n848), .ZN(n850) );
  XOR2_X1 U957 ( .A(KEYINPUT45), .B(n850), .Z(n851) );
  XNOR2_X1 U958 ( .A(KEYINPUT106), .B(n851), .ZN(n852) );
  NOR2_X1 U959 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U960 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U961 ( .A(G164), .B(G162), .ZN(n856) );
  XNOR2_X1 U962 ( .A(n857), .B(n856), .ZN(n873) );
  NAND2_X1 U963 ( .A1(G139), .A2(n858), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G103), .A2(n859), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G127), .A2(n862), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G115), .A2(n863), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n994) );
  XOR2_X1 U971 ( .A(n994), .B(n1009), .Z(n871) );
  XOR2_X1 U972 ( .A(G160), .B(n869), .Z(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n877) );
  XOR2_X1 U975 ( .A(n875), .B(n874), .Z(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U977 ( .A1(G37), .A2(n878), .ZN(G395) );
  XOR2_X1 U978 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n880) );
  XNOR2_X1 U979 ( .A(G171), .B(n942), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n881), .B(G286), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U983 ( .A(n884), .B(n960), .Z(n885) );
  NOR2_X1 U984 ( .A1(G37), .A2(n885), .ZN(G397) );
  XNOR2_X1 U985 ( .A(KEYINPUT103), .B(n886), .ZN(G319) );
  XNOR2_X1 U986 ( .A(G1996), .B(KEYINPUT41), .ZN(n896) );
  XOR2_X1 U987 ( .A(G1971), .B(G1956), .Z(n888) );
  XNOR2_X1 U988 ( .A(G1991), .B(G1961), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U990 ( .A(G1976), .B(G1981), .Z(n890) );
  XNOR2_X1 U991 ( .A(G1986), .B(G1966), .ZN(n889) );
  XNOR2_X1 U992 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U993 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U994 ( .A(KEYINPUT104), .B(G2474), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(G229) );
  XOR2_X1 U997 ( .A(G2100), .B(G2096), .Z(n898) );
  XNOR2_X1 U998 ( .A(KEYINPUT42), .B(G2678), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U1000 ( .A(KEYINPUT43), .B(G2072), .Z(n900) );
  XNOR2_X1 U1001 ( .A(G2067), .B(G2090), .ZN(n899) );
  XNOR2_X1 U1002 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U1003 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U1004 ( .A(G2084), .B(G2078), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(n904), .B(n903), .ZN(G227) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n905) );
  XOR2_X1 U1007 ( .A(KEYINPUT113), .B(n905), .Z(n912) );
  XNOR2_X1 U1008 ( .A(KEYINPUT111), .B(KEYINPUT49), .ZN(n907) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1010 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n908), .ZN(n909) );
  NOR2_X1 U1012 ( .A1(G401), .A2(n909), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(KEYINPUT112), .B(n910), .ZN(n911) );
  NAND2_X1 U1014 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1017 ( .A(KEYINPUT125), .B(KEYINPUT62), .ZN(n1026) );
  XOR2_X1 U1018 ( .A(G29), .B(KEYINPUT120), .Z(n936) );
  XOR2_X1 U1019 ( .A(G2090), .B(G35), .Z(n916) );
  XNOR2_X1 U1020 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n913) );
  XNOR2_X1 U1021 ( .A(n913), .B(G34), .ZN(n914) );
  XNOR2_X1 U1022 ( .A(G2084), .B(n914), .ZN(n915) );
  NAND2_X1 U1023 ( .A1(n916), .A2(n915), .ZN(n933) );
  XNOR2_X1 U1024 ( .A(G27), .B(n917), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT117), .B(G2072), .ZN(n918) );
  XNOR2_X1 U1026 ( .A(n918), .B(G33), .ZN(n925) );
  XOR2_X1 U1027 ( .A(n919), .B(KEYINPUT116), .Z(n920) );
  XNOR2_X1 U1028 ( .A(n920), .B(G25), .ZN(n921) );
  NAND2_X1 U1029 ( .A1(n921), .A2(G28), .ZN(n923) );
  XNOR2_X1 U1030 ( .A(G26), .B(G2067), .ZN(n922) );
  NOR2_X1 U1031 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1032 ( .A1(n925), .A2(n924), .ZN(n928) );
  XNOR2_X1 U1033 ( .A(G32), .B(G1996), .ZN(n926) );
  XNOR2_X1 U1034 ( .A(KEYINPUT118), .B(n926), .ZN(n927) );
  NOR2_X1 U1035 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1036 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1037 ( .A(KEYINPUT53), .B(n931), .Z(n932) );
  NOR2_X1 U1038 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1039 ( .A(n934), .B(KEYINPUT55), .ZN(n935) );
  NAND2_X1 U1040 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1041 ( .A1(n937), .A2(G11), .ZN(n938) );
  XNOR2_X1 U1042 ( .A(n938), .B(KEYINPUT121), .ZN(n1024) );
  XNOR2_X1 U1043 ( .A(G16), .B(KEYINPUT56), .ZN(n966) );
  XOR2_X1 U1044 ( .A(G168), .B(G1966), .Z(n939) );
  NOR2_X1 U1045 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1046 ( .A(KEYINPUT57), .B(n941), .Z(n964) );
  XOR2_X1 U1047 ( .A(G1348), .B(n942), .Z(n944) );
  XOR2_X1 U1048 ( .A(G171), .B(G1961), .Z(n943) );
  NOR2_X1 U1049 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1050 ( .A(KEYINPUT122), .B(n945), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(n947), .B(n946), .ZN(n948) );
  NOR2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(G1971), .A2(G303), .ZN(n950) );
  NAND2_X1 U1054 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1059 ( .A(G1341), .B(n960), .Z(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n993) );
  INV_X1 U1063 ( .A(G16), .ZN(n991) );
  XNOR2_X1 U1064 ( .A(G5), .B(n967), .ZN(n980) );
  XNOR2_X1 U1065 ( .A(G1348), .B(KEYINPUT59), .ZN(n968) );
  XNOR2_X1 U1066 ( .A(n968), .B(G4), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G1956), .B(G20), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(G6), .B(G1981), .ZN(n969) );
  NOR2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1071 ( .A(KEYINPUT123), .B(G1341), .Z(n973) );
  XNOR2_X1 U1072 ( .A(G19), .B(n973), .ZN(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1074 ( .A(KEYINPUT60), .B(n976), .Z(n978) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G21), .ZN(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(G1986), .B(G24), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(G23), .B(G1976), .ZN(n981) );
  NOR2_X1 U1080 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1081 ( .A(G1971), .B(KEYINPUT124), .Z(n983) );
  XNOR2_X1 U1082 ( .A(G22), .B(n983), .ZN(n984) );
  NAND2_X1 U1083 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1084 ( .A(KEYINPUT58), .B(n986), .ZN(n987) );
  NOR2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1086 ( .A(KEYINPUT61), .B(n989), .ZN(n990) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n1022) );
  XOR2_X1 U1089 ( .A(G2072), .B(n994), .Z(n996) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n995) );
  NOR2_X1 U1091 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1092 ( .A(KEYINPUT50), .B(n997), .Z(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1008) );
  XOR2_X1 U1094 ( .A(G2090), .B(G162), .Z(n1000) );
  NOR2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1096 ( .A(KEYINPUT51), .B(n1002), .Z(n1004) );
  NAND2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XOR2_X1 U1098 ( .A(G160), .B(G2084), .Z(n1005) );
  NOR2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(n1011), .B(KEYINPUT114), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(n1016), .B(KEYINPUT52), .ZN(n1018) );
  INV_X1 U1106 ( .A(KEYINPUT55), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(G29), .A2(n1019), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(KEYINPUT115), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(n1026), .B(n1025), .ZN(G311) );
  XOR2_X1 U1113 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

