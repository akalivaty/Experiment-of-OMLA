//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1232, new_n1233;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n449), .B1(new_n457), .B2(new_n454), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR3_X1   g036(.A1(new_n460), .A2(new_n461), .A3(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT70), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n465), .A2(G101), .B1(G137), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G113), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(new_n461), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g051(.A(KEYINPUT68), .B(G125), .C1(new_n472), .C2(new_n473), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n469), .B1(new_n478), .B2(KEYINPUT69), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  AOI211_X1 g055(.A(new_n480), .B(new_n463), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n481), .ZN(G160));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(G124), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n468), .A2(G136), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n463), .C1(new_n472), .C2(new_n473), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n499), .A2(new_n500), .A3(G138), .A4(new_n463), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n496), .B1(new_n498), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n511), .A2(G50), .B1(new_n517), .B2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n504), .A2(KEYINPUT71), .ZN(new_n520));
  OAI21_X1  g095(.A(G651), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n513), .A2(new_n514), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .A4(new_n509), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT72), .B1(new_n508), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n518), .B1(new_n527), .B2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  AND3_X1   g105(.A1(new_n524), .A2(G89), .A3(new_n526), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n511), .A2(G51), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n515), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(KEYINPUT74), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(KEYINPUT74), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(G651), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n524), .A2(new_n526), .A3(G90), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n511), .A2(G52), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT75), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n547), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(G171));
  NAND3_X1  g126(.A1(new_n524), .A2(new_n526), .A3(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n515), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n511), .A2(G43), .B1(new_n555), .B2(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT77), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(KEYINPUT6), .B2(new_n503), .ZN(new_n567));
  XNOR2_X1  g142(.A(KEYINPUT71), .B(KEYINPUT6), .ZN(new_n568));
  OAI211_X1 g143(.A(G53), .B(new_n567), .C1(new_n568), .C2(new_n503), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n521), .A2(new_n571), .A3(G53), .A4(new_n567), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n524), .A2(new_n526), .A3(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n515), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  AND3_X1   g155(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n524), .A2(new_n526), .A3(G89), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G286));
  NAND3_X1  g158(.A1(new_n524), .A2(new_n526), .A3(G87), .ZN(new_n584));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n503), .B1(new_n515), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n511), .B2(G49), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(G288));
  NAND3_X1  g163(.A1(new_n524), .A2(new_n526), .A3(G86), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT78), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n524), .A2(new_n526), .A3(new_n591), .A4(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n511), .A2(new_n594), .A3(G48), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n567), .B1(new_n568), .B2(new_n503), .ZN(new_n596));
  INV_X1    g171(.A(G48), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT79), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n515), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n595), .A2(new_n598), .B1(G651), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n593), .A2(new_n602), .ZN(G305));
  AND2_X1   g178(.A1(new_n524), .A2(new_n526), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G85), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n515), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n511), .A2(G47), .B1(new_n608), .B2(G651), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT81), .B(G66), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n523), .A2(new_n612), .B1(G79), .B2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G54), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n613), .A2(new_n503), .B1(new_n596), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n604), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n527), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n615), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n611), .A2(KEYINPUT80), .B1(G868), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(KEYINPUT80), .B2(new_n611), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT82), .Z(G284));
  XOR2_X1   g198(.A(new_n622), .B(KEYINPUT83), .Z(G321));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(G299), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n625), .B2(G168), .ZN(G280));
  XOR2_X1   g202(.A(G280), .B(KEYINPUT84), .Z(G297));
  XNOR2_X1  g203(.A(KEYINPUT85), .B(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n620), .B1(G860), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT86), .Z(G148));
  NAND2_X1  g206(.A1(new_n620), .A2(new_n629), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n465), .A2(new_n499), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT13), .Z(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n468), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n486), .A2(G123), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n463), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G2096), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n640), .A2(new_n641), .A3(new_n648), .ZN(G156));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n663), .A3(G14), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT87), .Z(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n639), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n647), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n680), .A2(KEYINPUT89), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(KEYINPUT89), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n678), .A2(new_n679), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  MUX2_X1   g264(.A(new_n689), .B(new_n688), .S(new_n684), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NOR2_X1   g274(.A1(G168), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n699), .B2(G21), .ZN(new_n701));
  INV_X1    g276(.A(G1966), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT103), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT31), .B(G11), .Z(new_n705));
  INV_X1    g280(.A(G28), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(KEYINPUT30), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT104), .ZN(new_n708));
  AOI21_X1  g283(.A(G29), .B1(new_n706), .B2(KEYINPUT30), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n646), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n701), .B2(new_n702), .ZN(new_n713));
  INV_X1    g288(.A(G1961), .ZN(new_n714));
  NAND2_X1  g289(.A1(G301), .A2(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n699), .A2(G5), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n704), .B(new_n713), .C1(new_n714), .C2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT105), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n699), .A2(G20), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT23), .Z(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G299), .B2(G16), .ZN(new_n723));
  INV_X1    g298(.A(G1956), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n711), .A2(G35), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n711), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT29), .Z(new_n728));
  INV_X1    g303(.A(G2090), .ZN(new_n729));
  INV_X1    g304(.A(G2072), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT25), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n468), .A2(G139), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n499), .A2(G127), .ZN(new_n737));
  AND2_X1   g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  OAI21_X1  g313(.A(G2105), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n736), .A2(G29), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G29), .B2(G33), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n728), .A2(new_n729), .B1(new_n730), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G27), .A2(G29), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G164), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2078), .ZN(new_n745));
  INV_X1    g320(.A(new_n741), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(G2072), .ZN(new_n747));
  OR4_X1    g322(.A1(new_n725), .A2(new_n742), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n717), .A2(new_n714), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n465), .A2(G105), .B1(G141), .B2(new_n468), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT26), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G129), .B2(new_n486), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(G29), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G29), .A2(G32), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(KEYINPUT100), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT100), .B2(new_n754), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT101), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT27), .B(G1996), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT102), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n758), .A2(new_n760), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n699), .A2(G19), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n558), .B2(new_n699), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT96), .B(G1341), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT97), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n764), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n711), .A2(G26), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT28), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n468), .A2(G140), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n486), .A2(G128), .ZN(new_n771));
  OR2_X1    g346(.A1(G104), .A2(G2105), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n772), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n770), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n769), .B1(new_n775), .B2(new_n711), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2067), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n728), .B2(new_n729), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n761), .A2(new_n762), .A3(new_n767), .A4(new_n778), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n748), .A2(new_n749), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n718), .A2(new_n719), .ZN(new_n781));
  NOR2_X1   g356(.A1(G4), .A2(G16), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n620), .B2(G16), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT95), .B(G1348), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G34), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G160), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2084), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n720), .A2(new_n780), .A3(new_n781), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n699), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n699), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT93), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n699), .A2(G23), .ZN(new_n798));
  INV_X1    g373(.A(G288), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n699), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT92), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT33), .B(G1976), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n699), .A2(G6), .ZN(new_n804));
  INV_X1    g379(.A(G305), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n699), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n797), .A2(new_n803), .A3(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n468), .A2(G131), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT90), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G107), .B2(new_n463), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT91), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n486), .A2(G119), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n813), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G25), .B(new_n819), .S(G29), .Z(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G1986), .ZN(new_n823));
  INV_X1    g398(.A(G290), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n699), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n699), .B2(G24), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n822), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n823), .B2(new_n826), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n810), .A2(new_n811), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n831), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n792), .B1(new_n832), .B2(new_n833), .ZN(G311));
  INV_X1    g409(.A(KEYINPUT106), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n833), .ZN(new_n836));
  INV_X1    g411(.A(new_n792), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI211_X1 g413(.A(KEYINPUT106), .B(new_n792), .C1(new_n832), .C2(new_n833), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(G150));
  NAND2_X1  g415(.A1(new_n620), .A2(G559), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT38), .Z(new_n842));
  NAND3_X1  g417(.A1(new_n524), .A2(new_n526), .A3(G93), .ZN(new_n843));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n515), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n511), .A2(G55), .B1(new_n846), .B2(G651), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n557), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n552), .A2(new_n556), .A3(new_n843), .A4(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n842), .B(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT107), .B(G860), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n843), .B2(new_n847), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(G145));
  NAND2_X1  g434(.A1(new_n736), .A2(new_n739), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT108), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n750), .A2(new_n753), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n637), .B(new_n819), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n491), .A2(new_n495), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n500), .B1(new_n468), .B2(G138), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n774), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n468), .A2(G142), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n486), .A2(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n463), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n872), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n489), .B(new_n646), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G160), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n865), .A2(new_n878), .A3(new_n866), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n882), .B1(new_n880), .B2(new_n883), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g464(.A1(new_n848), .A2(new_n625), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n824), .A2(G305), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G303), .B(G288), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n824), .A2(G305), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n893), .ZN(new_n896));
  INV_X1    g471(.A(new_n894), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n897), .B2(new_n891), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(KEYINPUT109), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(KEYINPUT109), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n632), .B(new_n851), .Z(new_n905));
  INV_X1    g480(.A(G299), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n620), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n620), .A2(new_n906), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n907), .B2(new_n908), .ZN(new_n912));
  INV_X1    g487(.A(new_n620), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n620), .A2(new_n906), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(KEYINPUT41), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n910), .B1(new_n905), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n904), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n890), .B1(new_n919), .B2(new_n625), .ZN(G295));
  OAI21_X1  g495(.A(new_n890), .B1(new_n919), .B2(new_n625), .ZN(G331));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n531), .B2(new_n537), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n849), .A2(new_n924), .A3(new_n850), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n924), .B1(new_n849), .B2(new_n850), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n581), .A2(KEYINPUT110), .A3(new_n582), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n547), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n928), .B(new_n544), .C1(new_n548), .C2(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n924), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n851), .A2(new_n932), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n933), .A2(new_n925), .B1(G171), .B2(new_n928), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n912), .B(new_n916), .C1(new_n931), .C2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n930), .B1(new_n926), .B2(new_n927), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n933), .A2(G171), .A3(new_n928), .A4(new_n925), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n909), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n899), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(G37), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(new_n899), .A3(new_n938), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n935), .A2(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n900), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n885), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT111), .B1(new_n939), .B2(G37), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n922), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n941), .A3(new_n950), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(KEYINPUT112), .A3(KEYINPUT43), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT112), .B1(new_n953), .B2(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n949), .A2(new_n940), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n952), .B1(new_n959), .B2(new_n922), .ZN(G397));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n479), .A2(new_n961), .A3(new_n481), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT45), .B1(new_n871), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1996), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT46), .ZN(new_n969));
  INV_X1    g544(.A(G2067), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n774), .B(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n971), .A2(new_n750), .A3(new_n753), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n965), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n974));
  XNOR2_X1  g549(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n965), .A2(new_n971), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT113), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n862), .B(G1996), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n966), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n821), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n819), .A2(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n979), .A2(new_n981), .B1(new_n970), .B2(new_n775), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n975), .B1(new_n982), .B2(new_n965), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n819), .B(new_n821), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n979), .B1(new_n965), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT126), .Z(new_n986));
  NAND2_X1  g561(.A1(new_n824), .A2(new_n823), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(new_n965), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT48), .Z(new_n989));
  AOI21_X1  g564(.A(new_n983), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT124), .ZN(new_n991));
  NAND2_X1  g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n965), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n985), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1981), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n593), .A2(new_n995), .A3(new_n602), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n602), .A2(new_n589), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G1981), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n468), .A2(G137), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n462), .A2(new_n464), .ZN(new_n1003));
  INV_X1    g578(.A(G101), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G125), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n466), .B2(new_n467), .ZN(new_n1007));
  OAI22_X1  g582(.A1(new_n1007), .A2(KEYINPUT68), .B1(new_n470), .B2(new_n461), .ZN(new_n1008));
  INV_X1    g583(.A(new_n477), .ZN(new_n1009));
  OAI21_X1  g584(.A(G2105), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1005), .B1(new_n1010), .B2(new_n480), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n478), .A2(KEYINPUT69), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G164), .A2(G1384), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1011), .A2(G40), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G8), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n996), .A2(new_n998), .A3(KEYINPUT49), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1001), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n799), .A2(G1976), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(G8), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT52), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT114), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n799), .B2(G1976), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1020), .A2(new_n1027), .A3(KEYINPUT52), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1018), .A2(new_n1022), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G303), .A2(G8), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT55), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1010), .A2(new_n480), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1033), .A2(G40), .A3(new_n1012), .A4(new_n469), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(G164), .B2(G1384), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n871), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n796), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n871), .A2(new_n1041), .A3(new_n963), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n962), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1039), .B1(new_n1044), .B2(G2090), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1032), .A2(new_n1045), .A3(G8), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1029), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1039), .B(KEYINPUT115), .C1(new_n1044), .C2(G2090), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1034), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n729), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT115), .B1(new_n1053), .B2(new_n1039), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1031), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT116), .B(new_n1031), .C1(new_n1050), .C2(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n498), .A2(new_n501), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n1035), .B(G1384), .C1(new_n1059), .C2(new_n868), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n964), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n962), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2084), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1062), .A2(new_n702), .B1(new_n1052), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1064), .A2(new_n1065), .A3(G286), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1048), .A2(new_n1057), .A3(new_n1058), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT63), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1045), .A2(G8), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1031), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1048), .A2(KEYINPUT63), .A3(new_n1066), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1029), .A2(new_n1046), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1018), .ZN(new_n1075));
  OR2_X1    g650(.A1(G288), .A2(G1976), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n996), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1016), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1058), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  AOI21_X1  g655(.A(G1971), .B1(new_n962), .B2(new_n1061), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1034), .A2(new_n1051), .A3(G2090), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(G8), .A3(new_n1049), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT116), .B1(new_n1084), .B2(new_n1031), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1015), .B1(new_n999), .B2(new_n1000), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1025), .B1(new_n1086), .B2(new_n1017), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1087), .A2(new_n1046), .A3(new_n1028), .A4(new_n1022), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1079), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G168), .A2(new_n1065), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT51), .B1(new_n1090), .B2(KEYINPUT119), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1091), .B(new_n1092), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1092), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1044), .A2(G2084), .B1(new_n1095), .B2(G1966), .ZN(new_n1096));
  OAI211_X1 g671(.A(G8), .B(new_n1094), .C1(new_n1096), .C2(G286), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1093), .A2(new_n1097), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(G2078), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n961), .B(new_n1102), .C1(new_n1005), .C2(KEYINPUT121), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(KEYINPUT121), .B2(new_n1005), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n478), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1061), .A2(new_n1105), .B1(new_n1044), .B2(new_n714), .ZN(new_n1106));
  INV_X1    g681(.A(G2078), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n962), .A2(new_n1061), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1100), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1108), .B2(new_n1100), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1106), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1099), .B1(new_n1113), .B2(G171), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1062), .A2(new_n1102), .B1(new_n1052), .B2(G1961), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1034), .A2(new_n1038), .A3(G2078), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT120), .B1(new_n1116), .B2(KEYINPUT53), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1117), .B2(new_n1110), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G301), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1098), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n714), .A2(new_n1044), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(G171), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1106), .B(G301), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n1121), .B(KEYINPUT54), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1118), .B2(G301), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT122), .B1(new_n1127), .B2(new_n1099), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1089), .B(new_n1120), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(G1348), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1044), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n962), .A2(new_n970), .A3(new_n1013), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n913), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n962), .A2(new_n1061), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n724), .B1(new_n1034), .B2(new_n1051), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G299), .B(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(G1956), .B1(new_n962), .B2(new_n1043), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1134), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1034), .A2(new_n1038), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1135), .A2(new_n1136), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1138), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1140), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n620), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT60), .A4(new_n913), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1153), .A2(new_n1154), .B1(new_n1152), .B2(new_n1151), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT58), .B(G1341), .Z(new_n1156));
  AOI22_X1  g731(.A1(new_n1095), .A2(new_n967), .B1(new_n1014), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT59), .B1(new_n1157), .B2(new_n557), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n962), .A2(new_n1061), .A3(new_n967), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1014), .A2(new_n1156), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1161), .A2(new_n1162), .A3(new_n558), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1138), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1135), .A2(new_n1136), .A3(new_n1145), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1145), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1169), .A2(new_n1170), .A3(new_n1138), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1139), .A2(KEYINPUT61), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1164), .B(new_n1168), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1155), .B1(new_n1173), .B2(KEYINPUT118), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1148), .A2(KEYINPUT61), .A3(new_n1139), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1175), .A2(new_n1176), .A3(new_n1168), .A4(new_n1164), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1150), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1073), .B(new_n1078), .C1(new_n1129), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1096), .A2(new_n1090), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1124), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1048), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT123), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1124), .B1(new_n1098), .B2(new_n1181), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1089), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1098), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT62), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1187), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n991), .B(new_n994), .C1(new_n1179), .C2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1162), .B1(new_n1161), .B2(new_n558), .ZN(new_n1197));
  AOI211_X1 g772(.A(KEYINPUT59), .B(new_n557), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1198));
  OAI22_X1  g773(.A1(new_n1196), .A2(KEYINPUT61), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1170), .A2(new_n1138), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1172), .B1(new_n1200), .B2(new_n1146), .ZN(new_n1201));
  OAI21_X1  g776(.A(KEYINPUT118), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1155), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1202), .A2(new_n1177), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1149), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1127), .A2(new_n1099), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1121), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1127), .A2(KEYINPUT122), .A3(new_n1099), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1113), .A2(G171), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1210), .A2(KEYINPUT54), .A3(new_n1119), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1191), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1212), .A2(new_n1186), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1205), .A2(new_n1209), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1187), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1214), .A2(new_n1215), .A3(new_n1073), .A4(new_n1078), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n991), .B1(new_n1216), .B2(new_n994), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n990), .B1(new_n1195), .B2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n1220));
  NOR3_X1   g794(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1221));
  OAI211_X1 g795(.A(new_n697), .B(new_n1221), .C1(new_n886), .C2(new_n887), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n1223));
  INV_X1    g797(.A(KEYINPUT112), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n958), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI211_X1 g799(.A(new_n1220), .B(new_n1222), .C1(new_n1225), .C2(new_n954), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1227));
  NAND3_X1  g801(.A1(new_n1227), .A2(new_n954), .A3(new_n957), .ZN(new_n1228));
  INV_X1    g802(.A(new_n1222), .ZN(new_n1229));
  AOI21_X1  g803(.A(KEYINPUT127), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g804(.A1(new_n1226), .A2(new_n1230), .ZN(G308));
  OAI21_X1  g805(.A(new_n1220), .B1(new_n959), .B2(new_n1222), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n1228), .A2(KEYINPUT127), .A3(new_n1229), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1232), .A2(new_n1233), .ZN(G225));
endmodule


