//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1323, new_n1324, new_n1325, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OR2_X1    g0004(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n206));
  NAND3_X1  g0006(.A1(new_n205), .A2(G50), .A3(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n210), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT65), .B(G68), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n222), .B1(G238), .B2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT66), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n227), .B(new_n228), .C1(new_n224), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n215), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n218), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT69), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT67), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT70), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G58), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(new_n213), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n209), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT8), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT8), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n213), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n258), .A2(new_n265), .B1(new_n253), .B2(new_n263), .ZN(new_n266));
  XOR2_X1   g0066(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n267));
  INV_X1    g0067(.A(new_n223), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT79), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT7), .B1(new_n274), .B2(new_n210), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT7), .ZN(new_n276));
  AOI211_X1 g0076(.A(new_n276), .B(G20), .C1(new_n271), .C2(new_n273), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n269), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n279), .B2(G20), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT79), .B1(new_n280), .B2(KEYINPUT7), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n268), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n201), .B1(new_n223), .B2(G58), .ZN(new_n283));
  INV_X1    g0083(.A(G159), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n283), .A2(new_n210), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n267), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n256), .ZN(new_n289));
  INV_X1    g0089(.A(G68), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n272), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n292));
  OAI211_X1 g0092(.A(KEYINPUT7), .B(new_n210), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(new_n280), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n289), .B1(new_n295), .B2(KEYINPUT16), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n266), .B1(new_n288), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  INV_X1    g0102(.A(new_n209), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n301), .A2(G232), .B1(new_n305), .B2(new_n300), .ZN(new_n306));
  INV_X1    g0106(.A(G1698), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n271), .A2(new_n273), .A3(G223), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G87), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n271), .A2(new_n273), .A3(G226), .A4(G1698), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT80), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n279), .A2(KEYINPUT80), .A3(G226), .A4(G1698), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n304), .A2(G1), .A3(G13), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n306), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G200), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n306), .B(G190), .C1(new_n315), .C2(new_n316), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n297), .A2(new_n321), .A3(KEYINPUT17), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT17), .ZN(new_n323));
  INV_X1    g0123(.A(new_n266), .ZN(new_n324));
  INV_X1    g0124(.A(new_n267), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT79), .B1(new_n280), .B2(new_n293), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n274), .A2(new_n210), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n269), .B1(new_n327), .B2(new_n276), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n223), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT65), .A2(G68), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT65), .A2(G68), .ZN(new_n331));
  OAI21_X1  g0131(.A(G58), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n202), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(G20), .B1(G159), .B2(new_n285), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n325), .B1(new_n329), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(G68), .B1(new_n275), .B2(new_n277), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT16), .A3(new_n334), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n256), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n324), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n323), .B1(new_n339), .B2(new_n320), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n322), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT18), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n317), .A2(G169), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n306), .B(G179), .C1(new_n315), .C2(new_n316), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n339), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n342), .B1(new_n339), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT81), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n343), .A2(new_n344), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT18), .B1(new_n297), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT81), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n339), .A2(new_n342), .A3(new_n345), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n341), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n285), .A2(G50), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT76), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n210), .A2(G33), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n223), .A2(new_n210), .B1(new_n220), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n256), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT11), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(KEYINPUT11), .B(new_n256), .C1(new_n356), .C2(new_n358), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n223), .B2(new_n253), .ZN(new_n364));
  OR3_X1    g0164(.A1(new_n253), .A2(KEYINPUT12), .A3(G68), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n290), .B1(new_n213), .B2(G20), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n364), .A2(new_n365), .B1(new_n257), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  OR2_X1    g0168(.A1(G226), .A2(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(G232), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G1698), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n271), .A2(new_n369), .A3(new_n273), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G97), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(KEYINPUT74), .A3(new_n298), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n300), .A2(new_n316), .A3(G274), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n316), .A2(G238), .A3(new_n299), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n316), .B1(new_n372), .B2(new_n373), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(KEYINPUT74), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT13), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  NOR2_X1   g0183(.A1(G226), .A2(G1698), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n370), .B2(G1698), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n279), .B1(G33), .B2(G97), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n316), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT13), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(new_n375), .A4(new_n378), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n368), .B1(new_n390), .B2(G200), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(KEYINPUT75), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n376), .A2(new_n377), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n380), .B2(KEYINPUT74), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n394), .A2(new_n387), .A3(new_n395), .A4(new_n388), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n392), .A2(G190), .A3(new_n396), .A4(new_n382), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n389), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n388), .B1(new_n394), .B2(new_n387), .ZN(new_n401));
  OAI21_X1  g0201(.A(G169), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT14), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n382), .B2(new_n389), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n392), .A2(G179), .A3(new_n396), .A4(new_n382), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n399), .B1(new_n368), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT8), .B(G58), .ZN(new_n411));
  INV_X1    g0211(.A(G150), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n411), .A2(new_n357), .B1(new_n412), .B2(new_n286), .ZN(new_n413));
  INV_X1    g0213(.A(G50), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n210), .B1(new_n201), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n256), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n213), .B2(G20), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n257), .A2(new_n417), .B1(new_n414), .B2(new_n254), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n301), .A2(G226), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n376), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n279), .A2(G222), .A3(new_n307), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n279), .A2(G223), .A3(G1698), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n423), .C1(new_n220), .C2(new_n279), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n421), .B1(new_n424), .B2(new_n298), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n419), .B1(new_n425), .B2(G169), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n298), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n376), .A3(new_n420), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G179), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT9), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n419), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g0232(.A(new_n432), .B(KEYINPUT73), .Z(new_n433));
  AND2_X1   g0233(.A1(new_n416), .A2(new_n418), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n428), .A2(G200), .B1(new_n434), .B2(KEYINPUT9), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n425), .A2(G190), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT10), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G200), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n425), .A2(new_n439), .B1(new_n419), .B2(new_n431), .ZN(new_n440));
  INV_X1    g0240(.A(G190), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n428), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT10), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n432), .B(KEYINPUT73), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n430), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n264), .A2(G77), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n258), .A2(new_n448), .B1(G77), .B2(new_n253), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n263), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT71), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT15), .B(G87), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(new_n357), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n270), .A2(G20), .ZN(new_n454));
  INV_X1    g0254(.A(G87), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n455), .A2(KEYINPUT15), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(KEYINPUT15), .ZN(new_n457));
  OAI211_X1 g0257(.A(KEYINPUT71), .B(new_n454), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n450), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n256), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT72), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(KEYINPUT72), .A3(new_n256), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n449), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n301), .A2(G244), .B1(new_n305), .B2(new_n300), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G232), .A2(G1698), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n307), .A2(G238), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n279), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n298), .C1(G107), .C2(new_n279), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n470), .A2(new_n439), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(G190), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n464), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n449), .ZN(new_n474));
  INV_X1    g0274(.A(new_n463), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT72), .B1(new_n459), .B2(new_n256), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(G169), .B1(new_n465), .B2(new_n469), .ZN(new_n478));
  INV_X1    g0278(.A(G179), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n470), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n354), .A2(new_n410), .A3(new_n447), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n213), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n253), .A2(new_n486), .A3(new_n209), .A4(new_n255), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G97), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n253), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n488), .A2(KEYINPUT83), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT83), .B1(new_n488), .B2(new_n490), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(G107), .B1(new_n326), .B2(new_n328), .ZN(new_n494));
  XNOR2_X1  g0294(.A(G97), .B(G107), .ZN(new_n495));
  NOR2_X1   g0295(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(KEYINPUT6), .B2(new_n489), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n498), .B(G20), .C1(new_n495), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n285), .A2(G77), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n493), .B1(new_n504), .B2(new_n256), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n271), .A2(new_n273), .A3(G244), .A4(new_n307), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n307), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n508), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n298), .ZN(new_n513));
  INV_X1    g0313(.A(G45), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G1), .ZN(new_n515));
  AND2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT5), .A2(G41), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(G257), .A3(new_n316), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT5), .B(G41), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n520), .A2(G274), .A3(new_n316), .A4(new_n515), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n513), .A2(new_n523), .A3(new_n479), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n522), .B1(new_n512), .B2(new_n298), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(G169), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n485), .B1(new_n505), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n493), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n278), .A2(new_n281), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n502), .B1(new_n529), .B2(G107), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n530), .B2(new_n289), .ZN(new_n531));
  AOI211_X1 g0331(.A(G179), .B(new_n522), .C1(new_n512), .C2(new_n298), .ZN(new_n532));
  AOI21_X1  g0332(.A(G169), .B1(new_n513), .B2(new_n523), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n534), .A3(KEYINPUT84), .ZN(new_n535));
  INV_X1    g0335(.A(new_n525), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n525), .A2(G190), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n505), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n527), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n271), .A2(new_n273), .A3(G244), .A4(G1698), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n271), .A2(new_n273), .A3(G238), .A4(new_n307), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G116), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n298), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n316), .A2(G274), .A3(new_n515), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n213), .A2(G45), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n316), .A2(G250), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n545), .A2(G190), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n439), .B1(new_n545), .B2(new_n550), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n454), .A2(new_n554), .A3(G97), .ZN(new_n555));
  NOR2_X1   g0355(.A1(G97), .A2(G107), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n455), .B1(new_n373), .B2(new_n210), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n557), .B2(new_n554), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n279), .A2(KEYINPUT85), .A3(new_n210), .A4(G68), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n271), .A2(new_n273), .A3(new_n210), .A4(G68), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT85), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n256), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n452), .A2(new_n254), .ZN(new_n565));
  INV_X1    g0365(.A(new_n487), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G87), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n545), .A2(G179), .A3(new_n550), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n549), .B1(new_n544), .B2(new_n298), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n404), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n452), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n564), .A2(new_n565), .A3(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n553), .A2(new_n568), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n271), .A2(new_n273), .A3(G250), .A4(new_n307), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT93), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n279), .A2(KEYINPUT93), .A3(G250), .A4(new_n307), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n279), .A2(G257), .A3(G1698), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G294), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n298), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n518), .A2(G264), .A3(new_n316), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n584), .A2(new_n521), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n441), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(KEYINPUT94), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT94), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n518), .A2(new_n589), .A3(G264), .A4(new_n316), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n583), .A2(new_n521), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n439), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n210), .B2(G107), .ZN(new_n596));
  INV_X1    g0396(.A(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(KEYINPUT23), .A3(G20), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT91), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n543), .B2(G20), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n210), .A2(KEYINPUT91), .A3(G33), .A4(G116), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n271), .A2(new_n273), .A3(new_n210), .A4(G87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT22), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT22), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n279), .A2(new_n606), .A3(new_n210), .A4(G87), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n256), .B1(new_n608), .B2(KEYINPUT24), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT24), .ZN(new_n610));
  AOI211_X1 g0410(.A(new_n610), .B(new_n603), .C1(new_n605), .C2(new_n607), .ZN(new_n611));
  OR3_X1    g0411(.A1(new_n253), .A2(KEYINPUT25), .A3(G107), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT25), .B1(new_n253), .B2(G107), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n597), .C2(new_n487), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n614), .A2(KEYINPUT92), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(KEYINPUT92), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n609), .A2(new_n611), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n575), .B1(new_n594), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n540), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT95), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n583), .A2(G179), .A3(new_n521), .A4(new_n591), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n404), .B1(new_n583), .B2(new_n585), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(KEYINPUT95), .B(new_n621), .C1(new_n586), .C2(new_n404), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n617), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n518), .A2(G270), .A3(new_n316), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n521), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT86), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT86), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n630), .A3(new_n521), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n271), .A2(new_n273), .A3(G264), .A4(G1698), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT87), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n279), .A2(KEYINPUT87), .A3(G264), .A4(G1698), .ZN(new_n636));
  INV_X1    g0436(.A(G303), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT88), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT88), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G303), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n274), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n279), .A2(G257), .A3(new_n307), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n635), .A2(new_n636), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(KEYINPUT89), .A3(new_n298), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n632), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT90), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n298), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n510), .B(new_n210), .C1(G33), .C2(new_n489), .ZN(new_n651));
  INV_X1    g0451(.A(G116), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G20), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n256), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n651), .A2(KEYINPUT20), .A3(new_n256), .A4(new_n653), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n253), .A2(G116), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n566), .B2(G116), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n479), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n646), .A2(new_n647), .A3(new_n650), .A4(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n650), .A2(new_n645), .A3(new_n632), .A4(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT90), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n650), .A2(new_n645), .A3(new_n632), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G200), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n658), .A2(new_n660), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n650), .A2(G190), .A3(new_n645), .A4(new_n632), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n668), .A2(new_n404), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT21), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n666), .A2(new_n671), .A3(KEYINPUT21), .ZN(new_n675));
  AND4_X1   g0475(.A1(new_n665), .A2(new_n670), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n484), .A2(new_n619), .A3(new_n626), .A4(new_n676), .ZN(G372));
  NOR2_X1   g0477(.A1(new_n346), .A2(new_n347), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n477), .A2(new_n480), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n409), .A2(new_n368), .B1(new_n398), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n678), .B1(new_n680), .B2(new_n341), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n438), .A2(new_n446), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n430), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n575), .A2(new_n684), .A3(new_n531), .A4(new_n534), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n571), .A2(KEYINPUT96), .A3(new_n574), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT96), .B1(new_n571), .B2(new_n574), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n505), .A2(new_n526), .A3(new_n485), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT84), .B1(new_n531), .B2(new_n534), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n575), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n689), .B1(new_n692), .B2(KEYINPUT26), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n527), .A2(new_n535), .A3(new_n539), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n617), .B1(new_n622), .B2(new_n623), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n665), .A2(new_n674), .A3(new_n675), .A4(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n617), .B1(new_n587), .B2(new_n593), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n553), .A2(new_n568), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n571), .A2(new_n574), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n694), .A2(new_n696), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n683), .B1(new_n483), .B2(new_n704), .ZN(G369));
  INV_X1    g0505(.A(G330), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n674), .A2(new_n675), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n707), .A2(new_n665), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n213), .A2(new_n210), .A3(G13), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(KEYINPUT27), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(KEYINPUT27), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G213), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G343), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OR3_X1    g0515(.A1(new_n708), .A2(new_n668), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n676), .B1(new_n668), .B2(new_n715), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n706), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n697), .B1(new_n617), .B2(new_n714), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n626), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n626), .A2(new_n715), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n708), .A2(new_n714), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n626), .A3(new_n719), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n695), .A2(new_n714), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT97), .Z(G399));
  INV_X1    g0530(.A(new_n216), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G41), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n556), .A2(new_n455), .A3(new_n652), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(G1), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n207), .B2(new_n733), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n531), .A2(new_n534), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n739), .B2(new_n700), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n688), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n700), .B1(new_n527), .B2(new_n535), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n741), .B1(new_n684), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n707), .A2(new_n626), .A3(new_n665), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n619), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n714), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(KEYINPUT99), .A3(KEYINPUT29), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n740), .A2(new_n688), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n742), .A2(new_n684), .ZN(new_n749));
  AND4_X1   g0549(.A1(new_n626), .A2(new_n665), .A3(new_n674), .A4(new_n675), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n701), .A2(new_n527), .A3(new_n535), .A4(new_n539), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n748), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(KEYINPUT29), .A3(new_n715), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT99), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n714), .B1(new_n693), .B2(new_n702), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(KEYINPUT29), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n747), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT30), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n545), .A2(G179), .A3(new_n550), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n760), .A2(new_n525), .A3(new_n583), .A4(new_n591), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n759), .B1(new_n666), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT98), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT98), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n764), .B(new_n759), .C1(new_n666), .C2(new_n761), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n666), .A2(new_n761), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT30), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n570), .A2(G179), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n592), .A2(new_n536), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n666), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n763), .A2(new_n765), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n714), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT31), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n767), .A2(new_n762), .A3(new_n770), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n715), .A2(new_n773), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n619), .A2(new_n676), .A3(new_n626), .A4(new_n715), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n706), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n758), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n738), .B1(new_n779), .B2(G1), .ZN(G364));
  AND2_X1   g0580(.A1(new_n210), .A2(G13), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n213), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n732), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n718), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n716), .A2(new_n717), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(G330), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT100), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n209), .B1(G20), .B2(new_n404), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n210), .A2(new_n479), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n210), .A2(G179), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n795), .A2(new_n441), .A3(G200), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n794), .A2(new_n290), .B1(new_n796), .B2(new_n597), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n479), .A2(new_n439), .A3(G190), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G20), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n489), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G190), .A2(G200), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n795), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n284), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT32), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n791), .A2(new_n803), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n279), .B1(new_n807), .B2(new_n220), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n791), .A2(G190), .A3(new_n439), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(G58), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n792), .A2(new_n441), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n795), .A2(G190), .A3(G200), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n812), .A2(G50), .B1(new_n814), .B2(G87), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n802), .A2(new_n806), .A3(new_n811), .A4(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n817), .A2(new_n796), .B1(new_n813), .B2(new_n637), .ZN(new_n818));
  XNOR2_X1  g0618(.A(KEYINPUT33), .B(G317), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(new_n793), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n804), .B(KEYINPUT103), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G329), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n274), .B1(new_n807), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G322), .B2(new_n810), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n812), .A2(G326), .B1(G294), .B2(new_n799), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n820), .A2(new_n822), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n790), .B1(new_n816), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n784), .B(KEYINPUT101), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n731), .A2(new_n274), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT102), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G355), .B1(new_n652), .B2(new_n731), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n251), .A2(new_n514), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n731), .A2(new_n279), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n207), .B2(G45), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n833), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(G13), .A2(G33), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(G20), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n789), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n828), .B(new_n830), .C1(new_n837), .C2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT104), .Z(new_n843));
  INV_X1    g0643(.A(new_n840), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n786), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n788), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G396));
  OAI21_X1  g0648(.A(KEYINPUT106), .B1(new_n464), .B2(new_n715), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT106), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n477), .A2(new_n850), .A3(new_n714), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n849), .A2(new_n473), .A3(new_n851), .A4(new_n481), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT107), .B1(new_n481), .B2(new_n715), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT107), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n679), .A2(new_n854), .A3(new_n714), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n756), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n756), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n776), .A2(new_n777), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(G330), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n784), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n860), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n789), .A2(new_n838), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n830), .B1(new_n220), .B2(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n455), .A2(new_n796), .B1(new_n813), .B2(new_n597), .ZN(new_n867));
  INV_X1    g0667(.A(G294), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n274), .B1(new_n807), .B2(new_n652), .C1(new_n868), .C2(new_n809), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n801), .B(new_n869), .C1(G303), .C2(new_n812), .ZN(new_n870));
  INV_X1    g0670(.A(new_n821), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n823), .B2(new_n871), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n867), .B(new_n872), .C1(G283), .C2(new_n793), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(KEYINPUT105), .ZN(new_n875));
  INV_X1    g0675(.A(new_n807), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n810), .A2(G143), .B1(new_n876), .B2(G159), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n812), .A2(G137), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n877), .B(new_n878), .C1(new_n412), .C2(new_n794), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT34), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n821), .A2(G132), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n414), .A2(new_n813), .B1(new_n796), .B2(new_n290), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n274), .B(new_n884), .C1(G58), .C2(new_n799), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n874), .A2(KEYINPUT105), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n875), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI221_X1 g0688(.A(new_n866), .B1(new_n839), .B2(new_n857), .C1(new_n888), .C2(new_n790), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n864), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(G384));
  OAI21_X1  g0691(.A(new_n498), .B1(new_n495), .B2(new_n499), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(G116), .B(new_n211), .C1(new_n893), .C2(KEYINPUT35), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT108), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(KEYINPUT35), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(KEYINPUT108), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT36), .Z(new_n900));
  NAND3_X1  g0700(.A1(new_n208), .A2(G77), .A3(new_n332), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n414), .A2(G68), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n213), .B(G13), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n297), .A2(new_n321), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n337), .B(new_n256), .C1(new_n295), .C2(new_n325), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n324), .ZN(new_n908));
  INV_X1    g0708(.A(new_n712), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n908), .B1(new_n345), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n905), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n339), .A2(new_n345), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n339), .A2(new_n909), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n906), .A2(new_n913), .A3(new_n914), .A4(new_n905), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n908), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n712), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n916), .B1(new_n354), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(KEYINPUT38), .B(new_n916), .C1(new_n354), .C2(new_n919), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n408), .B1(new_n406), .B2(new_n405), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n402), .A2(KEYINPUT14), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n368), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n368), .A2(new_n714), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n927), .A2(new_n398), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n927), .B2(new_n398), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n857), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n771), .A2(KEYINPUT31), .A3(new_n714), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT31), .B1(new_n771), .B2(new_n714), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n777), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT40), .B1(new_n924), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n350), .A2(new_n352), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n339), .B(new_n909), .C1(new_n937), .C2(new_n341), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n906), .A2(new_n913), .A3(new_n914), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT37), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n915), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n921), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n923), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n772), .A2(new_n773), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n771), .A2(KEYINPUT31), .A3(new_n714), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n777), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n927), .A2(new_n398), .A3(new_n928), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n368), .B(new_n714), .C1(new_n399), .C2(new_n409), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n856), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n947), .A2(KEYINPUT40), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n936), .B1(new_n944), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n484), .A2(new_n947), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n706), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n953), .B2(new_n955), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT39), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n944), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n923), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n927), .A2(new_n714), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n678), .A2(new_n909), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n929), .A2(new_n930), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n481), .A2(new_n714), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n859), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n963), .B1(new_n967), .B2(new_n924), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n683), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n758), .B2(new_n484), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n969), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n957), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n213), .B2(new_n781), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n957), .A2(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n904), .B1(new_n974), .B2(new_n975), .ZN(G367));
  INV_X1    g0776(.A(new_n835), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n238), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n841), .B1(new_n216), .B2(new_n452), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n829), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n800), .A2(new_n290), .ZN(new_n981));
  INV_X1    g0781(.A(G143), .ZN(new_n982));
  INV_X1    g0782(.A(new_n812), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n982), .A2(new_n983), .B1(new_n794), .B2(new_n284), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n981), .B(new_n984), .C1(G58), .C2(new_n814), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n810), .A2(G150), .ZN(new_n986));
  INV_X1    g0786(.A(new_n804), .ZN(new_n987));
  XNOR2_X1  g0787(.A(KEYINPUT115), .B(G137), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G50), .A2(new_n876), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n279), .B1(new_n796), .B2(new_n220), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT114), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n985), .A2(new_n986), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n274), .B1(new_n804), .B2(new_n993), .C1(new_n489), .C2(new_n796), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT113), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n800), .A2(new_n597), .ZN(new_n997));
  INV_X1    g0797(.A(new_n641), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n998), .A2(new_n809), .B1(new_n807), .B2(new_n817), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(G311), .C2(new_n812), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n814), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT46), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n813), .B2(new_n652), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1001), .B(new_n1003), .C1(new_n794), .C2(new_n868), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT112), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n995), .A2(KEYINPUT113), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n996), .A2(new_n1000), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1004), .A2(KEYINPUT112), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n992), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n980), .B1(new_n1010), .B2(new_n789), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n568), .A2(new_n715), .ZN(new_n1012));
  MUX2_X1   g0812(.A(new_n700), .B(new_n688), .S(new_n1012), .Z(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n840), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n694), .B1(new_n505), .B2(new_n715), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n531), .A2(new_n534), .A3(new_n714), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n726), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT42), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n527), .B(new_n535), .C1(new_n1024), .C2(new_n626), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1027), .B1(new_n715), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT109), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1018), .B(new_n1020), .C1(new_n1030), .C2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1031), .B(KEYINPUT109), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1035), .A2(new_n1017), .A3(new_n1013), .A4(new_n1029), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n723), .A2(new_n1024), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(KEYINPUT110), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT110), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1034), .A2(new_n1036), .A3(new_n1042), .A4(new_n1038), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n728), .A2(new_n1024), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT45), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT44), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1023), .B1(KEYINPUT111), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n728), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1048), .A2(KEYINPUT111), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n724), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1045), .B(KEYINPUT45), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1051), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1050), .B(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n723), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n726), .B1(new_n722), .B2(new_n725), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(new_n718), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n779), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n732), .B(KEYINPUT41), .Z(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n783), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1016), .B1(new_n1044), .B2(new_n1065), .ZN(G387));
  OR2_X1    g0866(.A1(new_n779), .A2(new_n1060), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n779), .A2(new_n1060), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n732), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n720), .A2(new_n721), .A3(new_n840), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n835), .B1(new_n243), .B2(new_n514), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n832), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1071), .B1(new_n735), .B2(new_n1072), .ZN(new_n1073));
  OR3_X1    g0873(.A1(new_n411), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1074));
  OAI21_X1  g0874(.A(KEYINPUT50), .B1(new_n411), .B2(G50), .ZN(new_n1075));
  AOI21_X1  g0875(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1074), .A2(new_n735), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1073), .A2(new_n1077), .B1(new_n597), .B2(new_n731), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n841), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n829), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n807), .A2(new_n290), .B1(new_n804), .B2(new_n412), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n274), .B(new_n1081), .C1(G50), .C2(new_n810), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n814), .A2(G77), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n793), .A2(new_n263), .B1(new_n572), .B2(new_n799), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n796), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n812), .A2(G159), .B1(new_n1085), .B2(G97), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n279), .B1(new_n987), .B2(G326), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n800), .A2(new_n817), .B1(new_n813), .B2(new_n868), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n810), .A2(G317), .B1(new_n876), .B2(new_n641), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n812), .A2(G322), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n823), .C2(new_n794), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1089), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1093), .B2(new_n1092), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT49), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1088), .B1(new_n652), .B2(new_n796), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1087), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT116), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n790), .B1(new_n1099), .B2(KEYINPUT116), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1080), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1060), .A2(new_n783), .B1(new_n1070), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1069), .A2(new_n1103), .ZN(G393));
  INV_X1    g0904(.A(new_n1058), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1024), .A2(new_n840), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n841), .B1(new_n489), .B2(new_n216), .C1(new_n248), .C2(new_n977), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT117), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n830), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n1108), .B2(new_n1107), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n983), .A2(new_n993), .B1(new_n823), .B2(new_n809), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT52), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n807), .A2(new_n868), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n279), .B(new_n1113), .C1(G322), .C2(new_n987), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n793), .A2(new_n641), .B1(new_n1085), .B2(G107), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n814), .A2(G283), .B1(new_n799), .B2(G116), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n983), .A2(new_n412), .B1(new_n284), .B2(new_n809), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT51), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n279), .B1(new_n804), .B2(new_n982), .C1(new_n411), .C2(new_n807), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n800), .A2(new_n220), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G87), .B2(new_n1085), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n793), .A2(G50), .B1(new_n814), .B2(new_n223), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1119), .A2(new_n1121), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n790), .B1(new_n1117), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1110), .A2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1105), .A2(new_n783), .B1(new_n1106), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1058), .A2(new_n1068), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n732), .B1(new_n1058), .B2(new_n1068), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(G390));
  NAND3_X1  g0931(.A1(new_n947), .A2(G330), .A3(new_n950), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n964), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n714), .B(new_n856), .C1(new_n693), .C2(new_n702), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n965), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n961), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n959), .A2(new_n960), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n944), .A2(new_n1137), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n752), .A2(new_n715), .A3(new_n857), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n964), .B1(new_n1140), .B2(new_n966), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1133), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n965), .B1(new_n756), .B2(new_n857), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1137), .B1(new_n1144), .B2(new_n964), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n923), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT39), .B1(new_n943), .B2(new_n923), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n778), .A2(new_n857), .A3(new_n1134), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1143), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n484), .A2(G330), .A3(new_n947), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n947), .A2(G330), .A3(new_n857), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n964), .ZN(new_n1155));
  AND4_X1   g0955(.A1(new_n966), .A2(new_n1155), .A3(new_n1140), .A4(new_n1150), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n964), .B1(new_n862), .B2(new_n856), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1144), .B1(new_n1157), .B2(new_n1132), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n971), .B(new_n1153), .C1(new_n1156), .C2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n733), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT118), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1143), .A2(new_n1151), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1140), .A2(new_n966), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n706), .B(new_n856), .C1(new_n776), .C2(new_n777), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n1134), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1132), .B1(new_n1164), .B2(new_n1134), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1144), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1155), .A2(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AND4_X1   g0968(.A1(KEYINPUT99), .A2(new_n752), .A3(KEYINPUT29), .A4(new_n715), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT99), .B1(new_n746), .B2(KEYINPUT29), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n757), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n683), .B(new_n1153), .C1(new_n1172), .C2(new_n483), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1161), .B1(new_n1162), .B2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1152), .A2(new_n1159), .A3(KEYINPUT118), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1160), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n838), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1122), .B1(G283), .B2(new_n812), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n597), .B2(new_n794), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n871), .A2(new_n868), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n274), .B1(new_n807), .B2(new_n489), .C1(new_n652), .C2(new_n809), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n290), .A2(new_n796), .B1(new_n813), .B2(new_n455), .ZN(new_n1183));
  OR4_X1    g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n814), .A2(G150), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT53), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n821), .A2(G125), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT54), .B(G143), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n279), .B1(new_n807), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G132), .B2(new_n810), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n793), .A2(new_n988), .B1(new_n1085), .B2(G50), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n812), .A2(G128), .B1(G159), .B2(new_n799), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1187), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1184), .B1(new_n1186), .B2(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1194), .A2(new_n789), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n830), .B(new_n1195), .C1(new_n411), .C2(new_n865), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1162), .A2(new_n783), .B1(new_n1178), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1177), .A2(new_n1197), .ZN(G378));
  INV_X1    g0998(.A(KEYINPUT119), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n434), .A2(new_n712), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n447), .A2(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n430), .B(new_n1200), .C1(new_n438), .C2(new_n446), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n430), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n446), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n444), .B1(new_n443), .B2(new_n445), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1200), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n447), .A2(new_n1201), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1204), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1199), .B1(new_n1206), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1205), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1204), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(KEYINPUT119), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n838), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n812), .A2(G125), .ZN(new_n1220));
  INV_X1    g1020(.A(G132), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(new_n794), .B2(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n810), .A2(G128), .B1(new_n876), .B2(G137), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n813), .B2(new_n1188), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(G150), .C2(new_n799), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1085), .A2(G159), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G33), .B(G41), .C1(new_n987), .C2(G124), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n279), .A2(G41), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n807), .B2(new_n452), .C1(new_n597), .C2(new_n809), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n981), .B(new_n1233), .C1(G77), .C2(new_n814), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n817), .B2(new_n871), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n796), .A2(new_n259), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n489), .A2(new_n794), .B1(new_n983), .B2(new_n652), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1232), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1241), .B(new_n414), .C1(G33), .C2(G41), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1231), .A2(new_n1239), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n789), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n783), .B(new_n732), .C1(new_n414), .C2(new_n865), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1219), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n962), .A2(new_n968), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1206), .A2(new_n1213), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n906), .A2(new_n913), .A3(new_n914), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n911), .B1(new_n1251), .B2(new_n905), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n341), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT81), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n351), .B1(new_n350), .B2(new_n352), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1252), .B1(new_n1256), .B2(new_n918), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT38), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n923), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n935), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT40), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n706), .B1(new_n952), .B2(new_n944), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1250), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT38), .B1(new_n938), .B2(new_n941), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1257), .B2(KEYINPUT38), .ZN(new_n1266));
  OAI21_X1  g1066(.A(G330), .B1(new_n1266), .B2(new_n951), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n936), .A2(new_n1267), .A3(new_n1218), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1248), .B1(new_n1264), .B2(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1262), .A2(new_n1263), .A3(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1249), .B1(new_n936), .B2(new_n1267), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n969), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1247), .B1(new_n1274), .B2(new_n783), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1173), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1274), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT120), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1269), .B2(new_n1273), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1273), .A2(new_n1279), .ZN(new_n1281));
  OAI21_X1  g1081(.A(KEYINPUT57), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT118), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1174), .A2(new_n1161), .A3(new_n1151), .A4(new_n1143), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1173), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n732), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1275), .B1(new_n1278), .B2(new_n1286), .ZN(G375));
  OAI21_X1  g1087(.A(KEYINPUT121), .B1(new_n1168), .B2(new_n782), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n983), .A2(new_n868), .B1(new_n813), .B2(new_n489), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(G116), .B2(new_n793), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n821), .A2(G303), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n274), .B1(new_n807), .B2(new_n597), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(G283), .B2(new_n810), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1085), .A2(G77), .B1(new_n572), .B2(new_n799), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n983), .A2(new_n1221), .B1(new_n813), .B2(new_n284), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(G50), .B2(new_n799), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n821), .A2(G128), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n279), .B1(new_n807), .B2(new_n412), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n810), .B2(new_n988), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1188), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1236), .B1(new_n793), .B2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1297), .A2(new_n1298), .A3(new_n1300), .A4(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n790), .B1(new_n1295), .B2(new_n1303), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n830), .B(new_n1304), .C1(new_n290), .C2(new_n865), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(new_n1134), .B2(new_n839), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1288), .A2(new_n1306), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1168), .A2(KEYINPUT121), .A3(new_n782), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1159), .A2(new_n1064), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1309), .B1(new_n1310), .B2(new_n1311), .ZN(G381));
  NOR2_X1   g1112(.A1(G387), .A2(G390), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1177), .A2(new_n1197), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n847), .A2(new_n890), .A3(new_n1069), .A4(new_n1103), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT122), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(KEYINPUT122), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1317), .A2(G381), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1313), .A2(new_n1314), .A3(new_n1316), .A4(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1319), .A2(G375), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT123), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1320), .B(new_n1321), .ZN(G407));
  NAND2_X1  g1122(.A1(new_n713), .A2(G213), .ZN(new_n1323));
  OR3_X1    g1123(.A1(G375), .A2(G378), .A3(new_n1323), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(KEYINPUT124), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(G407), .A2(G213), .A3(new_n1325), .ZN(G409));
  INV_X1    g1126(.A(new_n1323), .ZN(new_n1327));
  OAI211_X1 g1127(.A(G378), .B(new_n1275), .C1(new_n1278), .C2(new_n1286), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1274), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1285), .A2(new_n1063), .A3(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n783), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1246), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1314), .B1(new_n1330), .B2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1327), .B1(new_n1328), .B2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1310), .B1(KEYINPUT60), .B2(new_n1159), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1168), .A2(new_n1173), .A3(KEYINPUT60), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n732), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1309), .B1(new_n1335), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n890), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1309), .B(G384), .C1(new_n1335), .C2(new_n1337), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1334), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT63), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G396), .A2(G393), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(G396), .A2(G393), .ZN(new_n1348));
  OAI221_X1 g1148(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .C1(new_n1347), .C2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1348), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(G390), .A2(new_n1350), .A3(new_n1346), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1349), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(G387), .ZN(new_n1353));
  INV_X1    g1153(.A(G387), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1354), .A2(new_n1351), .A3(new_n1349), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1353), .A2(new_n1355), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1356), .A2(KEYINPUT61), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1327), .A2(KEYINPUT125), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1339), .A2(new_n1340), .A3(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1327), .A2(G2897), .ZN(new_n1360));
  XOR2_X1   g1160(.A(new_n1360), .B(KEYINPUT126), .Z(new_n1361));
  NAND2_X1  g1161(.A1(new_n1359), .A2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1361), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1339), .A2(new_n1340), .A3(new_n1358), .A4(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1362), .A2(new_n1364), .ZN(new_n1365));
  OR2_X1    g1165(.A1(new_n1334), .A2(new_n1365), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1342), .ZN(new_n1367));
  NAND4_X1  g1167(.A1(new_n1345), .A2(new_n1357), .A3(new_n1366), .A4(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT62), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1334), .A2(new_n1369), .A3(new_n1342), .ZN(new_n1370));
  XNOR2_X1  g1170(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1371), .B1(new_n1334), .B2(new_n1365), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1369), .B1(new_n1334), .B2(new_n1342), .ZN(new_n1373));
  NOR3_X1   g1173(.A1(new_n1370), .A2(new_n1372), .A3(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1356), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1368), .B1(new_n1374), .B2(new_n1375), .ZN(G405));
  NAND2_X1  g1176(.A1(G375), .A2(new_n1314), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1377), .A2(new_n1328), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1378), .A2(new_n1342), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1377), .A2(new_n1328), .A3(new_n1341), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  XNOR2_X1  g1181(.A(new_n1381), .B(new_n1356), .ZN(G402));
endmodule


