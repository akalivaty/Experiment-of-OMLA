//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G116), .ZN(new_n210));
  INV_X1    g0010(.A(G270), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n212), .B(new_n218), .C1(G58), .C2(G232), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G1), .B2(G20), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G1), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n226), .A2(new_n223), .A3(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR3_X1   g0029(.A1(new_n221), .A2(new_n225), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G226), .B(G232), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n211), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  INV_X1    g0040(.A(G50), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n210), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  OAI21_X1  g0047(.A(new_n226), .B1(G41), .B2(G45), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  OAI21_X1  g0054(.A(KEYINPUT66), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n251), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT66), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G222), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G223), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n262), .B1(new_n202), .B2(new_n260), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  OAI211_X1 g0066(.A(G1), .B(G13), .C1(new_n253), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n250), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n267), .A2(new_n248), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G226), .ZN(new_n271));
  AOI21_X1  g0071(.A(G169), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n201), .A2(new_n203), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n223), .A2(G33), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT67), .ZN(new_n279));
  XOR2_X1   g0079(.A(KEYINPUT8), .B(G58), .Z(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n274), .B1(new_n275), .B2(new_n277), .C1(new_n279), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n224), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n285), .A2(new_n223), .A3(G1), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n282), .A2(new_n284), .B1(new_n241), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n284), .B1(new_n226), .B2(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G50), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OR3_X1    g0091(.A1(new_n272), .A2(KEYINPUT68), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT68), .B1(new_n272), .B2(new_n291), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n269), .A2(new_n271), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n290), .B(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n269), .B2(new_n271), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(G190), .B2(new_n294), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT70), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n300), .A2(new_n303), .A3(new_n304), .A4(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n269), .A2(G190), .A3(new_n271), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n294), .B2(new_n301), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n306), .B(new_n307), .C1(new_n309), .C2(new_n299), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n297), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT76), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT17), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n280), .A2(new_n286), .ZN(new_n315));
  INV_X1    g0115(.A(new_n288), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n280), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT16), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n255), .A2(new_n223), .A3(new_n259), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT74), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n251), .A2(KEYINPUT74), .A3(G33), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n256), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n214), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G58), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n214), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n329), .B2(new_n203), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n276), .A2(G159), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n318), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n284), .ZN(new_n334));
  AOI21_X1  g0134(.A(G20), .B1(new_n256), .B2(new_n257), .ZN(new_n335));
  OAI21_X1  g0135(.A(G68), .B1(new_n335), .B2(new_n320), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n320), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n332), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n334), .B1(new_n339), .B2(KEYINPUT16), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n317), .B1(new_n333), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n264), .A2(new_n261), .ZN(new_n342));
  INV_X1    g0142(.A(G226), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G1698), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n256), .A2(new_n342), .A3(new_n257), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G87), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n250), .B1(new_n347), .B2(new_n268), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n270), .A2(G232), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT75), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n301), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n350), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n341), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n312), .A2(new_n313), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n314), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n314), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n341), .B2(new_n358), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n341), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n351), .A2(new_n366), .A3(new_n353), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n355), .A2(new_n295), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(new_n370), .A3(KEYINPUT18), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n341), .B2(new_n369), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n364), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT13), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n258), .B1(new_n256), .B2(new_n257), .ZN(new_n378));
  OAI211_X1 g0178(.A(G226), .B(new_n261), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT71), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n260), .A2(new_n381), .A3(G226), .A4(new_n261), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G97), .ZN(new_n384));
  INV_X1    g0184(.A(G232), .ZN(new_n385));
  AOI211_X1 g0185(.A(new_n385), .B(new_n261), .C1(new_n255), .C2(new_n259), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n250), .B1(new_n388), .B2(new_n268), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n270), .A2(G238), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n376), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n386), .B1(new_n380), .B2(new_n382), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n267), .B1(new_n393), .B2(new_n384), .ZN(new_n394));
  INV_X1    g0194(.A(new_n390), .ZN(new_n395));
  NOR4_X1   g0195(.A1(new_n394), .A2(KEYINPUT13), .A3(new_n395), .A4(new_n250), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n397), .A3(G190), .ZN(new_n398));
  OAI21_X1  g0198(.A(G200), .B1(new_n391), .B2(new_n396), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT11), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n276), .A2(G50), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT72), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n402), .B1(new_n223), .B2(G68), .C1(new_n202), .C2(new_n279), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT73), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(new_n284), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n403), .B2(new_n284), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n407), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT11), .A3(new_n405), .ZN(new_n410));
  INV_X1    g0210(.A(new_n286), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(G68), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT12), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n316), .A2(new_n214), .B1(new_n412), .B2(KEYINPUT12), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n408), .A2(new_n410), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n398), .A2(new_n399), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n311), .A2(new_n375), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n411), .A2(G77), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n316), .A2(new_n202), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n280), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT15), .B(G87), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n278), .B2(new_n424), .ZN(new_n425));
  AOI211_X1 g0225(.A(new_n421), .B(new_n422), .C1(new_n425), .C2(new_n284), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT69), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n260), .A2(G232), .A3(new_n261), .ZN(new_n428));
  INV_X1    g0228(.A(G107), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n428), .B1(new_n429), .B2(new_n260), .C1(new_n263), .C2(new_n215), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n250), .B1(new_n430), .B2(new_n268), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n270), .A2(G244), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n427), .B1(new_n433), .B2(G179), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n431), .A2(KEYINPUT69), .A3(new_n295), .A4(new_n432), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n426), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n366), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(G169), .B1(new_n391), .B2(new_n396), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT14), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n392), .A2(G179), .A3(new_n397), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(G169), .C1(new_n391), .C2(new_n396), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n439), .B1(new_n445), .B2(new_n416), .ZN(new_n446));
  INV_X1    g0246(.A(new_n433), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G190), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(new_n426), .C1(new_n301), .C2(new_n447), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n420), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n226), .A2(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(G264), .A3(new_n267), .ZN(new_n457));
  INV_X1    g0257(.A(G250), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n261), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n217), .A2(G1698), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n256), .A2(new_n459), .A3(new_n257), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G294), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n268), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT84), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n455), .A2(G274), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(G179), .A4(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n457), .A2(new_n464), .A3(new_n467), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT84), .B1(new_n469), .B2(G169), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n295), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT85), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n468), .B(KEYINPUT85), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n256), .A2(new_n257), .A3(new_n223), .A4(G87), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT82), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT22), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(KEYINPUT22), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT82), .ZN(new_n481));
  OR2_X1    g0281(.A1(KEYINPUT22), .A2(G20), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n255), .B2(new_n259), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n479), .A2(new_n481), .B1(new_n483), .B2(G87), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT23), .B1(new_n429), .B2(G20), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n429), .A2(KEYINPUT23), .A3(G20), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n253), .A2(new_n210), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n223), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT83), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n481), .A2(new_n479), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n377), .A2(new_n378), .ZN(new_n494));
  INV_X1    g0294(.A(G87), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n494), .A2(new_n495), .A3(new_n482), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n492), .B(new_n489), .C1(new_n493), .C2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n491), .A2(new_n497), .A3(KEYINPUT24), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  OAI211_X1 g0299(.A(KEYINPUT83), .B(new_n499), .C1(new_n484), .C2(new_n490), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n284), .A3(new_n500), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n284), .B(new_n286), .C1(new_n226), .C2(G33), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT25), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n411), .B2(G107), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n429), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n502), .A2(G107), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n476), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n469), .A2(new_n301), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(G190), .B2(new_n469), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n501), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT86), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n501), .A2(new_n506), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n474), .A3(new_n475), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT86), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n501), .A2(new_n506), .A3(new_n509), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n255), .A2(G303), .A3(new_n259), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n252), .A2(new_n254), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n261), .A2(G264), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n217), .A2(new_n261), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n267), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n455), .A2(new_n268), .A3(new_n211), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT81), .B1(new_n525), .B2(new_n467), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT81), .ZN(new_n527));
  INV_X1    g0327(.A(new_n467), .ZN(new_n528));
  NOR4_X1   g0328(.A1(new_n523), .A2(new_n527), .A3(new_n524), .A4(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(G200), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n411), .A2(G116), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n502), .A2(G116), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G283), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT77), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(new_n223), .C1(G33), .C2(new_n216), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n334), .B1(G20), .B2(new_n210), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT20), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n532), .B(new_n533), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n524), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n518), .A2(new_n522), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n467), .B(new_n542), .C1(new_n543), .C2(new_n267), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n527), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n523), .A2(new_n528), .A3(new_n524), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n530), .B(new_n541), .C1(new_n356), .C2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(G169), .B(new_n540), .C1(new_n526), .C2(new_n529), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT21), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n548), .A2(KEYINPUT21), .A3(G169), .A4(new_n540), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n540), .A2(G179), .A3(new_n546), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n549), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n556));
  INV_X1    g0356(.A(G244), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(G1698), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n260), .A2(KEYINPUT4), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n519), .A2(new_n558), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n556), .A2(new_n559), .A3(new_n562), .A4(new_n535), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n268), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n455), .A2(new_n268), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G257), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n467), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G200), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n277), .A2(new_n202), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT6), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n216), .A2(new_n429), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(new_n206), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n429), .A2(KEYINPUT6), .A3(G97), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n575), .A2(new_n223), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n325), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n320), .B2(new_n319), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n570), .B(new_n576), .C1(new_n578), .C2(new_n429), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(new_n284), .B1(new_n216), .B2(new_n286), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n502), .A2(G97), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n564), .A2(G190), .A3(new_n467), .A4(new_n566), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n568), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n284), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n286), .A2(new_n216), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n581), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n567), .A2(new_n366), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n564), .A2(new_n295), .A3(new_n467), .A4(new_n566), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n519), .A2(new_n223), .A3(G68), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n223), .B1(new_n384), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(G87), .B2(new_n207), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n278), .B2(new_n216), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(KEYINPUT79), .B(new_n592), .C1(new_n278), .C2(new_n216), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n591), .A2(new_n594), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n284), .B1(new_n286), .B2(new_n424), .ZN(new_n600));
  INV_X1    g0400(.A(new_n502), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n424), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n226), .A2(G45), .A3(G274), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n458), .B1(new_n451), .B2(KEYINPUT78), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n604), .B(new_n267), .C1(KEYINPUT78), .C2(new_n451), .ZN(new_n605));
  NOR2_X1   g0405(.A1(G238), .A2(G1698), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n557), .B2(G1698), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n488), .B1(new_n519), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n603), .B(new_n605), .C1(new_n608), .C2(new_n267), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n366), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n609), .A2(G179), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n602), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n609), .A2(new_n356), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n502), .A2(G87), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(G200), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n613), .A2(new_n600), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT80), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT80), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n612), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n555), .A2(new_n590), .A3(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n450), .A2(new_n517), .A3(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n297), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n371), .A2(new_n373), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n446), .A2(new_n418), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n364), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n305), .A2(new_n310), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n624), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT87), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n512), .A2(new_n472), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT87), .A4(new_n554), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n590), .A2(new_n510), .A3(new_n617), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT26), .B1(new_n621), .B2(new_n589), .ZN(new_n639));
  INV_X1    g0439(.A(new_n617), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(new_n587), .A3(new_n588), .A4(new_n586), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n612), .B1(new_n641), .B2(KEYINPUT26), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n450), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n630), .A2(new_n645), .ZN(G369));
  XOR2_X1   g0446(.A(new_n555), .B(KEYINPUT88), .Z(new_n647));
  NOR2_X1   g0447(.A1(new_n285), .A2(G20), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n226), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n541), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n647), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G330), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n633), .A2(new_n635), .A3(new_n656), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n512), .A2(new_n654), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n517), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n513), .B2(new_n655), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n512), .A2(new_n472), .A3(new_n655), .ZN(new_n666));
  INV_X1    g0466(.A(new_n631), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n654), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n517), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(G399));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  INV_X1    g0471(.A(new_n227), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G1), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n222), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n671), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n671), .B2(new_n676), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT28), .Z(new_n681));
  NAND2_X1  g0481(.A1(new_n644), .A2(new_n655), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT92), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT29), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n642), .B1(new_n636), .B2(new_n637), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n654), .B1(new_n686), .B2(new_n639), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT92), .B1(new_n687), .B2(KEYINPUT29), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n589), .A2(new_n617), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n612), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n667), .A2(new_n513), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n637), .B2(new_n692), .ZN(new_n693));
  OR3_X1    g0493(.A1(new_n621), .A2(KEYINPUT26), .A3(new_n589), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n654), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n685), .A2(new_n688), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n622), .A2(new_n511), .A3(new_n516), .A4(new_n655), .ZN(new_n698));
  INV_X1    g0498(.A(new_n566), .ZN(new_n699));
  AOI211_X1 g0499(.A(new_n699), .B(new_n609), .C1(new_n563), .C2(new_n268), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n544), .B2(new_n295), .ZN(new_n702));
  INV_X1    g0502(.A(new_n469), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n546), .A2(KEYINPUT90), .A3(G179), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n700), .A2(new_n702), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n469), .A2(new_n295), .A3(new_n609), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n548), .A2(new_n567), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT91), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n548), .A2(new_n567), .A3(KEYINPUT91), .A4(new_n709), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n707), .A2(new_n708), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n654), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n698), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n697), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n681), .B1(new_n722), .B2(G1), .ZN(G364));
  NAND2_X1  g0523(.A1(new_n648), .A2(G45), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n674), .A2(G1), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n661), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n657), .A2(new_n660), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(G330), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n224), .B1(G20), .B2(new_n366), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n223), .A2(G179), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n356), .A3(G200), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G107), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(G190), .A3(G200), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n735), .B(new_n260), .C1(new_n495), .C2(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT98), .Z(new_n738));
  NOR2_X1   g0538(.A1(G190), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n732), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G159), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT97), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT32), .ZN(new_n744));
  NAND2_X1  g0544(.A1(G20), .A2(G179), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT96), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n356), .A2(G200), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n223), .B1(new_n750), .B2(new_n295), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT99), .Z(new_n752));
  OAI22_X1  g0552(.A1(new_n214), .A2(new_n749), .B1(new_n752), .B2(new_n216), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n747), .A2(new_n356), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(new_n750), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n754), .A2(G50), .B1(new_n756), .B2(G58), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n746), .A2(new_n739), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n202), .B2(new_n758), .ZN(new_n759));
  OR4_X1    g0559(.A1(new_n738), .A2(new_n744), .A3(new_n753), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  INV_X1    g0561(.A(G329), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n751), .A2(new_n761), .B1(new_n740), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  INV_X1    g0564(.A(G322), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n758), .B1(new_n755), .B2(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n763), .B(new_n766), .C1(G283), .C2(new_n734), .ZN(new_n767));
  INV_X1    g0567(.A(new_n736), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n260), .B1(G303), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT100), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n769), .A2(new_n770), .B1(new_n754), .B2(G326), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT101), .B(G317), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT33), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n748), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n767), .A2(new_n771), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n731), .B1(new_n760), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT94), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT95), .Z(new_n780));
  AOI21_X1  g0580(.A(new_n730), .B1(new_n780), .B2(new_n223), .ZN(new_n781));
  INV_X1    g0581(.A(G45), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n677), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n256), .A2(new_n257), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n227), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT93), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n783), .B(new_n786), .C1(new_n243), .C2(new_n782), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n494), .A2(new_n672), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G355), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n787), .B(new_n789), .C1(G116), .C2(new_n227), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n777), .B1(new_n781), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n780), .A2(new_n223), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n726), .B(new_n791), .C1(new_n728), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n729), .A2(new_n793), .ZN(G396));
  INV_X1    g0594(.A(new_n758), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n754), .A2(G137), .B1(new_n795), .B2(G159), .ZN(new_n796));
  INV_X1    g0596(.A(G143), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n797), .B2(new_n755), .C1(new_n275), .C2(new_n749), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT102), .Z(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT34), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n733), .A2(new_n214), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n519), .B1(new_n751), .B2(new_n328), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(G50), .C2(new_n768), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n800), .B(new_n803), .C1(new_n804), .C2(new_n740), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n494), .B1(new_n764), .B2(new_n740), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n210), .A2(new_n758), .B1(new_n755), .B2(new_n761), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(G87), .C2(new_n734), .ZN(new_n808));
  INV_X1    g0608(.A(new_n752), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n809), .A2(G97), .B1(G283), .B2(new_n748), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n754), .A2(G303), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n768), .A2(G107), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n808), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n731), .B1(new_n805), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n779), .A2(new_n730), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n725), .B(new_n814), .C1(new_n202), .C2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT103), .Z(new_n817));
  INV_X1    g0617(.A(new_n780), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n426), .A2(new_n655), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT104), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n436), .A2(new_n820), .A3(new_n437), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n436), .B2(new_n437), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n449), .B(new_n819), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n439), .A2(new_n654), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n817), .B1(new_n818), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n449), .ZN(new_n827));
  INV_X1    g0627(.A(new_n822), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n436), .A2(new_n820), .A3(new_n437), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n644), .A2(new_n655), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n687), .B2(new_n825), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(new_n721), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n725), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n826), .A2(new_n834), .ZN(G384));
  INV_X1    g0635(.A(KEYINPUT35), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n223), .B(new_n224), .C1(new_n575), .C2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n837), .B(G116), .C1(new_n836), .C2(new_n575), .ZN(new_n838));
  XNOR2_X1  g0638(.A(KEYINPUT105), .B(KEYINPUT36), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n201), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n214), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n329), .A2(new_n222), .A3(new_n202), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n285), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n840), .B1(new_n226), .B2(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT106), .Z(new_n846));
  NAND2_X1  g0646(.A1(new_n445), .A2(new_n416), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n416), .A2(new_n654), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(new_n419), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n416), .B(new_n654), .C1(new_n445), .C2(new_n418), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n698), .A2(new_n717), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n825), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT107), .B1(new_n341), .B2(new_n652), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT107), .ZN(new_n857));
  INV_X1    g0657(.A(new_n652), .ZN(new_n858));
  INV_X1    g0658(.A(new_n332), .ZN(new_n859));
  INV_X1    g0659(.A(new_n338), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n860), .B2(new_n336), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n284), .B1(new_n861), .B2(new_n318), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n578), .B2(new_n214), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(new_n318), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n857), .B(new_n858), .C1(new_n864), .C2(new_n317), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n856), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n855), .B1(new_n866), .B2(KEYINPUT108), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n365), .A2(new_n370), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n868), .A3(new_n359), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n867), .B(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT109), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n361), .B2(new_n363), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n359), .A2(new_n314), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n341), .A2(new_n358), .B1(new_n312), .B2(new_n313), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n873), .B(KEYINPUT109), .C1(new_n874), .C2(new_n314), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n872), .A2(new_n625), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n866), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n317), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n339), .A2(KEYINPUT16), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n881), .B2(new_n862), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n370), .B2(new_n858), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n883), .A2(KEYINPUT37), .A3(new_n359), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n869), .B2(new_n855), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n858), .B(new_n882), .C1(new_n364), .C2(new_n374), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT40), .B1(new_n854), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n853), .A2(new_n825), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n885), .A2(new_n886), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n890), .A2(new_n895), .A3(new_n896), .A4(new_n851), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n450), .A2(new_n853), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n898), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n893), .B2(new_n894), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT110), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n847), .A2(new_n654), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n876), .A2(new_n877), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n867), .A2(new_n868), .A3(new_n359), .A4(new_n866), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT108), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(new_n856), .B2(new_n865), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n869), .B1(new_n855), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n892), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n903), .A3(new_n894), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT110), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n885), .B2(new_n886), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT39), .B1(new_n887), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n905), .A2(new_n906), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n821), .A2(new_n822), .A3(new_n654), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n831), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n851), .A3(new_n895), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n374), .A2(new_n652), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n919), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n901), .B(new_n925), .Z(new_n926));
  NAND4_X1  g0726(.A1(new_n450), .A2(new_n685), .A3(new_n688), .A4(new_n696), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n630), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n648), .A2(new_n226), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n846), .B1(new_n929), .B2(new_n930), .ZN(G367));
  INV_X1    g0731(.A(G137), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n260), .B1(new_n932), .B2(new_n740), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n275), .A2(new_n755), .B1(new_n758), .B2(new_n201), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n933), .B(new_n934), .C1(G58), .C2(new_n768), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n809), .A2(G68), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n734), .A2(G77), .ZN(new_n937));
  AOI22_X1  g0737(.A1(G143), .A2(new_n754), .B1(new_n748), .B2(G159), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G303), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n755), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(G317), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n784), .B1(new_n740), .B2(new_n942), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n751), .A2(new_n429), .B1(new_n733), .B2(new_n216), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(G283), .C2(new_n795), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G294), .A2(new_n748), .B1(new_n754), .B2(G311), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT114), .B1(new_n736), .B2(new_n210), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT46), .Z(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n939), .B1(new_n941), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT47), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n725), .B1(new_n951), .B2(new_n730), .ZN(new_n952));
  INV_X1    g0752(.A(new_n786), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n781), .B1(new_n227), .B2(new_n424), .C1(new_n238), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n600), .A2(new_n614), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n654), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n640), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n612), .B2(new_n956), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n952), .B(new_n954), .C1(new_n792), .C2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n724), .A2(G1), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n669), .A2(new_n666), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n589), .A2(new_n655), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n586), .A2(new_n654), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n583), .A2(new_n589), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT44), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n961), .A2(new_n966), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n665), .A2(KEYINPUT113), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n669), .B1(new_n664), .B2(new_n668), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n661), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n722), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n722), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n673), .B(KEYINPUT41), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n960), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n669), .A2(new_n964), .ZN(new_n980));
  XNOR2_X1  g0780(.A(KEYINPUT112), .B(KEYINPUT42), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n964), .A2(new_n513), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n983), .A2(new_n589), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n982), .B1(new_n654), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n958), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n985), .A2(new_n986), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n991), .B2(new_n985), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n665), .A2(new_n966), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n993), .B(new_n994), .Z(new_n995));
  OAI21_X1  g0795(.A(new_n959), .B1(new_n979), .B2(new_n995), .ZN(G387));
  OR2_X1    g0796(.A1(new_n975), .A2(new_n722), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(new_n673), .A3(new_n976), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n953), .B1(new_n235), .B2(G45), .ZN(new_n999));
  INV_X1    g0799(.A(new_n675), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n788), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n281), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT50), .B1(new_n281), .B2(G50), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1002), .A2(new_n1003), .A3(new_n782), .A4(new_n675), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G68), .B2(G77), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n1001), .A2(new_n1005), .B1(G107), .B2(new_n227), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n781), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n664), .A2(new_n792), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n754), .A2(G322), .B1(new_n795), .B2(G303), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n764), .B2(new_n749), .C1(new_n942), .C2(new_n755), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT48), .ZN(new_n1011));
  INV_X1    g0811(.A(G283), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n751), .C1(new_n761), .C2(new_n736), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n740), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(G326), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n519), .B1(new_n734), .B2(G116), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n281), .A2(new_n749), .B1(new_n752), .B2(new_n424), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G50), .A2(new_n756), .B1(new_n795), .B2(G68), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n768), .A2(G77), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n519), .B1(new_n275), .B2(new_n740), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G97), .B2(new_n734), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1021), .B(new_n1026), .C1(G159), .C2(new_n754), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT115), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n731), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1008), .A2(new_n725), .A3(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n975), .A2(new_n960), .B1(new_n1007), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n998), .A2(new_n1031), .ZN(G393));
  NAND3_X1  g0832(.A1(new_n968), .A2(new_n665), .A3(new_n970), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n960), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n665), .B1(new_n968), .B2(new_n970), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n781), .B1(new_n216), .B2(new_n227), .C1(new_n246), .C2(new_n953), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n965), .A2(new_n792), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT116), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n519), .B1(new_n797), .B2(new_n740), .C1(new_n758), .C2(new_n281), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n733), .A2(new_n495), .B1(new_n736), .B2(new_n214), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n201), .B2(new_n749), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT51), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n754), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1048), .A2(new_n275), .B1(new_n755), .B2(new_n741), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n1047), .B2(new_n1049), .C1(new_n202), .C2(new_n752), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n754), .A2(G317), .B1(new_n756), .B2(G311), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  OAI21_X1  g0853(.A(new_n494), .B1(new_n758), .B2(new_n761), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n735), .B1(new_n210), .B2(new_n751), .C1(new_n1012), .C2(new_n736), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(G303), .C2(new_n748), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1053), .B(new_n1056), .C1(new_n765), .C2(new_n740), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n725), .B1(new_n1058), .B2(new_n730), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n1041), .A2(new_n1042), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1037), .B1(new_n1038), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n976), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n673), .C1(new_n973), .C2(new_n976), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1061), .A2(new_n1063), .A3(KEYINPUT117), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(G390));
  NAND3_X1  g0868(.A1(new_n450), .A2(G330), .A3(new_n853), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n630), .A2(new_n927), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT118), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n890), .A2(new_n1071), .A3(G330), .A4(new_n851), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n851), .A2(G330), .A3(new_n825), .A4(new_n853), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(KEYINPUT118), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n849), .A2(new_n850), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n825), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1075), .B1(new_n721), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1072), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n922), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n853), .A2(new_n825), .A3(G330), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1075), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n920), .B1(new_n695), .B2(new_n830), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n851), .A2(new_n720), .A3(G330), .A4(new_n825), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1070), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n906), .B1(new_n922), .B2(new_n851), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n905), .B2(new_n918), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n906), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n887), .B2(new_n879), .C1(new_n1082), .C2(new_n1075), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1088), .A2(new_n1091), .A3(new_n1083), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n922), .A2(new_n851), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1089), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n915), .B1(new_n914), .B2(new_n917), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1093), .B1(new_n1098), .B2(new_n1090), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1086), .B1(new_n1092), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1093), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1083), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1098), .A2(new_n1103), .A3(new_n1090), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1084), .B1(new_n1078), .B2(new_n922), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1102), .B(new_n1104), .C1(new_n1070), .C2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1100), .A2(new_n1106), .A3(new_n673), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT119), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1100), .A2(new_n1106), .A3(KEYINPUT119), .A4(new_n673), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n280), .A2(new_n779), .A3(new_n730), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n818), .B1(new_n905), .B2(new_n918), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n260), .B1(new_n201), .B2(new_n733), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n809), .B2(G159), .ZN(new_n1115));
  OAI21_X1  g0915(.A(KEYINPUT53), .B1(new_n736), .B2(new_n275), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT54), .B(G143), .Z(new_n1117));
  NAND2_X1  g0917(.A1(new_n795), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n756), .A2(G132), .ZN(new_n1119));
  OR3_X1    g0919(.A1(new_n736), .A2(KEYINPUT53), .A3(new_n275), .ZN(new_n1120));
  AND4_X1   g0920(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1016), .A2(G125), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G128), .A2(new_n754), .B1(new_n748), .B2(G137), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1115), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n809), .A2(G77), .B1(G283), .B2(new_n754), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n801), .B(new_n260), .C1(G294), .C2(new_n1016), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n216), .A2(new_n758), .B1(new_n755), .B2(new_n210), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G87), .B2(new_n768), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n749), .A2(new_n429), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1124), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1112), .B(new_n1113), .C1(new_n730), .C2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1132), .A2(new_n726), .B1(new_n1133), .B2(new_n960), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1111), .A2(new_n1134), .ZN(G378));
  OAI21_X1  g0935(.A(new_n311), .B1(new_n291), .B2(new_n652), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT55), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n290), .B(new_n858), .C1(new_n628), .C2(new_n624), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT56), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1137), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1142));
  OR3_X1    g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1141), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n780), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n815), .A2(new_n201), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n424), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n748), .A2(G97), .B1(new_n795), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT121), .Z(new_n1151));
  NAND2_X1  g0951(.A1(new_n756), .A2(G107), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n734), .A2(G58), .ZN(new_n1153));
  AOI21_X1  g0953(.A(G41), .B1(new_n1016), .B2(G283), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1152), .A2(new_n784), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n936), .B(new_n1023), .C1(new_n210), .C2(new_n1048), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1151), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT122), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT58), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(KEYINPUT58), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n754), .A2(G125), .B1(new_n795), .B2(G137), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G150), .B2(new_n809), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n756), .A2(G128), .B1(new_n768), .B2(new_n1117), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT123), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(new_n804), .C2(new_n749), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1169));
  AOI21_X1  g0969(.A(G33), .B1(new_n1016), .B2(G124), .ZN(new_n1170));
  AOI21_X1  g0970(.A(G41), .B1(new_n734), .B2(G159), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(KEYINPUT3), .A2(G33), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G50), .B1(new_n1173), .B2(new_n266), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT120), .Z(new_n1175));
  NAND4_X1  g0975(.A1(new_n1159), .A2(new_n1160), .A3(new_n1172), .A4(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n725), .B1(new_n1176), .B2(new_n730), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1147), .A2(new_n1148), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n658), .B1(new_n889), .B2(new_n897), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n925), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n898), .A2(G330), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1181), .A2(new_n923), .A3(new_n919), .A4(new_n924), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1180), .A2(new_n1146), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1146), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1178), .B1(new_n1185), .B2(new_n1035), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1070), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1100), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n674), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1145), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1180), .A2(new_n1182), .A3(new_n1146), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(KEYINPUT57), .A3(new_n1188), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1186), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(G375));
  NAND2_X1  g0998(.A1(new_n1075), .A2(new_n779), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n809), .A2(G50), .B1(new_n748), .B2(new_n1117), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n754), .A2(G132), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n795), .A2(G150), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n784), .B1(new_n1016), .B2(G128), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n1153), .C1(new_n741), .C2(new_n736), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G137), .B2(new_n756), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n809), .A2(new_n1149), .B1(G294), .B2(new_n754), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n937), .B(new_n494), .C1(new_n940), .C2(new_n740), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n429), .A2(new_n758), .B1(new_n755), .B2(new_n1012), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1207), .B(new_n1210), .C1(new_n216), .C2(new_n736), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n749), .A2(new_n210), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1206), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1213), .A2(new_n730), .B1(new_n214), .B2(new_n815), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1199), .A2(new_n726), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1105), .B2(new_n1035), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1105), .A2(new_n1070), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1217), .A2(new_n978), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1086), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1216), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(G381));
  OR2_X1    g1021(.A1(new_n979), .A2(new_n995), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1222), .A2(new_n959), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(G381), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1107), .A2(new_n1134), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(G375), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G384), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G393), .A2(G396), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(G407));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1226), .B2(new_n653), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(G407), .A2(new_n1231), .ZN(G409));
  AOI21_X1  g1032(.A(new_n1070), .B1(new_n1133), .B2(new_n1086), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1190), .B1(new_n1185), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n673), .A3(new_n1196), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1178), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1195), .B2(new_n960), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(G378), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1195), .A2(new_n978), .A3(new_n1188), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1225), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1230), .A2(G343), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1105), .A2(new_n1070), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1086), .B1(new_n1245), .B2(KEYINPUT60), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n674), .B1(new_n1217), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1216), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT125), .B1(new_n1249), .B2(G384), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1217), .A2(new_n1247), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1105), .A2(KEYINPUT60), .A3(new_n1070), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1251), .A2(new_n1219), .A3(new_n673), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1216), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT125), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1256), .A3(new_n1227), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1249), .A2(G384), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1250), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1242), .A2(new_n1244), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1243), .A2(G2897), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1259), .B(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1240), .B1(new_n1197), .B2(G378), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1264), .B1(new_n1243), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1242), .A2(new_n1268), .A3(new_n1244), .A4(new_n1260), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1262), .A2(new_n1266), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(G393), .A2(G396), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(new_n1228), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT127), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1272), .B(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G390), .A2(G387), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1223), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1223), .A2(new_n1275), .B1(new_n1273), .B2(new_n1272), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1270), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1261), .A2(KEYINPUT63), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1242), .A2(new_n1282), .A3(new_n1244), .A4(new_n1260), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1223), .A2(new_n1275), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1272), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1285), .B1(KEYINPUT127), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1276), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT126), .B1(new_n1265), .B2(new_n1243), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1242), .A2(new_n1290), .A3(new_n1244), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1264), .A3(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1284), .A2(new_n1267), .A3(new_n1288), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1280), .A2(new_n1293), .ZN(G405));
  OAI21_X1  g1094(.A(new_n1238), .B1(new_n1197), .B2(new_n1225), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(new_n1260), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1296), .B(new_n1279), .ZN(G402));
endmodule


