

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735;

  XNOR2_X1 U373 ( .A(n405), .B(n530), .ZN(n558) );
  INV_X1 U374 ( .A(G953), .ZN(n723) );
  NOR2_X2 U375 ( .A1(n731), .A2(KEYINPUT65), .ZN(n594) );
  XNOR2_X2 U376 ( .A(n528), .B(n527), .ZN(n545) );
  INV_X1 U377 ( .A(n714), .ZN(n352) );
  NOR2_X2 U378 ( .A1(n644), .A2(n596), .ZN(n582) );
  XNOR2_X1 U379 ( .A(n555), .B(n402), .ZN(n656) );
  XNOR2_X1 U380 ( .A(n364), .B(G131), .ZN(n477) );
  XNOR2_X1 U381 ( .A(n381), .B(G110), .ZN(n480) );
  XOR2_X1 U382 ( .A(G122), .B(G104), .Z(n460) );
  XOR2_X1 U383 ( .A(G116), .B(G107), .Z(n451) );
  NOR2_X1 U384 ( .A1(n628), .A2(n733), .ZN(n595) );
  INV_X1 U385 ( .A(KEYINPUT66), .ZN(n364) );
  NOR2_X1 U386 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U387 ( .A(n731), .B(KEYINPUT65), .ZN(n390) );
  NOR2_X1 U388 ( .A1(G953), .A2(G237), .ZN(n511) );
  XNOR2_X1 U389 ( .A(G107), .B(G104), .ZN(n481) );
  NOR2_X1 U390 ( .A1(n523), .A2(n611), .ZN(n528) );
  INV_X1 U391 ( .A(KEYINPUT87), .ZN(n525) );
  XNOR2_X1 U392 ( .A(n470), .B(n354), .ZN(n560) );
  NOR2_X1 U393 ( .A1(G902), .A2(n694), .ZN(n470) );
  INV_X1 U394 ( .A(KEYINPUT104), .ZN(n366) );
  NAND2_X1 U395 ( .A1(n658), .A2(n353), .ZN(n655) );
  INV_X1 U396 ( .A(G469), .ZN(n403) );
  XNOR2_X1 U397 ( .A(n439), .B(KEYINPUT68), .ZN(n516) );
  XNOR2_X1 U398 ( .A(n438), .B(n373), .ZN(n439) );
  XNOR2_X1 U399 ( .A(n374), .B(G119), .ZN(n373) );
  XNOR2_X1 U400 ( .A(n490), .B(n413), .ZN(n720) );
  INV_X1 U401 ( .A(n491), .ZN(n413) );
  INV_X1 U402 ( .A(G902), .ZN(n517) );
  XNOR2_X1 U403 ( .A(n477), .B(n476), .ZN(n396) );
  INV_X1 U404 ( .A(G134), .ZN(n476) );
  XNOR2_X1 U405 ( .A(n459), .B(n414), .ZN(n490) );
  INV_X1 U406 ( .A(KEYINPUT10), .ZN(n414) );
  INV_X1 U407 ( .A(n490), .ZN(n385) );
  XNOR2_X1 U408 ( .A(G113), .B(G143), .ZN(n466) );
  INV_X1 U409 ( .A(G101), .ZN(n483) );
  INV_X1 U410 ( .A(n730), .ZN(n417) );
  INV_X1 U411 ( .A(n535), .ZN(n408) );
  INV_X1 U412 ( .A(KEYINPUT72), .ZN(n406) );
  INV_X1 U413 ( .A(KEYINPUT30), .ZN(n518) );
  XNOR2_X1 U414 ( .A(n514), .B(n433), .ZN(n432) );
  XNOR2_X1 U415 ( .A(n513), .B(n512), .ZN(n514) );
  INV_X1 U416 ( .A(KEYINPUT45), .ZN(n419) );
  INV_X1 U417 ( .A(KEYINPUT86), .ZN(n381) );
  INV_X1 U418 ( .A(KEYINPUT16), .ZN(n380) );
  XNOR2_X1 U419 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n494) );
  XOR2_X1 U420 ( .A(KEYINPUT89), .B(KEYINPUT79), .Z(n495) );
  XNOR2_X1 U421 ( .A(G119), .B(G128), .ZN(n492) );
  XOR2_X1 U422 ( .A(KEYINPUT90), .B(G110), .Z(n493) );
  XNOR2_X1 U423 ( .A(n450), .B(n356), .ZN(n370) );
  XNOR2_X1 U424 ( .A(G134), .B(G122), .ZN(n448) );
  XNOR2_X1 U425 ( .A(n425), .B(n709), .ZN(n523) );
  XNOR2_X1 U426 ( .A(n442), .B(n443), .ZN(n425) );
  XNOR2_X1 U427 ( .A(n562), .B(n376), .ZN(n678) );
  XNOR2_X1 U428 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n376) );
  INV_X1 U429 ( .A(KEYINPUT112), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n551), .B(KEYINPUT106), .ZN(n570) );
  NAND2_X1 U431 ( .A1(n388), .A2(n387), .ZN(n386) );
  INV_X1 U432 ( .A(n550), .ZN(n387) );
  NAND2_X1 U433 ( .A1(n363), .A2(n362), .ZN(n581) );
  NOR2_X1 U434 ( .A1(n580), .A2(n358), .ZN(n362) );
  INV_X1 U435 ( .A(n579), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n537), .B(n375), .ZN(n538) );
  XNOR2_X1 U437 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n375) );
  OR2_X1 U438 ( .A1(n588), .A2(n550), .ZN(n537) );
  XNOR2_X1 U439 ( .A(n502), .B(KEYINPUT25), .ZN(n503) );
  NOR2_X1 U440 ( .A1(G902), .A2(n705), .ZN(n504) );
  XNOR2_X1 U441 ( .A(n377), .B(KEYINPUT22), .ZN(n608) );
  NAND2_X1 U442 ( .A1(n372), .A2(n371), .ZN(n377) );
  AND2_X1 U443 ( .A1(n587), .A2(n353), .ZN(n371) );
  INV_X1 U444 ( .A(n601), .ZN(n372) );
  INV_X1 U445 ( .A(KEYINPUT1), .ZN(n402) );
  AND2_X1 U446 ( .A1(n680), .A2(G472), .ZN(n409) );
  NAND2_X1 U447 ( .A1(n703), .A2(G210), .ZN(n422) );
  OR2_X1 U448 ( .A1(G237), .A2(G902), .ZN(n524) );
  XNOR2_X1 U449 ( .A(G137), .B(G116), .ZN(n509) );
  INV_X1 U450 ( .A(KEYINPUT44), .ZN(n423) );
  AND2_X1 U451 ( .A1(n392), .A2(n355), .ZN(n391) );
  INV_X1 U452 ( .A(KEYINPUT3), .ZN(n374) );
  NOR2_X1 U453 ( .A1(n682), .A2(n522), .ZN(n398) );
  XOR2_X1 U454 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n449) );
  INV_X1 U455 ( .A(KEYINPUT4), .ZN(n440) );
  XOR2_X1 U456 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n441) );
  XOR2_X1 U457 ( .A(G146), .B(G125), .Z(n459) );
  XOR2_X1 U458 ( .A(KEYINPUT38), .B(n545), .Z(n646) );
  XNOR2_X1 U459 ( .A(n401), .B(KEYINPUT70), .ZN(n599) );
  OR2_X1 U460 ( .A1(n656), .A2(n655), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n431), .B(n367), .ZN(n600) );
  INV_X1 U462 ( .A(G472), .ZN(n367) );
  XNOR2_X1 U463 ( .A(n384), .B(n469), .ZN(n694) );
  XNOR2_X1 U464 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U465 ( .A(n465), .B(n385), .ZN(n384) );
  XNOR2_X1 U466 ( .A(n515), .B(n487), .ZN(n690) );
  XNOR2_X1 U467 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U468 ( .A1(n352), .A2(n399), .ZN(n680) );
  NOR2_X1 U469 ( .A1(n682), .A2(n400), .ZN(n399) );
  XNOR2_X1 U470 ( .A(n368), .B(KEYINPUT71), .ZN(n546) );
  NAND2_X1 U471 ( .A1(n520), .A2(n521), .ZN(n368) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n521) );
  XNOR2_X1 U473 ( .A(n553), .B(n539), .ZN(n579) );
  XNOR2_X1 U474 ( .A(n560), .B(KEYINPUT99), .ZN(n532) );
  AND2_X1 U475 ( .A1(n561), .A2(n532), .ZN(n559) );
  NOR2_X1 U476 ( .A1(n655), .A2(n508), .ZN(n598) );
  XNOR2_X1 U477 ( .A(n516), .B(n426), .ZN(n709) );
  XNOR2_X1 U478 ( .A(n480), .B(n380), .ZN(n437) );
  XNOR2_X1 U479 ( .A(n415), .B(n720), .ZN(n705) );
  XNOR2_X1 U480 ( .A(n498), .B(n499), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n447), .B(n370), .ZN(n454) );
  XNOR2_X1 U482 ( .A(KEYINPUT108), .B(n575), .ZN(n732) );
  XNOR2_X1 U483 ( .A(n564), .B(n565), .ZN(n735) );
  OR2_X1 U484 ( .A1(n563), .A2(n678), .ZN(n564) );
  XNOR2_X1 U485 ( .A(n404), .B(KEYINPUT40), .ZN(n734) );
  NAND2_X1 U486 ( .A1(n558), .A2(n559), .ZN(n404) );
  XNOR2_X1 U487 ( .A(n570), .B(n365), .ZN(n552) );
  XNOR2_X1 U488 ( .A(n586), .B(KEYINPUT82), .ZN(n424) );
  AND2_X1 U489 ( .A1(n591), .A2(n379), .ZN(n378) );
  NOR2_X1 U490 ( .A1(n563), .A2(n579), .ZN(n634) );
  XNOR2_X1 U491 ( .A(n559), .B(KEYINPUT105), .ZN(n636) );
  XNOR2_X1 U492 ( .A(n361), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U493 ( .A1(n411), .A2(n410), .ZN(n361) );
  XNOR2_X1 U494 ( .A(n412), .B(n359), .ZN(n411) );
  INV_X1 U495 ( .A(KEYINPUT122), .ZN(n427) );
  NAND2_X1 U496 ( .A1(n429), .A2(n410), .ZN(n428) );
  XNOR2_X1 U497 ( .A(n430), .B(n693), .ZN(n429) );
  NAND2_X1 U498 ( .A1(n421), .A2(n410), .ZN(n369) );
  XNOR2_X1 U499 ( .A(n422), .B(n616), .ZN(n421) );
  INV_X1 U500 ( .A(n656), .ZN(n379) );
  XNOR2_X1 U501 ( .A(n507), .B(n506), .ZN(n353) );
  XOR2_X1 U502 ( .A(n458), .B(n457), .Z(n354) );
  AND2_X1 U503 ( .A1(n610), .A2(n619), .ZN(n355) );
  XNOR2_X1 U504 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n356) );
  AND2_X1 U505 ( .A1(n595), .A2(n423), .ZN(n357) );
  AND2_X1 U506 ( .A1(G898), .A2(G953), .ZN(n358) );
  XOR2_X1 U507 ( .A(n618), .B(KEYINPUT62), .Z(n359) );
  XOR2_X1 U508 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n360) );
  INV_X1 U509 ( .A(KEYINPUT2), .ZN(n400) );
  INV_X1 U510 ( .A(n708), .ZN(n410) );
  NAND2_X1 U511 ( .A1(n598), .A2(n408), .ZN(n407) );
  NAND2_X1 U512 ( .A1(n391), .A2(n389), .ZN(n420) );
  NOR2_X1 U513 ( .A1(n697), .A2(n708), .ZN(n382) );
  NAND2_X1 U514 ( .A1(n398), .A2(n352), .ZN(n397) );
  INV_X1 U515 ( .A(n606), .ZN(n388) );
  NAND2_X1 U516 ( .A1(n734), .A2(n735), .ZN(n566) );
  INV_X1 U517 ( .A(n600), .ZN(n661) );
  XNOR2_X1 U518 ( .A(n600), .B(n366), .ZN(n534) );
  XNOR2_X1 U519 ( .A(n369), .B(n360), .ZN(G51) );
  NOR2_X1 U520 ( .A1(n636), .A2(n386), .ZN(n551) );
  NAND2_X1 U521 ( .A1(n617), .A2(n517), .ZN(n431) );
  XNOR2_X1 U522 ( .A(n515), .B(n432), .ZN(n617) );
  XNOR2_X2 U523 ( .A(n581), .B(KEYINPUT0), .ZN(n601) );
  AND2_X1 U524 ( .A1(n590), .A2(n378), .ZN(n593) );
  XNOR2_X1 U525 ( .A(n436), .B(n437), .ZN(n426) );
  XNOR2_X1 U526 ( .A(n382), .B(n698), .ZN(G60) );
  NAND2_X1 U527 ( .A1(n357), .A2(n390), .ZN(n389) );
  XNOR2_X1 U528 ( .A(n383), .B(KEYINPUT107), .ZN(n571) );
  NAND2_X1 U529 ( .A1(n570), .A2(n645), .ZN(n383) );
  AND2_X1 U530 ( .A1(n732), .A2(n417), .ZN(n416) );
  NAND2_X1 U531 ( .A1(n393), .A2(KEYINPUT44), .ZN(n392) );
  NAND2_X1 U532 ( .A1(n595), .A2(n594), .ZN(n393) );
  NAND2_X2 U533 ( .A1(n395), .A2(n394), .ZN(n515) );
  NAND2_X1 U534 ( .A1(n719), .A2(G146), .ZN(n394) );
  OR2_X2 U535 ( .A1(n719), .A2(G146), .ZN(n395) );
  XNOR2_X2 U536 ( .A(n478), .B(n396), .ZN(n719) );
  XNOR2_X2 U537 ( .A(n452), .B(n440), .ZN(n478) );
  NAND2_X2 U538 ( .A1(n397), .A2(n614), .ZN(n615) );
  AND2_X4 U539 ( .A1(n615), .A2(n680), .ZN(n703) );
  XNOR2_X2 U540 ( .A(n488), .B(n403), .ZN(n555) );
  NAND2_X1 U541 ( .A1(n546), .A2(n646), .ZN(n405) );
  NAND2_X1 U542 ( .A1(n409), .A2(n615), .ZN(n412) );
  NAND2_X1 U543 ( .A1(n418), .A2(n416), .ZN(n682) );
  XNOR2_X1 U544 ( .A(n569), .B(KEYINPUT48), .ZN(n418) );
  XNOR2_X2 U545 ( .A(n420), .B(n419), .ZN(n714) );
  XNOR2_X2 U546 ( .A(n585), .B(n424), .ZN(n731) );
  XNOR2_X1 U547 ( .A(n428), .B(n427), .ZN(G54) );
  NAND2_X1 U548 ( .A1(n703), .A2(G469), .ZN(n430) );
  INV_X1 U549 ( .A(n516), .ZN(n433) );
  XNOR2_X1 U550 ( .A(n459), .B(n435), .ZN(n443) );
  NOR2_X2 U551 ( .A1(n690), .A2(G902), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n478), .B(n441), .ZN(n442) );
  NAND2_X1 U553 ( .A1(n534), .A2(n645), .ZN(n519) );
  XNOR2_X1 U554 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n434) );
  AND2_X1 U555 ( .A1(G224), .A2(n723), .ZN(n435) );
  XNOR2_X1 U556 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U557 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n529), .B(KEYINPUT83), .ZN(n530) );
  XNOR2_X1 U560 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U561 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U562 ( .A1(G952), .A2(n723), .ZN(n708) );
  XOR2_X1 U563 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n445) );
  XNOR2_X1 U564 ( .A(n451), .B(n460), .ZN(n436) );
  XNOR2_X1 U565 ( .A(G113), .B(G101), .ZN(n438) );
  XOR2_X2 U566 ( .A(G143), .B(G128), .Z(n452) );
  XNOR2_X1 U567 ( .A(n523), .B(KEYINPUT77), .ZN(n444) );
  XNOR2_X1 U568 ( .A(n445), .B(n444), .ZN(n616) );
  XNOR2_X1 U569 ( .A(KEYINPUT102), .B(G478), .ZN(n456) );
  NAND2_X1 U570 ( .A1(G234), .A2(n723), .ZN(n446) );
  XOR2_X1 U571 ( .A(KEYINPUT8), .B(n446), .Z(n489) );
  NAND2_X1 U572 ( .A1(G217), .A2(n489), .ZN(n447) );
  XNOR2_X1 U573 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U574 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U575 ( .A(n454), .B(n453), .ZN(n699) );
  NOR2_X1 U576 ( .A1(G902), .A2(n699), .ZN(n455) );
  XNOR2_X1 U577 ( .A(n456), .B(n455), .ZN(n561) );
  XOR2_X1 U578 ( .A(KEYINPUT98), .B(KEYINPUT13), .Z(n458) );
  XNOR2_X1 U579 ( .A(KEYINPUT97), .B(G475), .ZN(n457) );
  XNOR2_X1 U580 ( .A(n460), .B(KEYINPUT96), .ZN(n464) );
  XOR2_X1 U581 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n462) );
  XNOR2_X1 U582 ( .A(G140), .B(KEYINPUT11), .ZN(n461) );
  XNOR2_X1 U583 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U584 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U585 ( .A(n466), .B(n477), .ZN(n468) );
  NAND2_X1 U586 ( .A1(G214), .A2(n511), .ZN(n467) );
  NOR2_X1 U587 ( .A1(n561), .A2(n532), .ZN(n629) );
  INV_X1 U588 ( .A(n629), .ZN(n639) );
  XNOR2_X1 U589 ( .A(KEYINPUT103), .B(n639), .ZN(n533) );
  NAND2_X1 U590 ( .A1(G234), .A2(G237), .ZN(n471) );
  XNOR2_X1 U591 ( .A(n471), .B(KEYINPUT14), .ZN(n673) );
  NAND2_X1 U592 ( .A1(G953), .A2(n517), .ZN(n472) );
  NAND2_X1 U593 ( .A1(n673), .A2(n472), .ZN(n474) );
  NOR2_X1 U594 ( .A1(G953), .A2(G952), .ZN(n473) );
  NOR2_X1 U595 ( .A1(n474), .A2(n473), .ZN(n578) );
  NAND2_X1 U596 ( .A1(G953), .A2(G900), .ZN(n475) );
  NAND2_X1 U597 ( .A1(n578), .A2(n475), .ZN(n535) );
  XNOR2_X1 U598 ( .A(G137), .B(G140), .ZN(n479) );
  XNOR2_X1 U599 ( .A(n479), .B(KEYINPUT67), .ZN(n491) );
  XNOR2_X1 U600 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U601 ( .A(n491), .B(n482), .ZN(n486) );
  NAND2_X1 U602 ( .A1(G227), .A2(n723), .ZN(n484) );
  INV_X1 U603 ( .A(n555), .ZN(n508) );
  NAND2_X1 U604 ( .A1(n489), .A2(G221), .ZN(n499) );
  XNOR2_X1 U605 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U606 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U607 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n501) );
  XOR2_X1 U608 ( .A(KEYINPUT15), .B(n517), .Z(n522) );
  NAND2_X1 U609 ( .A1(G234), .A2(n522), .ZN(n500) );
  XNOR2_X1 U610 ( .A(n501), .B(n500), .ZN(n505) );
  NAND2_X1 U611 ( .A1(n505), .A2(G217), .ZN(n502) );
  XNOR2_X2 U612 ( .A(n504), .B(n503), .ZN(n658) );
  XOR2_X1 U613 ( .A(KEYINPUT21), .B(KEYINPUT92), .Z(n507) );
  NAND2_X1 U614 ( .A1(n505), .A2(G221), .ZN(n506) );
  XOR2_X1 U615 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n510) );
  XOR2_X1 U616 ( .A(n510), .B(n509), .Z(n513) );
  NAND2_X1 U617 ( .A1(n511), .A2(G210), .ZN(n512) );
  NAND2_X1 U618 ( .A1(G214), .A2(n524), .ZN(n645) );
  INV_X1 U619 ( .A(n522), .ZN(n611) );
  NAND2_X1 U620 ( .A1(G210), .A2(n524), .ZN(n526) );
  INV_X1 U621 ( .A(KEYINPUT39), .ZN(n529) );
  NAND2_X1 U622 ( .A1(n533), .A2(n558), .ZN(n531) );
  XNOR2_X1 U623 ( .A(n531), .B(KEYINPUT113), .ZN(n730) );
  NOR2_X1 U624 ( .A1(n559), .A2(n533), .ZN(n650) );
  NOR2_X1 U625 ( .A1(KEYINPUT69), .A2(n650), .ZN(n540) );
  INV_X1 U626 ( .A(n534), .ZN(n588) );
  NOR2_X1 U627 ( .A1(n658), .A2(n535), .ZN(n536) );
  NAND2_X1 U628 ( .A1(n353), .A2(n536), .ZN(n550) );
  NAND2_X1 U629 ( .A1(n555), .A2(n538), .ZN(n563) );
  XNOR2_X1 U630 ( .A(KEYINPUT73), .B(KEYINPUT19), .ZN(n539) );
  NAND2_X1 U631 ( .A1(n545), .A2(n645), .ZN(n553) );
  NAND2_X1 U632 ( .A1(n540), .A2(n634), .ZN(n541) );
  XOR2_X1 U633 ( .A(n541), .B(KEYINPUT47), .Z(n544) );
  AND2_X1 U634 ( .A1(KEYINPUT69), .A2(n650), .ZN(n542) );
  NAND2_X1 U635 ( .A1(n542), .A2(n634), .ZN(n543) );
  NAND2_X1 U636 ( .A1(n544), .A2(n543), .ZN(n549) );
  INV_X1 U637 ( .A(n545), .ZN(n573) );
  NOR2_X1 U638 ( .A1(n561), .A2(n560), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n546), .A2(n583), .ZN(n547) );
  NOR2_X1 U640 ( .A1(n573), .A2(n547), .ZN(n632) );
  XNOR2_X1 U641 ( .A(n632), .B(KEYINPUT78), .ZN(n548) );
  NOR2_X1 U642 ( .A1(n549), .A2(n548), .ZN(n557) );
  XNOR2_X1 U643 ( .A(KEYINPUT6), .B(n661), .ZN(n606) );
  NOR2_X1 U644 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U645 ( .A(n554), .B(KEYINPUT36), .ZN(n556) );
  NAND2_X1 U646 ( .A1(n556), .A2(n379), .ZN(n643) );
  NAND2_X1 U647 ( .A1(n557), .A2(n643), .ZN(n568) );
  XOR2_X1 U648 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n565) );
  NAND2_X1 U649 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U650 ( .A1(n561), .A2(n560), .ZN(n648) );
  NOR2_X1 U651 ( .A1(n649), .A2(n648), .ZN(n562) );
  XNOR2_X1 U652 ( .A(n566), .B(KEYINPUT46), .ZN(n567) );
  NAND2_X1 U653 ( .A1(n571), .A2(n656), .ZN(n572) );
  XNOR2_X1 U654 ( .A(n572), .B(KEYINPUT43), .ZN(n574) );
  NAND2_X1 U655 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U656 ( .A1(n599), .A2(n606), .ZN(n577) );
  XNOR2_X1 U657 ( .A(KEYINPUT84), .B(KEYINPUT33), .ZN(n576) );
  XNOR2_X1 U658 ( .A(n577), .B(n576), .ZN(n644) );
  INV_X1 U659 ( .A(n578), .ZN(n580) );
  XNOR2_X1 U660 ( .A(n601), .B(KEYINPUT88), .ZN(n596) );
  XNOR2_X1 U661 ( .A(n582), .B(KEYINPUT34), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U663 ( .A(KEYINPUT74), .B(KEYINPUT35), .ZN(n586) );
  INV_X1 U664 ( .A(n648), .ZN(n587) );
  NOR2_X1 U665 ( .A1(n608), .A2(n658), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n588), .A2(n590), .ZN(n589) );
  NOR2_X1 U667 ( .A1(n379), .A2(n589), .ZN(n628) );
  XNOR2_X1 U668 ( .A(KEYINPUT76), .B(n606), .ZN(n591) );
  XOR2_X1 U669 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n592) );
  XNOR2_X1 U670 ( .A(n593), .B(n592), .ZN(n733) );
  NOR2_X1 U671 ( .A1(n661), .A2(n596), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n622) );
  OR2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n664) );
  NOR2_X1 U674 ( .A1(n664), .A2(n601), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT31), .ZN(n603) );
  XNOR2_X1 U676 ( .A(KEYINPUT94), .B(n603), .ZN(n640) );
  NAND2_X1 U677 ( .A1(n622), .A2(n640), .ZN(n605) );
  INV_X1 U678 ( .A(n650), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n658), .A2(n606), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n656), .A2(n609), .ZN(n619) );
  XOR2_X1 U683 ( .A(KEYINPUT81), .B(n611), .Z(n612) );
  NAND2_X1 U684 ( .A1(n612), .A2(KEYINPUT2), .ZN(n613) );
  XNOR2_X1 U685 ( .A(KEYINPUT64), .B(n613), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n617), .B(KEYINPUT85), .ZN(n618) );
  XNOR2_X1 U687 ( .A(G101), .B(n619), .ZN(G3) );
  NOR2_X1 U688 ( .A1(n636), .A2(n622), .ZN(n620) );
  XOR2_X1 U689 ( .A(KEYINPUT114), .B(n620), .Z(n621) );
  XNOR2_X1 U690 ( .A(G104), .B(n621), .ZN(G6) );
  NOR2_X1 U691 ( .A1(n639), .A2(n622), .ZN(n627) );
  XOR2_X1 U692 ( .A(KEYINPUT116), .B(KEYINPUT27), .Z(n624) );
  XNOR2_X1 U693 ( .A(G107), .B(KEYINPUT26), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U695 ( .A(KEYINPUT115), .B(n625), .ZN(n626) );
  XNOR2_X1 U696 ( .A(n627), .B(n626), .ZN(G9) );
  XOR2_X1 U697 ( .A(G110), .B(n628), .Z(G12) );
  XOR2_X1 U698 ( .A(G128), .B(KEYINPUT29), .Z(n631) );
  NAND2_X1 U699 ( .A1(n634), .A2(n629), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n631), .B(n630), .ZN(G30) );
  XOR2_X1 U701 ( .A(G143), .B(n632), .Z(G45) );
  INV_X1 U702 ( .A(n636), .ZN(n633) );
  NAND2_X1 U703 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n635), .B(G146), .ZN(G48) );
  NOR2_X1 U705 ( .A1(n640), .A2(n636), .ZN(n638) );
  XNOR2_X1 U706 ( .A(G113), .B(KEYINPUT117), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n638), .B(n637), .ZN(G15) );
  NOR2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U709 ( .A(G116), .B(n641), .Z(G18) );
  XOR2_X1 U710 ( .A(G125), .B(KEYINPUT37), .Z(n642) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(G27) );
  XNOR2_X1 U712 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n672) );
  BUF_X1 U713 ( .A(n644), .Z(n677) );
  NOR2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n652) );
  NOR2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U717 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U718 ( .A1(n677), .A2(n653), .ZN(n654) );
  XOR2_X1 U719 ( .A(KEYINPUT118), .B(n654), .Z(n670) );
  NAND2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U721 ( .A(n657), .B(KEYINPUT50), .ZN(n663) );
  NOR2_X1 U722 ( .A1(n658), .A2(n353), .ZN(n659) );
  XOR2_X1 U723 ( .A(KEYINPUT49), .B(n659), .Z(n660) );
  NOR2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n665) );
  NAND2_X1 U726 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U727 ( .A(KEYINPUT51), .B(n666), .Z(n668) );
  INV_X1 U728 ( .A(n678), .ZN(n667) );
  NAND2_X1 U729 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U730 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U731 ( .A(n672), .B(n671), .ZN(n675) );
  NAND2_X1 U732 ( .A1(G952), .A2(n673), .ZN(n674) );
  NOR2_X1 U733 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U734 ( .A1(G953), .A2(n676), .ZN(n688) );
  NOR2_X1 U735 ( .A1(n678), .A2(n677), .ZN(n686) );
  NAND2_X1 U736 ( .A1(n714), .A2(n400), .ZN(n679) );
  XNOR2_X1 U737 ( .A(n679), .B(KEYINPUT80), .ZN(n681) );
  NAND2_X1 U738 ( .A1(n681), .A2(n680), .ZN(n684) );
  INV_X1 U739 ( .A(n682), .ZN(n721) );
  NOR2_X1 U740 ( .A1(n721), .A2(KEYINPUT2), .ZN(n683) );
  NOR2_X1 U741 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U742 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U743 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U744 ( .A(KEYINPUT53), .B(n689), .Z(G75) );
  XOR2_X1 U745 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n692) );
  XNOR2_X1 U746 ( .A(n690), .B(KEYINPUT121), .ZN(n691) );
  XNOR2_X1 U747 ( .A(n692), .B(n691), .ZN(n693) );
  NAND2_X1 U748 ( .A1(n703), .A2(G475), .ZN(n696) );
  XNOR2_X1 U749 ( .A(n694), .B(n434), .ZN(n695) );
  XNOR2_X1 U750 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n698) );
  XOR2_X1 U751 ( .A(n699), .B(KEYINPUT125), .Z(n701) );
  NAND2_X1 U752 ( .A1(n703), .A2(G478), .ZN(n700) );
  XNOR2_X1 U753 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U754 ( .A1(n708), .A2(n702), .ZN(G63) );
  NAND2_X1 U755 ( .A1(n703), .A2(G217), .ZN(n704) );
  XNOR2_X1 U756 ( .A(n704), .B(KEYINPUT126), .ZN(n706) );
  XNOR2_X1 U757 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U758 ( .A1(n708), .A2(n707), .ZN(G66) );
  INV_X1 U759 ( .A(G898), .ZN(n713) );
  NAND2_X1 U760 ( .A1(n713), .A2(G953), .ZN(n710) );
  NAND2_X1 U761 ( .A1(n710), .A2(n709), .ZN(n718) );
  NAND2_X1 U762 ( .A1(G953), .A2(G224), .ZN(n711) );
  XOR2_X1 U763 ( .A(KEYINPUT61), .B(n711), .Z(n712) );
  NOR2_X1 U764 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U765 ( .A1(G953), .A2(n714), .ZN(n715) );
  NOR2_X1 U766 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(G69) );
  XNOR2_X1 U768 ( .A(n719), .B(n720), .ZN(n725) );
  INV_X1 U769 ( .A(n725), .ZN(n722) );
  XOR2_X1 U770 ( .A(n722), .B(n721), .Z(n724) );
  NAND2_X1 U771 ( .A1(n724), .A2(n723), .ZN(n729) );
  XOR2_X1 U772 ( .A(G227), .B(n725), .Z(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n727), .A2(G953), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n729), .A2(n728), .ZN(G72) );
  XOR2_X1 U776 ( .A(G134), .B(n730), .Z(G36) );
  XOR2_X1 U777 ( .A(n731), .B(G122), .Z(G24) );
  XNOR2_X1 U778 ( .A(G140), .B(n732), .ZN(G42) );
  XOR2_X1 U779 ( .A(G119), .B(n733), .Z(G21) );
  XNOR2_X1 U780 ( .A(G131), .B(n734), .ZN(G33) );
  XNOR2_X1 U781 ( .A(G137), .B(n735), .ZN(G39) );
endmodule

