//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT66), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(new_n465), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n461), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT71), .ZN(G160));
  NAND2_X1  g054(.A1(new_n466), .A2(KEYINPUT72), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n471), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(KEYINPUT3), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n461), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n488), .A2(new_n470), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  NOR2_X1   g071(.A1(new_n470), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n466), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n484), .A2(new_n461), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n503), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n474), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n502), .B1(new_n506), .B2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  XOR2_X1   g085(.A(KEYINPUT73), .B(G651), .Z(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT74), .A3(G543), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n518), .A2(new_n520), .B1(KEYINPUT5), .B2(new_n517), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n521), .B1(new_n513), .B2(new_n514), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n510), .A2(new_n515), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n511), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT76), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  INV_X1    g106(.A(new_n522), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  INV_X1    g108(.A(new_n515), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n543), .A2(new_n515), .B1(new_n522), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n511), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(G171));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n549), .A2(new_n515), .B1(new_n522), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n511), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G651), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n522), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n515), .B2(new_n564), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G299));
  OR2_X1    g143(.A1(new_n545), .A2(new_n547), .ZN(G301));
  OAI21_X1  g144(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI221_X1 g147(.A(new_n570), .B1(new_n522), .B2(new_n571), .C1(new_n572), .C2(new_n515), .ZN(G288));
  NAND2_X1  g148(.A1(new_n521), .A2(G61), .ZN(new_n574));
  INV_X1    g149(.A(G73), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n517), .ZN(new_n576));
  INV_X1    g151(.A(new_n511), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g153(.A(G86), .B(new_n521), .C1(new_n513), .C2(new_n514), .ZN(new_n579));
  OAI211_X1 g154(.A(G48), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G305));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n582), .A2(new_n515), .B1(new_n522), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n511), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n522), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n515), .B2(KEYINPUT78), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(KEYINPUT78), .B2(new_n515), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n562), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n592), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  OR3_X1    g176(.A1(G168), .A2(KEYINPUT79), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT79), .B1(G168), .B2(new_n601), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n602), .B(new_n603), .C1(G868), .C2(new_n567), .ZN(G297));
  OAI211_X1 g179(.A(new_n602), .B(new_n603), .C1(G868), .C2(new_n567), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n489), .A2(G135), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n491), .A2(G123), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  INV_X1    g189(.A(G111), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n614), .A2(KEYINPUT81), .B1(new_n615), .B2(G2105), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(KEYINPUT81), .B2(new_n614), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n612), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(G2096), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(G2096), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n467), .A2(new_n470), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(new_n473), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(G156));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2430), .Z(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n632), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT84), .Z(new_n644));
  OAI21_X1  g219(.A(G14), .B1(new_n641), .B2(new_n642), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(G401));
  XNOR2_X1  g221(.A(G2084), .B(G2090), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT85), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT86), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  AOI211_X1 g229(.A(new_n648), .B(new_n652), .C1(new_n654), .C2(new_n651), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT18), .ZN(new_n657));
  INV_X1    g232(.A(new_n651), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n655), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT91), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT92), .ZN(new_n679));
  XOR2_X1   g254(.A(G1981), .B(G1986), .Z(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n679), .B(new_n684), .ZN(G229));
  NAND2_X1  g260(.A1(G166), .A2(G16), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G16), .B2(G22), .ZN(new_n687));
  INV_X1    g262(.A(G1971), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(G6), .A2(G16), .ZN(new_n690));
  INV_X1    g265(.A(G305), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G16), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT32), .ZN(new_n693));
  INV_X1    g268(.A(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n687), .A2(new_n688), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G23), .ZN(new_n698));
  INV_X1    g273(.A(G288), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT33), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n689), .A2(new_n695), .A3(new_n696), .A4(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT34), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(KEYINPUT34), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(G25), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n489), .A2(G131), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n491), .A2(G119), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n470), .A2(G107), .ZN(new_n710));
  OAI21_X1  g285(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n708), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT93), .Z(new_n713));
  AOI21_X1  g288(.A(new_n707), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT35), .B(G1991), .Z(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n697), .A2(G24), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n587), .B2(new_n697), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1986), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n716), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n704), .A2(new_n705), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT36), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n697), .A2(G4), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n598), .B2(new_n697), .ZN(new_n725));
  INV_X1    g300(.A(G1348), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n489), .A2(G140), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n491), .A2(G128), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n470), .A2(G116), .ZN(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n706), .A2(G26), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT95), .B(G2067), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n697), .A2(G19), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n554), .B2(new_n697), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT94), .B(G1341), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n727), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT96), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n706), .A2(G32), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n489), .A2(G141), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT97), .Z(new_n747));
  NAND3_X1  g322(.A1(new_n467), .A2(G105), .A3(new_n470), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  AOI211_X1 g327(.A(new_n749), .B(new_n752), .C1(G129), .C2(new_n491), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n745), .B1(new_n755), .B2(new_n706), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n706), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n706), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G2078), .ZN(new_n761));
  NOR2_X1   g336(.A1(G171), .A2(new_n697), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G5), .B2(new_n697), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n764), .B2(new_n763), .ZN(new_n766));
  OR2_X1    g341(.A1(G29), .A2(G33), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n489), .A2(G139), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n770), .C1(new_n470), .C2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(new_n706), .ZN(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT100), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(G28), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n706), .B1(new_n779), .B2(G28), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n778), .B1(new_n780), .B2(new_n781), .C1(new_n760), .C2(G2078), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n775), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n766), .B(new_n783), .C1(new_n706), .C2(new_n620), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n758), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(G168), .A2(G16), .ZN(new_n786));
  NOR2_X1   g361(.A1(G16), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(KEYINPUT99), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT99), .B2(new_n786), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1966), .ZN(new_n790));
  INV_X1    g365(.A(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(G29), .B1(new_n791), .B2(KEYINPUT24), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(KEYINPUT24), .B2(new_n791), .ZN(new_n793));
  INV_X1    g368(.A(G160), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n706), .ZN(new_n795));
  INV_X1    g370(.A(G2084), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n790), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n706), .A2(G35), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G162), .B2(new_n706), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2090), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n697), .A2(G20), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT23), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n567), .B2(new_n697), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT101), .ZN(new_n807));
  INV_X1    g382(.A(G1956), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n799), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n723), .A2(new_n744), .A3(new_n785), .A4(new_n810), .ZN(G150));
  INV_X1    g386(.A(G150), .ZN(G311));
  INV_X1    g387(.A(KEYINPUT103), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n532), .A2(G93), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT102), .B(G55), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n534), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n511), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n554), .ZN(new_n821));
  INV_X1    g396(.A(new_n819), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n814), .A2(new_n816), .A3(KEYINPUT103), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n817), .A2(new_n819), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n825), .A2(KEYINPUT103), .A3(new_n554), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT38), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n598), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n825), .A2(new_n832), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n620), .B(new_n495), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT104), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n620), .B(G162), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n794), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n712), .B(new_n626), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n491), .A2(G130), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT106), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n489), .A2(G142), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n470), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n845), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT107), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  AOI221_X4 g429(.A(KEYINPUT105), .B1(new_n474), .B2(new_n507), .C1(new_n505), .C2(KEYINPUT4), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n506), .B2(new_n508), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n501), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n732), .B(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(new_n754), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n772), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n844), .B(new_n862), .C1(new_n861), .C2(new_n852), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n854), .A2(new_n861), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n844), .B1(new_n867), .B2(new_n862), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT40), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n865), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(new_n872), .ZN(G395));
  XNOR2_X1  g448(.A(new_n827), .B(new_n608), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n598), .A2(G299), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n592), .A2(new_n595), .A3(new_n597), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n567), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(KEYINPUT41), .B1(new_n876), .B2(new_n567), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n876), .A2(KEYINPUT108), .A3(new_n567), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n875), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n879), .B1(new_n888), .B2(new_n874), .ZN(new_n889));
  XNOR2_X1  g464(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(G288), .B(KEYINPUT109), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G290), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT110), .ZN(new_n894));
  NAND2_X1  g469(.A1(G303), .A2(G305), .ZN(new_n895));
  NAND2_X1  g470(.A1(G166), .A2(new_n691), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n894), .A3(new_n895), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n892), .B(new_n587), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n894), .B1(new_n896), .B2(new_n895), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n891), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G868), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(G868), .B2(new_n825), .ZN(G295));
  OAI21_X1  g481(.A(new_n905), .B1(G868), .B2(new_n825), .ZN(G331));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  INV_X1    g484(.A(new_n827), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT114), .ZN(new_n911));
  NAND3_X1  g486(.A1(G168), .A2(KEYINPUT112), .A3(G171), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT112), .ZN(new_n913));
  NAND2_X1  g488(.A1(G301), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(G171), .A2(KEYINPUT112), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(G286), .A3(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n912), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n827), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n916), .A2(new_n824), .A3(new_n826), .A4(new_n912), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT114), .ZN(new_n921));
  AND4_X1   g496(.A1(new_n878), .A2(new_n917), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT113), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n919), .A2(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n888), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n919), .A2(new_n920), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n876), .A2(KEYINPUT108), .A3(new_n567), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT108), .B1(new_n876), .B2(new_n567), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT41), .B1(new_n929), .B2(new_n875), .ZN(new_n930));
  OAI211_X1 g505(.A(KEYINPUT113), .B(new_n926), .C1(new_n930), .C2(new_n882), .ZN(new_n931));
  AOI211_X1 g506(.A(new_n902), .B(new_n922), .C1(new_n925), .C2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n922), .B1(new_n931), .B2(new_n925), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n864), .B1(new_n933), .B2(new_n903), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT115), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g511(.A(KEYINPUT115), .B(new_n864), .C1(new_n933), .C2(new_n903), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n909), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(new_n903), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n917), .A2(new_n919), .A3(new_n921), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n878), .A2(new_n887), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n884), .A2(new_n885), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n941), .B1(new_n942), .B2(new_n881), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n919), .A2(new_n878), .A3(new_n920), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n946), .B2(new_n902), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n939), .A2(new_n947), .A3(new_n909), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT116), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT116), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n939), .A2(new_n947), .A3(new_n950), .A4(new_n909), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n908), .B1(new_n938), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT43), .B1(new_n936), .B2(new_n937), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n939), .A2(KEYINPUT43), .A3(new_n947), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(KEYINPUT4), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n466), .B2(new_n504), .ZN(new_n959));
  INV_X1    g534(.A(new_n508), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT105), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n506), .A2(new_n856), .A3(new_n508), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n502), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n478), .A2(G40), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n964), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n754), .A2(G1996), .A3(new_n966), .ZN(new_n968));
  XOR2_X1   g543(.A(new_n968), .B(KEYINPUT117), .Z(new_n969));
  XOR2_X1   g544(.A(new_n732), .B(G2067), .Z(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n754), .B2(G1996), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n966), .ZN(new_n972));
  INV_X1    g547(.A(new_n715), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n713), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n732), .A2(G2067), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n967), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n967), .B1(new_n755), .B2(new_n970), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT46), .B1(new_n967), .B2(G1996), .ZN(new_n980));
  OR3_X1    g555(.A1(new_n967), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT47), .Z(new_n983));
  XNOR2_X1  g558(.A(new_n712), .B(new_n973), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n966), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n969), .A2(new_n972), .A3(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n967), .A2(G1986), .A3(G290), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n988));
  XNOR2_X1  g563(.A(new_n987), .B(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n983), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n978), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G305), .A2(G1981), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n578), .A2(new_n694), .A3(new_n579), .A4(new_n580), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n993), .A2(KEYINPUT49), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT49), .B1(new_n993), .B2(new_n994), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n963), .B2(G1384), .ZN(new_n999));
  INV_X1    g574(.A(new_n965), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n858), .A2(KEYINPUT118), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(G8), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1003), .B(G8), .C1(new_n1005), .C2(G288), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1005), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1004), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1006), .A2(KEYINPUT120), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n1006), .B2(KEYINPUT120), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1009), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT119), .ZN(new_n1015));
  NAND3_X1  g590(.A1(G303), .A2(G8), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G166), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(G164), .A2(G1384), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n1000), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n688), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n999), .A2(new_n1027), .A3(new_n1002), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n965), .B1(new_n1021), .B2(KEYINPUT50), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1026), .B1(G2090), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1013), .A2(G8), .A3(new_n1020), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1004), .A2(new_n1005), .A3(new_n699), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n994), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(G8), .A3(new_n1003), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1020), .A2(new_n1031), .A3(G8), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1013), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT45), .B1(new_n999), .B2(new_n1002), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(new_n965), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n858), .A2(KEYINPUT118), .A3(new_n1001), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT118), .B1(new_n858), .B2(new_n1001), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1022), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT121), .A3(new_n1000), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1021), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT45), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1041), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1966), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1030), .A2(G2084), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1017), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT63), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1031), .A2(G8), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1019), .B1(G303), .B2(G8), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n1018), .B2(new_n1015), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1054), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1038), .A2(G168), .A3(new_n1053), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1027), .B1(new_n999), .B2(new_n1002), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1000), .B1(new_n1021), .B2(KEYINPUT50), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2090), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1062), .A2(new_n1063), .B1(new_n688), .B2(new_n1025), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1057), .B1(new_n1064), .B2(new_n1017), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1013), .A2(new_n1065), .A3(new_n1037), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1053), .A2(G168), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1054), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1036), .B1(new_n1059), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G286), .A2(G8), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT124), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1053), .A2(KEYINPUT51), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1071), .B(KEYINPUT125), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT123), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1077), .B(new_n1051), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1075), .B1(new_n1079), .B2(G8), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1047), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n999), .A2(new_n1002), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n965), .B1(new_n1082), .B2(new_n1022), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1083), .B2(KEYINPUT121), .ZN(new_n1084));
  AOI21_X1  g659(.A(G1966), .B1(new_n1084), .B2(new_n1041), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1077), .B1(new_n1085), .B2(new_n1051), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1050), .A2(KEYINPUT123), .A3(new_n1052), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1071), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT51), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1073), .B1(new_n1080), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n567), .B(KEYINPUT57), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n808), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1023), .A2(new_n1024), .A3(new_n1000), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1030), .A2(new_n726), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1003), .A2(G2067), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n876), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1092), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1095), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT58), .B(G1341), .Z(new_n1102));
  NAND2_X1  g677(.A1(new_n1003), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1025), .B2(G1996), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1104), .A2(KEYINPUT59), .A3(new_n554), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT59), .B1(new_n1104), .B2(new_n554), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1100), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(new_n1095), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1095), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(KEYINPUT61), .A3(new_n1100), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1348), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n1115), .B2(new_n1097), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1115), .A2(new_n1097), .A3(new_n1114), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n876), .A2(KEYINPUT122), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n598), .B(KEYINPUT122), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1101), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(G171), .B(KEYINPUT54), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1025), .B2(G2078), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1030), .A2(new_n764), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1124), .A2(G2078), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n964), .B2(KEYINPUT45), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n965), .B(new_n1129), .C1(KEYINPUT45), .C2(new_n964), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1123), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1127), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1123), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1128), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1132), .B(new_n1133), .C1(new_n1048), .C2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1066), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1122), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1069), .B1(new_n1090), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1079), .B2(new_n1071), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1086), .A2(G8), .A3(new_n1087), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1074), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1072), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1143), .A2(KEYINPUT62), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1132), .B1(new_n1048), .B2(new_n1134), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1038), .A2(G171), .A3(new_n1065), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1143), .B2(KEYINPUT62), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1138), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n986), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n587), .B(G1986), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n967), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n992), .B1(new_n1148), .B2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g727(.A1(new_n938), .A2(new_n952), .ZN(new_n1154));
  INV_X1    g728(.A(new_n458), .ZN(new_n1155));
  NOR4_X1   g729(.A1(G401), .A2(new_n1155), .A3(G227), .A4(G229), .ZN(new_n1156));
  OAI21_X1  g730(.A(new_n1156), .B1(new_n865), .B2(new_n868), .ZN(new_n1157));
  NOR2_X1   g731(.A1(new_n1154), .A2(new_n1157), .ZN(G308));
  OAI221_X1 g732(.A(new_n1156), .B1(new_n868), .B2(new_n865), .C1(new_n938), .C2(new_n952), .ZN(G225));
endmodule


