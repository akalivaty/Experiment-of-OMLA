

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786;

  XNOR2_X2 U366 ( .A(n492), .B(G902), .ZN(n535) );
  XOR2_X2 U367 ( .A(KEYINPUT59), .B(n680), .Z(n681) );
  XNOR2_X2 U368 ( .A(n675), .B(KEYINPUT122), .ZN(n676) );
  XOR2_X2 U369 ( .A(KEYINPUT90), .B(n665), .Z(n759) );
  XNOR2_X2 U370 ( .A(n375), .B(n568), .ZN(n757) );
  INV_X1 U371 ( .A(G140), .ZN(n474) );
  NOR2_X1 U372 ( .A1(n674), .A2(G902), .ZN(n399) );
  NAND2_X1 U373 ( .A1(n588), .A2(n587), .ZN(n699) );
  NAND2_X2 U374 ( .A1(n403), .A2(n402), .ZN(n406) );
  NOR2_X2 U375 ( .A1(n729), .A2(n726), .ZN(n624) );
  AND2_X2 U376 ( .A1(n405), .A2(n404), .ZN(n371) );
  NAND2_X2 U377 ( .A1(n413), .A2(KEYINPUT65), .ZN(n412) );
  INV_X2 U378 ( .A(n605), .ZN(n606) );
  XNOR2_X2 U379 ( .A(n516), .B(n515), .ZN(n741) );
  NAND2_X2 U380 ( .A1(n465), .A2(n606), .ZN(n516) );
  NOR2_X2 U381 ( .A1(n741), .A2(n583), .ZN(n546) );
  XNOR2_X1 U382 ( .A(n394), .B(n393), .ZN(n650) );
  NOR2_X1 U383 ( .A1(n590), .A2(n410), .ZN(n439) );
  OR2_X1 U384 ( .A1(n644), .A2(n395), .ZN(n394) );
  NOR2_X1 U385 ( .A1(n699), .A2(n631), .ZN(n632) );
  NAND2_X1 U386 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U387 ( .A1(n397), .A2(n618), .ZN(n619) );
  NAND2_X1 U388 ( .A1(n434), .A2(n352), .ZN(n397) );
  XNOR2_X1 U389 ( .A(n640), .B(n382), .ZN(n724) );
  XNOR2_X1 U390 ( .A(n558), .B(n557), .ZN(n587) );
  NAND2_X1 U391 ( .A1(n751), .A2(G469), .ZN(n422) );
  XNOR2_X1 U392 ( .A(n554), .B(n345), .ZN(n556) );
  XNOR2_X1 U393 ( .A(n555), .B(n553), .ZN(n345) );
  XNOR2_X1 U394 ( .A(n539), .B(KEYINPUT79), .ZN(n540) );
  XNOR2_X1 U395 ( .A(n474), .B(G137), .ZN(n483) );
  INV_X1 U396 ( .A(n370), .ZN(n343) );
  NOR2_X1 U397 ( .A1(n440), .A2(n343), .ZN(n436) );
  INV_X1 U398 ( .A(n344), .ZN(n442) );
  NOR2_X1 U399 ( .A1(n666), .A2(KEYINPUT87), .ZN(n344) );
  XNOR2_X2 U400 ( .A(n451), .B(n450), .ZN(n574) );
  NAND2_X1 U401 ( .A1(n668), .A2(n650), .ZN(n651) );
  NAND2_X1 U402 ( .A1(n424), .A2(n368), .ZN(n668) );
  XNOR2_X1 U403 ( .A(n346), .B(n634), .ZN(n652) );
  NAND2_X1 U404 ( .A1(n783), .A2(n785), .ZN(n346) );
  XNOR2_X2 U405 ( .A(n347), .B(KEYINPUT35), .ZN(n666) );
  NAND2_X1 U406 ( .A1(n571), .A2(n396), .ZN(n347) );
  BUF_X1 U407 ( .A(n666), .Z(n348) );
  INV_X1 U408 ( .A(n454), .ZN(n349) );
  NAND2_X1 U409 ( .A1(n414), .A2(n412), .ZN(n364) );
  XNOR2_X1 U410 ( .A(n645), .B(n540), .ZN(n635) );
  INV_X1 U411 ( .A(KEYINPUT15), .ZN(n492) );
  NAND2_X1 U412 ( .A1(n419), .A2(n418), .ZN(n417) );
  INV_X1 U413 ( .A(G469), .ZN(n419) );
  INV_X1 U414 ( .A(KEYINPUT0), .ZN(n450) );
  NAND2_X1 U415 ( .A1(n635), .A2(n545), .ZN(n451) );
  OR2_X1 U416 ( .A1(n643), .A2(n388), .ZN(n387) );
  NAND2_X1 U417 ( .A1(n396), .A2(n391), .ZN(n388) );
  AND2_X1 U418 ( .A1(n392), .A2(n390), .ZN(n389) );
  OR2_X1 U419 ( .A1(n396), .A2(n391), .ZN(n390) );
  NAND2_X1 U420 ( .A1(n411), .A2(n444), .ZN(n410) );
  XOR2_X1 U421 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n561) );
  XNOR2_X1 U422 ( .A(G122), .B(KEYINPUT9), .ZN(n560) );
  NOR2_X1 U423 ( .A1(n659), .A2(n468), .ZN(n467) );
  INV_X1 U424 ( .A(KEYINPUT38), .ZN(n382) );
  OR2_X1 U425 ( .A1(n712), .A2(n466), .ZN(n464) );
  XNOR2_X1 U426 ( .A(G134), .B(G131), .ZN(n473) );
  XNOR2_X1 U427 ( .A(n429), .B(n503), .ZN(n532) );
  XNOR2_X1 U428 ( .A(n431), .B(n430), .ZN(n429) );
  INV_X1 U429 ( .A(G101), .ZN(n430) );
  INV_X1 U430 ( .A(KEYINPUT107), .ZN(n612) );
  XNOR2_X1 U431 ( .A(n428), .B(n427), .ZN(n616) );
  XNOR2_X1 U432 ( .A(n385), .B(n384), .ZN(n637) );
  INV_X1 U433 ( .A(KEYINPUT28), .ZN(n384) );
  NAND2_X1 U434 ( .A1(n381), .A2(n353), .ZN(n576) );
  INV_X1 U435 ( .A(n664), .ZN(n453) );
  AND2_X1 U436 ( .A1(n457), .A2(n358), .ZN(n455) );
  OR2_X1 U437 ( .A1(n664), .A2(G210), .ZN(n456) );
  INV_X1 U438 ( .A(KEYINPUT83), .ZN(n391) );
  AND2_X1 U439 ( .A1(n447), .A2(n445), .ZN(n444) );
  NAND2_X1 U440 ( .A1(KEYINPUT87), .A2(n448), .ZN(n445) );
  NAND2_X1 U441 ( .A1(n449), .A2(n448), .ZN(n447) );
  NAND2_X1 U442 ( .A1(G953), .A2(G902), .ZN(n599) );
  NAND2_X1 U443 ( .A1(n389), .A2(n387), .ZN(n395) );
  INV_X1 U444 ( .A(KEYINPUT47), .ZN(n363) );
  INV_X1 U445 ( .A(KEYINPUT76), .ZN(n393) );
  NOR2_X1 U446 ( .A1(n437), .A2(n436), .ZN(n443) );
  XNOR2_X1 U447 ( .A(KEYINPUT82), .B(KEYINPUT91), .ZN(n523) );
  XOR2_X1 U448 ( .A(KEYINPUT18), .B(KEYINPUT89), .Z(n524) );
  XNOR2_X1 U449 ( .A(n518), .B(n517), .ZN(n521) );
  INV_X1 U450 ( .A(KEYINPUT17), .ZN(n517) );
  OR2_X1 U451 ( .A1(G902), .A2(G237), .ZN(n538) );
  XOR2_X1 U452 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n494) );
  NAND2_X1 U453 ( .A1(G902), .A2(G469), .ZN(n421) );
  INV_X1 U454 ( .A(KEYINPUT48), .ZN(n426) );
  XNOR2_X1 U455 ( .A(G119), .B(KEYINPUT3), .ZN(n431) );
  XNOR2_X1 U456 ( .A(G113), .B(G104), .ZN(n553) );
  XOR2_X1 U457 ( .A(G131), .B(G140), .Z(n548) );
  XNOR2_X1 U458 ( .A(G143), .B(G122), .ZN(n547) );
  NAND2_X1 U459 ( .A1(G237), .A2(G234), .ZN(n541) );
  INV_X1 U460 ( .A(KEYINPUT30), .ZN(n427) );
  INV_X1 U461 ( .A(n617), .ZN(n435) );
  XNOR2_X1 U462 ( .A(G146), .B(G137), .ZN(n507) );
  INV_X1 U463 ( .A(KEYINPUT77), .ZN(n506) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n674) );
  AND2_X1 U465 ( .A1(n559), .A2(G221), .ZN(n400) );
  XNOR2_X1 U466 ( .A(G116), .B(G107), .ZN(n563) );
  NOR2_X1 U467 ( .A1(n659), .A2(n657), .ZN(n469) );
  AND2_X1 U468 ( .A1(n664), .A2(G210), .ZN(n458) );
  NOR2_X1 U469 ( .A1(n583), .A2(n718), .ZN(n582) );
  AND2_X1 U470 ( .A1(n623), .A2(n709), .ZN(n573) );
  XNOR2_X1 U471 ( .A(n531), .B(n530), .ZN(n533) );
  XNOR2_X1 U472 ( .A(KEYINPUT81), .B(G146), .ZN(n478) );
  XNOR2_X1 U473 ( .A(n612), .B(KEYINPUT43), .ZN(n613) );
  BUF_X1 U474 ( .A(n702), .Z(n409) );
  INV_X1 U475 ( .A(KEYINPUT108), .ZN(n432) );
  INV_X1 U476 ( .A(n627), .ZN(n408) );
  INV_X1 U477 ( .A(KEYINPUT56), .ZN(n459) );
  NAND2_X1 U478 ( .A1(n455), .A2(n452), .ZN(n460) );
  NAND2_X1 U479 ( .A1(n454), .A2(n453), .ZN(n452) );
  AND2_X1 U480 ( .A1(n406), .A2(n466), .ZN(n350) );
  NOR2_X1 U481 ( .A1(n643), .A2(n642), .ZN(n351) );
  AND2_X1 U482 ( .A1(n616), .A2(n712), .ZN(n352) );
  INV_X1 U483 ( .A(G902), .ZN(n418) );
  INV_X1 U484 ( .A(KEYINPUT1), .ZN(n407) );
  AND2_X1 U485 ( .A1(n580), .A2(n625), .ZN(n353) );
  AND2_X1 U486 ( .A1(n577), .A2(n368), .ZN(n354) );
  AND2_X1 U487 ( .A1(n368), .A2(n712), .ZN(n355) );
  AND2_X1 U488 ( .A1(n581), .A2(n580), .ZN(n356) );
  INV_X1 U489 ( .A(n686), .ZN(n411) );
  XOR2_X1 U490 ( .A(KEYINPUT68), .B(KEYINPUT22), .Z(n357) );
  AND2_X1 U491 ( .A1(n456), .A2(n759), .ZN(n358) );
  INV_X1 U492 ( .A(KEYINPUT87), .ZN(n572) );
  INV_X1 U493 ( .A(KEYINPUT44), .ZN(n448) );
  NAND2_X1 U494 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n359) );
  INV_X1 U495 ( .A(n657), .ZN(n658) );
  OR2_X1 U496 ( .A1(n469), .A2(n660), .ZN(n360) );
  INV_X1 U497 ( .A(KEYINPUT66), .ZN(n449) );
  AND2_X1 U498 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n361) );
  NAND2_X1 U499 ( .A1(n572), .A2(KEYINPUT44), .ZN(n362) );
  XNOR2_X1 U500 ( .A(n656), .B(n359), .ZN(n470) );
  INV_X1 U501 ( .A(n470), .ZN(n413) );
  XNOR2_X1 U502 ( .A(n363), .B(n639), .ZN(n644) );
  NAND2_X1 U503 ( .A1(n414), .A2(n412), .ZN(n365) );
  BUF_X1 U504 ( .A(n635), .Z(n366) );
  NAND2_X1 U505 ( .A1(n414), .A2(n412), .ZN(n756) );
  XNOR2_X1 U506 ( .A(n576), .B(KEYINPUT67), .ZN(n367) );
  NAND2_X1 U507 ( .A1(n371), .A2(n406), .ZN(n368) );
  NAND2_X1 U508 ( .A1(n371), .A2(n406), .ZN(n398) );
  INV_X1 U509 ( .A(n579), .ZN(n369) );
  NAND2_X1 U510 ( .A1(n367), .A2(n579), .ZN(n370) );
  NAND2_X1 U511 ( .A1(n591), .A2(n361), .ZN(n438) );
  NOR2_X1 U512 ( .A1(n697), .A2(n638), .ZN(n639) );
  INV_X1 U513 ( .A(n583), .ZN(n372) );
  AND2_X1 U514 ( .A1(n422), .A2(n373), .ZN(n403) );
  AND2_X1 U515 ( .A1(n421), .A2(n407), .ZN(n373) );
  NAND2_X1 U516 ( .A1(n422), .A2(n421), .ZN(n420) );
  NOR2_X1 U517 ( .A1(n627), .A2(n435), .ZN(n434) );
  INV_X1 U518 ( .A(n413), .ZN(n374) );
  BUF_X1 U519 ( .A(n567), .Z(n375) );
  BUF_X1 U520 ( .A(n661), .Z(n376) );
  BUF_X1 U521 ( .A(n764), .Z(n377) );
  NAND2_X1 U522 ( .A1(n378), .A2(n379), .ZN(n380) );
  NAND2_X1 U523 ( .A1(n398), .A2(n386), .ZN(n378) );
  NAND2_X1 U524 ( .A1(n350), .A2(n371), .ZN(n379) );
  NAND2_X1 U525 ( .A1(n380), .A2(n464), .ZN(n465) );
  NAND2_X1 U526 ( .A1(n381), .A2(n354), .ZN(n578) );
  AND2_X1 U527 ( .A1(n381), .A2(n356), .ZN(n686) );
  XNOR2_X2 U528 ( .A(n575), .B(n357), .ZN(n381) );
  XNOR2_X1 U529 ( .A(n383), .B(n463), .ZN(n462) );
  NAND2_X1 U530 ( .A1(n443), .A2(n446), .ZN(n383) );
  NOR2_X1 U531 ( .A1(n626), .A2(n625), .ZN(n385) );
  AND2_X2 U532 ( .A1(n708), .A2(n709), .ZN(n712) );
  NAND2_X1 U533 ( .A1(n438), .A2(n439), .ZN(n437) );
  OR2_X2 U534 ( .A1(n609), .A2(n699), .ZN(n425) );
  XNOR2_X1 U535 ( .A(n614), .B(n613), .ZN(n615) );
  NAND2_X1 U536 ( .A1(n416), .A2(KEYINPUT1), .ZN(n404) );
  NAND2_X1 U537 ( .A1(n712), .A2(n466), .ZN(n386) );
  NAND2_X1 U538 ( .A1(n643), .A2(KEYINPUT83), .ZN(n392) );
  INV_X1 U539 ( .A(n642), .ZN(n396) );
  NOR2_X1 U540 ( .A1(n397), .A2(n641), .ZN(n433) );
  INV_X1 U541 ( .A(n368), .ZN(n580) );
  NOR2_X1 U542 ( .A1(n368), .A2(n712), .ZN(n713) );
  NOR2_X1 U543 ( .A1(n611), .A2(n368), .ZN(n614) );
  XNOR2_X2 U544 ( .A(n399), .B(n498), .ZN(n708) );
  XNOR2_X1 U545 ( .A(n488), .B(n772), .ZN(n401) );
  INV_X1 U546 ( .A(n416), .ZN(n402) );
  NOR2_X1 U547 ( .A1(n416), .A2(n420), .ZN(n627) );
  NAND2_X1 U548 ( .A1(n420), .A2(KEYINPUT1), .ZN(n405) );
  NAND2_X1 U549 ( .A1(n366), .A2(n408), .ZN(n636) );
  XNOR2_X1 U550 ( .A(n527), .B(n528), .ZN(n534) );
  XNOR2_X1 U551 ( .A(n597), .B(n596), .ZN(n764) );
  AND2_X2 U552 ( .A1(n415), .A2(n360), .ZN(n414) );
  NAND2_X1 U553 ( .A1(n470), .A2(n467), .ZN(n415) );
  NOR2_X1 U554 ( .A1(n751), .A2(n417), .ZN(n416) );
  XNOR2_X2 U555 ( .A(n461), .B(n481), .ZN(n751) );
  NAND2_X1 U556 ( .A1(n365), .A2(G217), .ZN(n677) );
  XNOR2_X1 U557 ( .A(n423), .B(n679), .ZN(G66) );
  NAND2_X1 U558 ( .A1(n678), .A2(n759), .ZN(n423) );
  XNOR2_X1 U559 ( .A(n649), .B(KEYINPUT36), .ZN(n424) );
  INV_X1 U560 ( .A(n626), .ZN(n607) );
  XNOR2_X1 U561 ( .A(n604), .B(KEYINPUT73), .ZN(n626) );
  XNOR2_X2 U562 ( .A(n425), .B(KEYINPUT105), .ZN(n646) );
  XNOR2_X1 U563 ( .A(n653), .B(n426), .ZN(n654) );
  INV_X2 U564 ( .A(G953), .ZN(n776) );
  NAND2_X1 U565 ( .A1(n715), .A2(n723), .ZN(n428) );
  XNOR2_X2 U566 ( .A(n513), .B(G472), .ZN(n715) );
  XNOR2_X1 U567 ( .A(n433), .B(n432), .ZN(n643) );
  NAND2_X1 U568 ( .A1(n784), .A2(n449), .ZN(n440) );
  NAND2_X1 U569 ( .A1(n442), .A2(n441), .ZN(n446) );
  NAND2_X1 U570 ( .A1(n666), .A2(n362), .ZN(n441) );
  NAND2_X1 U571 ( .A1(n693), .A2(n784), .ZN(n591) );
  XNOR2_X2 U572 ( .A(n629), .B(KEYINPUT42), .ZN(n785) );
  NOR2_X2 U573 ( .A1(n648), .A2(n647), .ZN(n649) );
  INV_X1 U574 ( .A(n574), .ZN(n583) );
  INV_X1 U575 ( .A(n365), .ZN(n454) );
  NAND2_X1 U576 ( .A1(n364), .A2(n458), .ZN(n457) );
  XNOR2_X1 U577 ( .A(n460), .B(n459), .ZN(G51) );
  XNOR2_X1 U578 ( .A(n461), .B(n773), .ZN(n778) );
  XNOR2_X2 U579 ( .A(n511), .B(n475), .ZN(n461) );
  NAND2_X1 U580 ( .A1(n462), .A2(n595), .ZN(n597) );
  INV_X1 U581 ( .A(KEYINPUT86), .ZN(n463) );
  INV_X1 U582 ( .A(KEYINPUT103), .ZN(n466) );
  NAND2_X1 U583 ( .A1(n374), .A2(n658), .ZN(n747) );
  NAND2_X1 U584 ( .A1(n658), .A2(n660), .ZN(n468) );
  XNOR2_X2 U585 ( .A(n578), .B(KEYINPUT32), .ZN(n784) );
  XOR2_X1 U586 ( .A(n496), .B(n495), .Z(n471) );
  INV_X1 U587 ( .A(n519), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U590 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U591 ( .A(n497), .B(n471), .ZN(n498) );
  XNOR2_X1 U592 ( .A(n529), .B(G122), .ZN(n531) );
  XNOR2_X2 U593 ( .A(G143), .B(KEYINPUT64), .ZN(n472) );
  XNOR2_X2 U594 ( .A(n472), .B(G128), .ZN(n567) );
  XNOR2_X2 U595 ( .A(n567), .B(KEYINPUT4), .ZN(n526) );
  XNOR2_X2 U596 ( .A(n526), .B(n473), .ZN(n511) );
  INV_X1 U597 ( .A(n483), .ZN(n475) );
  XNOR2_X1 U598 ( .A(G110), .B(G107), .ZN(n476) );
  XNOR2_X1 U599 ( .A(n476), .B(G104), .ZN(n530) );
  NAND2_X1 U600 ( .A1(n776), .A2(G227), .ZN(n477) );
  XNOR2_X1 U601 ( .A(n477), .B(G101), .ZN(n479) );
  XNOR2_X1 U602 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U603 ( .A(n530), .B(n480), .ZN(n481) );
  XNOR2_X1 U604 ( .A(KEYINPUT72), .B(KEYINPUT10), .ZN(n482) );
  XNOR2_X2 U605 ( .A(G125), .B(G146), .ZN(n519) );
  XOR2_X1 U606 ( .A(n482), .B(n519), .Z(n772) );
  XNOR2_X1 U607 ( .A(n483), .B(KEYINPUT23), .ZN(n487) );
  XOR2_X1 U608 ( .A(KEYINPUT24), .B(G110), .Z(n485) );
  XNOR2_X1 U609 ( .A(G128), .B(G119), .ZN(n484) );
  XNOR2_X1 U610 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U611 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U612 ( .A(KEYINPUT8), .B(KEYINPUT71), .Z(n490) );
  NAND2_X1 U613 ( .A1(G234), .A2(n776), .ZN(n489) );
  XNOR2_X1 U614 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U615 ( .A(KEYINPUT84), .B(n491), .Z(n559) );
  INV_X1 U616 ( .A(n535), .ZN(n659) );
  NAND2_X1 U617 ( .A1(G234), .A2(n659), .ZN(n493) );
  XNOR2_X1 U618 ( .A(n494), .B(n493), .ZN(n499) );
  NAND2_X1 U619 ( .A1(G217), .A2(n499), .ZN(n497) );
  XOR2_X1 U620 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n496) );
  XNOR2_X1 U621 ( .A(KEYINPUT94), .B(KEYINPUT96), .ZN(n495) );
  NAND2_X1 U622 ( .A1(n499), .A2(G221), .ZN(n502) );
  XNOR2_X1 U623 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n500) );
  XNOR2_X1 U624 ( .A(n500), .B(KEYINPUT21), .ZN(n501) );
  XNOR2_X1 U625 ( .A(n502), .B(n501), .ZN(n709) );
  XNOR2_X1 U626 ( .A(G116), .B(G113), .ZN(n503) );
  XOR2_X1 U627 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n505) );
  NOR2_X2 U628 ( .A1(G953), .A2(G237), .ZN(n549) );
  NAND2_X1 U629 ( .A1(n549), .A2(G210), .ZN(n504) );
  XNOR2_X1 U630 ( .A(n505), .B(n504), .ZN(n509) );
  XNOR2_X1 U631 ( .A(n532), .B(n510), .ZN(n512) );
  XNOR2_X1 U632 ( .A(n511), .B(n512), .ZN(n669) );
  NAND2_X1 U633 ( .A1(n669), .A2(n418), .ZN(n513) );
  XNOR2_X1 U634 ( .A(n715), .B(KEYINPUT6), .ZN(n605) );
  INV_X1 U635 ( .A(KEYINPUT74), .ZN(n514) );
  XNOR2_X1 U636 ( .A(n514), .B(KEYINPUT33), .ZN(n515) );
  NAND2_X1 U637 ( .A1(G224), .A2(n776), .ZN(n518) );
  XNOR2_X1 U638 ( .A(n522), .B(KEYINPUT92), .ZN(n528) );
  XNOR2_X1 U639 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U640 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U641 ( .A(KEYINPUT75), .B(KEYINPUT16), .Z(n529) );
  XNOR2_X1 U642 ( .A(n533), .B(n532), .ZN(n762) );
  XNOR2_X1 U643 ( .A(n534), .B(n762), .ZN(n661) );
  NOR2_X1 U644 ( .A1(n661), .A2(n535), .ZN(n537) );
  NAND2_X1 U645 ( .A1(G210), .A2(n538), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n537), .B(n536), .ZN(n598) );
  NAND2_X1 U647 ( .A1(G214), .A2(n538), .ZN(n723) );
  NAND2_X1 U648 ( .A1(n598), .A2(n723), .ZN(n645) );
  XNOR2_X1 U649 ( .A(KEYINPUT19), .B(KEYINPUT69), .ZN(n539) );
  XNOR2_X1 U650 ( .A(n541), .B(KEYINPUT93), .ZN(n542) );
  XNOR2_X1 U651 ( .A(KEYINPUT14), .B(n542), .ZN(n738) );
  AND2_X1 U652 ( .A1(n776), .A2(G952), .ZN(n601) );
  NOR2_X1 U653 ( .A1(G898), .A2(n599), .ZN(n543) );
  NOR2_X1 U654 ( .A1(n601), .A2(n543), .ZN(n544) );
  NOR2_X1 U655 ( .A1(n738), .A2(n544), .ZN(n545) );
  XNOR2_X1 U656 ( .A(n546), .B(KEYINPUT34), .ZN(n571) );
  XNOR2_X1 U657 ( .A(n548), .B(n547), .ZN(n555) );
  XOR2_X1 U658 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n551) );
  NAND2_X1 U659 ( .A1(n549), .A2(G214), .ZN(n550) );
  XNOR2_X1 U660 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U661 ( .A(n552), .B(KEYINPUT11), .Z(n554) );
  XNOR2_X1 U662 ( .A(n772), .B(n556), .ZN(n680) );
  NAND2_X1 U663 ( .A1(n680), .A2(n418), .ZN(n558) );
  XOR2_X1 U664 ( .A(KEYINPUT13), .B(G475), .Z(n557) );
  NAND2_X1 U665 ( .A1(G217), .A2(n559), .ZN(n566) );
  XNOR2_X1 U666 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U667 ( .A(n562), .B(G134), .Z(n564) );
  XNOR2_X1 U668 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U669 ( .A(n566), .B(n565), .ZN(n568) );
  NAND2_X1 U670 ( .A1(n757), .A2(n418), .ZN(n570) );
  XNOR2_X1 U671 ( .A(G478), .B(KEYINPUT102), .ZN(n569) );
  XNOR2_X1 U672 ( .A(n570), .B(n569), .ZN(n586) );
  NAND2_X1 U673 ( .A1(n587), .A2(n586), .ZN(n642) );
  NOR2_X1 U674 ( .A1(n586), .A2(n587), .ZN(n623) );
  INV_X1 U675 ( .A(n708), .ZN(n579) );
  NAND2_X1 U676 ( .A1(n367), .A2(n579), .ZN(n693) );
  NOR2_X1 U677 ( .A1(n606), .A2(n369), .ZN(n577) );
  NOR2_X1 U678 ( .A1(n606), .A2(n579), .ZN(n581) );
  NAND2_X1 U679 ( .A1(n355), .A2(n715), .ZN(n718) );
  XNOR2_X1 U680 ( .A(n582), .B(KEYINPUT31), .ZN(n702) );
  INV_X1 U681 ( .A(n715), .ZN(n625) );
  NAND2_X1 U682 ( .A1(n712), .A2(n625), .ZN(n584) );
  NOR2_X1 U683 ( .A1(n584), .A2(n627), .ZN(n585) );
  NAND2_X1 U684 ( .A1(n372), .A2(n585), .ZN(n690) );
  NAND2_X1 U685 ( .A1(n702), .A2(n690), .ZN(n589) );
  INV_X1 U686 ( .A(n586), .ZN(n588) );
  OR2_X1 U687 ( .A1(n588), .A2(n587), .ZN(n703) );
  NAND2_X1 U688 ( .A1(n703), .A2(n699), .ZN(n728) );
  AND2_X1 U689 ( .A1(n589), .A2(n728), .ZN(n590) );
  BUF_X1 U690 ( .A(n591), .Z(n592) );
  NOR2_X1 U691 ( .A1(n592), .A2(KEYINPUT44), .ZN(n594) );
  INV_X1 U692 ( .A(n348), .ZN(n593) );
  NAND2_X1 U693 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U694 ( .A(KEYINPUT45), .ZN(n596) );
  BUF_X1 U695 ( .A(n598), .Z(n640) );
  NOR2_X1 U696 ( .A1(G900), .A2(n599), .ZN(n600) );
  NOR2_X1 U697 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U698 ( .A1(n602), .A2(n738), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n617), .A2(n709), .ZN(n603) );
  NOR2_X1 U700 ( .A1(n708), .A2(n603), .ZN(n604) );
  NAND2_X1 U701 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U702 ( .A(n608), .B(KEYINPUT104), .ZN(n609) );
  NAND2_X1 U703 ( .A1(n646), .A2(n723), .ZN(n610) );
  XNOR2_X1 U704 ( .A(KEYINPUT106), .B(n610), .ZN(n611) );
  NOR2_X1 U705 ( .A1(n640), .A2(n615), .ZN(n707) );
  INV_X1 U706 ( .A(n724), .ZN(n618) );
  XNOR2_X1 U707 ( .A(KEYINPUT39), .B(n619), .ZN(n631) );
  INV_X1 U708 ( .A(n631), .ZN(n621) );
  INV_X1 U709 ( .A(n703), .ZN(n620) );
  NAND2_X1 U710 ( .A1(n621), .A2(n620), .ZN(n706) );
  INV_X1 U711 ( .A(n706), .ZN(n622) );
  OR2_X1 U712 ( .A1(n707), .A2(n622), .ZN(n655) );
  XOR2_X1 U713 ( .A(KEYINPUT46), .B(KEYINPUT85), .Z(n634) );
  NAND2_X1 U714 ( .A1(n724), .A2(n723), .ZN(n729) );
  INV_X1 U715 ( .A(n623), .ZN(n726) );
  XOR2_X1 U716 ( .A(KEYINPUT41), .B(n624), .Z(n721) );
  NOR2_X1 U717 ( .A1(n637), .A2(n627), .ZN(n628) );
  NAND2_X1 U718 ( .A1(n721), .A2(n628), .ZN(n629) );
  XOR2_X1 U719 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n630) );
  XNOR2_X1 U720 ( .A(KEYINPUT40), .B(n630), .ZN(n633) );
  XOR2_X1 U721 ( .A(n633), .B(n632), .Z(n783) );
  OR2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n697) );
  NAND2_X1 U723 ( .A1(KEYINPUT70), .A2(n728), .ZN(n638) );
  INV_X1 U724 ( .A(n640), .ZN(n641) );
  BUF_X1 U725 ( .A(n645), .Z(n648) );
  XNOR2_X1 U726 ( .A(KEYINPUT111), .B(n646), .ZN(n647) );
  NOR2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  OR2_X2 U728 ( .A1(n655), .A2(n654), .ZN(n774) );
  NOR2_X2 U729 ( .A1(n764), .A2(n774), .ZN(n656) );
  NOR2_X1 U730 ( .A1(KEYINPUT2), .A2(KEYINPUT78), .ZN(n657) );
  INV_X1 U731 ( .A(KEYINPUT65), .ZN(n660) );
  XNOR2_X1 U732 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n376), .B(KEYINPUT88), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X1 U735 ( .A1(n776), .A2(G952), .ZN(n665) );
  XOR2_X1 U736 ( .A(n348), .B(G122), .Z(G24) );
  XOR2_X1 U737 ( .A(G125), .B(KEYINPUT37), .Z(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(G27) );
  NAND2_X1 U739 ( .A1(n756), .A2(G472), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n669), .B(KEYINPUT62), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n672), .A2(n759), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n673), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U744 ( .A(KEYINPUT124), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n674), .B(KEYINPUT123), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n364), .A2(G475), .ZN(n682) );
  XNOR2_X1 U748 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n683), .A2(n759), .ZN(n685) );
  XOR2_X1 U750 ( .A(KEYINPUT120), .B(KEYINPUT60), .Z(n684) );
  XNOR2_X1 U751 ( .A(n685), .B(n684), .ZN(G60) );
  XOR2_X1 U752 ( .A(G101), .B(n686), .Z(G3) );
  NOR2_X1 U753 ( .A1(n699), .A2(n690), .ZN(n687) );
  XOR2_X1 U754 ( .A(G104), .B(n687), .Z(G6) );
  XOR2_X1 U755 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n689) );
  XNOR2_X1 U756 ( .A(G107), .B(KEYINPUT112), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n689), .B(n688), .ZN(n692) );
  NOR2_X1 U758 ( .A1(n703), .A2(n690), .ZN(n691) );
  XOR2_X1 U759 ( .A(n692), .B(n691), .Z(G9) );
  XNOR2_X1 U760 ( .A(n370), .B(G110), .ZN(G12) );
  NOR2_X1 U761 ( .A1(n703), .A2(n697), .ZN(n695) );
  XNOR2_X1 U762 ( .A(KEYINPUT113), .B(KEYINPUT29), .ZN(n694) );
  XNOR2_X1 U763 ( .A(n695), .B(n694), .ZN(n696) );
  XOR2_X1 U764 ( .A(G128), .B(n696), .Z(G30) );
  XOR2_X1 U765 ( .A(G143), .B(n351), .Z(G45) );
  NOR2_X1 U766 ( .A1(n699), .A2(n697), .ZN(n698) );
  XOR2_X1 U767 ( .A(G146), .B(n698), .Z(G48) );
  NOR2_X1 U768 ( .A1(n699), .A2(n409), .ZN(n700) );
  XOR2_X1 U769 ( .A(KEYINPUT114), .B(n700), .Z(n701) );
  XNOR2_X1 U770 ( .A(G113), .B(n701), .ZN(G15) );
  NOR2_X1 U771 ( .A1(n703), .A2(n409), .ZN(n705) );
  XNOR2_X1 U772 ( .A(G116), .B(KEYINPUT115), .ZN(n704) );
  XNOR2_X1 U773 ( .A(n705), .B(n704), .ZN(G18) );
  XNOR2_X1 U774 ( .A(G134), .B(n706), .ZN(G36) );
  XOR2_X1 U775 ( .A(G140), .B(n707), .Z(G42) );
  NOR2_X1 U776 ( .A1(n709), .A2(n369), .ZN(n710) );
  XNOR2_X1 U777 ( .A(n710), .B(KEYINPUT116), .ZN(n711) );
  XNOR2_X1 U778 ( .A(n711), .B(KEYINPUT49), .ZN(n717) );
  XNOR2_X1 U779 ( .A(n713), .B(KEYINPUT50), .ZN(n714) );
  NOR2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U782 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U783 ( .A(KEYINPUT51), .B(n720), .ZN(n722) );
  INV_X1 U784 ( .A(n721), .ZN(n740) );
  NOR2_X1 U785 ( .A1(n722), .A2(n740), .ZN(n735) );
  NOR2_X1 U786 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U787 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U788 ( .A(KEYINPUT117), .B(n727), .Z(n732) );
  INV_X1 U789 ( .A(n728), .ZN(n730) );
  NOR2_X1 U790 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U791 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U792 ( .A1(n741), .A2(n733), .ZN(n734) );
  NOR2_X1 U793 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U794 ( .A(n736), .B(KEYINPUT52), .ZN(n737) );
  NOR2_X1 U795 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U796 ( .A1(G952), .A2(n739), .ZN(n743) );
  OR2_X1 U797 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U798 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U799 ( .A(n744), .B(KEYINPUT118), .ZN(n745) );
  NOR2_X1 U800 ( .A1(n745), .A2(G953), .ZN(n746) );
  AND2_X1 U801 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U802 ( .A(n748), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U803 ( .A(n759), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n349), .A2(G469), .ZN(n753) );
  XNOR2_X1 U805 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n749) );
  XNOR2_X1 U806 ( .A(n749), .B(KEYINPUT57), .ZN(n750) );
  XNOR2_X1 U807 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U808 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U809 ( .A1(n755), .A2(n754), .ZN(G54) );
  NAND2_X1 U810 ( .A1(n756), .A2(G478), .ZN(n758) );
  XNOR2_X1 U811 ( .A(n758), .B(n757), .ZN(n760) );
  NAND2_X1 U812 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U813 ( .A(n761), .B(KEYINPUT121), .ZN(G63) );
  INV_X1 U814 ( .A(G898), .ZN(n767) );
  NAND2_X1 U815 ( .A1(n767), .A2(G953), .ZN(n763) );
  NAND2_X1 U816 ( .A1(n763), .A2(n762), .ZN(n771) );
  NOR2_X1 U817 ( .A1(n377), .A2(G953), .ZN(n769) );
  NAND2_X1 U818 ( .A1(G953), .A2(G224), .ZN(n765) );
  XOR2_X1 U819 ( .A(KEYINPUT61), .B(n765), .Z(n766) );
  NOR2_X1 U820 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U821 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U822 ( .A(n771), .B(n770), .ZN(G69) );
  XOR2_X1 U823 ( .A(n772), .B(KEYINPUT125), .Z(n773) );
  XNOR2_X1 U824 ( .A(n778), .B(KEYINPUT126), .ZN(n775) );
  XNOR2_X1 U825 ( .A(n775), .B(n774), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n777), .A2(n776), .ZN(n782) );
  XNOR2_X1 U827 ( .A(G227), .B(n778), .ZN(n779) );
  NAND2_X1 U828 ( .A1(n779), .A2(G900), .ZN(n780) );
  NAND2_X1 U829 ( .A1(n780), .A2(G953), .ZN(n781) );
  NAND2_X1 U830 ( .A1(n782), .A2(n781), .ZN(G72) );
  XNOR2_X1 U831 ( .A(G131), .B(n783), .ZN(G33) );
  XNOR2_X1 U832 ( .A(G119), .B(n784), .ZN(G21) );
  XOR2_X1 U833 ( .A(n785), .B(G137), .Z(n786) );
  XNOR2_X1 U834 ( .A(KEYINPUT127), .B(n786), .ZN(G39) );
endmodule

