

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  XOR2_X1 U321 ( .A(n382), .B(n381), .Z(n289) );
  NOR2_X1 U322 ( .A1(n421), .A2(n420), .ZN(n422) );
  XNOR2_X1 U323 ( .A(n387), .B(n386), .ZN(n388) );
  NOR2_X1 U324 ( .A1(n510), .A2(n424), .ZN(n563) );
  XNOR2_X1 U325 ( .A(n389), .B(n388), .ZN(n391) );
  INV_X1 U326 ( .A(G190GAT), .ZN(n442) );
  XNOR2_X1 U327 ( .A(n392), .B(n569), .ZN(n554) );
  XNOR2_X1 U328 ( .A(n442), .B(KEYINPUT58), .ZN(n443) );
  XNOR2_X1 U329 ( .A(n444), .B(n443), .ZN(G1351GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n291) );
  XNOR2_X1 U331 ( .A(G92GAT), .B(KEYINPUT78), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U333 ( .A(G50GAT), .B(G162GAT), .Z(n319) );
  XOR2_X1 U334 ( .A(n292), .B(n319), .Z(n294) );
  XNOR2_X1 U335 ( .A(G218GAT), .B(G106GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n299) );
  XNOR2_X1 U337 ( .A(G99GAT), .B(G85GAT), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n295), .B(KEYINPUT73), .ZN(n380) );
  XOR2_X1 U339 ( .A(G36GAT), .B(G190GAT), .Z(n346) );
  XOR2_X1 U340 ( .A(n380), .B(n346), .Z(n297) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U343 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U344 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n301) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(G29GAT), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(KEYINPUT7), .B(n302), .Z(n377) );
  XOR2_X1 U348 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n304) );
  XNOR2_X1 U349 ( .A(G134GAT), .B(KEYINPUT66), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n377), .B(n305), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n548) );
  XOR2_X1 U353 ( .A(KEYINPUT89), .B(G204GAT), .Z(n309) );
  NAND2_X1 U354 ( .A1(G228GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U356 ( .A(n310), .B(KEYINPUT23), .Z(n314) );
  XNOR2_X1 U357 ( .A(G106GAT), .B(G78GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n311), .B(G148GAT), .ZN(n383) );
  XNOR2_X1 U359 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n312), .B(KEYINPUT2), .ZN(n337) );
  XNOR2_X1 U361 ( .A(n383), .B(n337), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U363 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n316) );
  XNOR2_X1 U364 ( .A(KEYINPUT22), .B(KEYINPUT88), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U366 ( .A(n318), .B(n317), .Z(n321) );
  XOR2_X1 U367 ( .A(G141GAT), .B(G22GAT), .Z(n363) );
  XNOR2_X1 U368 ( .A(n363), .B(n319), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U370 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n323) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G211GAT), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n325) );
  XOR2_X1 U373 ( .A(G218GAT), .B(KEYINPUT21), .Z(n324) );
  XOR2_X1 U374 ( .A(n325), .B(n324), .Z(n357) );
  XOR2_X1 U375 ( .A(n326), .B(n357), .Z(n455) );
  XOR2_X1 U376 ( .A(KEYINPUT4), .B(G57GAT), .Z(n328) );
  XNOR2_X1 U377 ( .A(G1GAT), .B(G120GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n345) );
  XOR2_X1 U379 ( .A(G148GAT), .B(G127GAT), .Z(n330) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(G141GAT), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n332) );
  XOR2_X1 U382 ( .A(G162GAT), .B(G85GAT), .Z(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n341) );
  XNOR2_X1 U384 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n333), .B(KEYINPUT5), .ZN(n334) );
  XOR2_X1 U386 ( .A(n334), .B(KEYINPUT90), .Z(n339) );
  XOR2_X1 U387 ( .A(KEYINPUT0), .B(KEYINPUT81), .Z(n336) );
  XNOR2_X1 U388 ( .A(G113GAT), .B(G134GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n428) );
  XNOR2_X1 U390 ( .A(n428), .B(n337), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n343) );
  NAND2_X1 U393 ( .A1(G225GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U395 ( .A(n345), .B(n344), .Z(n465) );
  INV_X1 U396 ( .A(n465), .ZN(n510) );
  XOR2_X1 U397 ( .A(G8GAT), .B(G183GAT), .Z(n396) );
  XOR2_X1 U398 ( .A(n346), .B(n396), .Z(n348) );
  NAND2_X1 U399 ( .A1(G226GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U401 ( .A(G92GAT), .B(G64GAT), .Z(n350) );
  XNOR2_X1 U402 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U404 ( .A(G176GAT), .B(n351), .ZN(n390) );
  XNOR2_X1 U405 ( .A(n352), .B(n390), .ZN(n360) );
  XNOR2_X1 U406 ( .A(KEYINPUT17), .B(KEYINPUT82), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n353), .B(KEYINPUT19), .ZN(n354) );
  XOR2_X1 U408 ( .A(n354), .B(KEYINPUT83), .Z(n356) );
  XNOR2_X1 U409 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n440) );
  INV_X1 U411 ( .A(n357), .ZN(n358) );
  XOR2_X1 U412 ( .A(n440), .B(n358), .Z(n359) );
  XOR2_X1 U413 ( .A(n360), .B(n359), .Z(n512) );
  INV_X1 U414 ( .A(n512), .ZN(n469) );
  XOR2_X1 U415 ( .A(KEYINPUT47), .B(KEYINPUT111), .Z(n414) );
  XOR2_X1 U416 ( .A(KEYINPUT70), .B(KEYINPUT67), .Z(n362) );
  XNOR2_X1 U417 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n367) );
  XOR2_X1 U419 ( .A(G50GAT), .B(G36GAT), .Z(n365) );
  XNOR2_X1 U420 ( .A(n363), .B(KEYINPUT68), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U422 ( .A(n367), .B(n366), .Z(n369) );
  NAND2_X1 U423 ( .A1(G229GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U425 ( .A(G113GAT), .B(G15GAT), .Z(n371) );
  XNOR2_X1 U426 ( .A(G169GAT), .B(G197GAT), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U428 ( .A(n373), .B(n372), .Z(n379) );
  XOR2_X1 U429 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n375) );
  XNOR2_X1 U430 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n564) );
  XNOR2_X1 U434 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n392) );
  XOR2_X1 U435 ( .A(n380), .B(KEYINPUT76), .Z(n382) );
  NAND2_X1 U436 ( .A1(G230GAT), .A2(G233GAT), .ZN(n381) );
  XOR2_X1 U437 ( .A(G57GAT), .B(KEYINPUT13), .Z(n397) );
  XNOR2_X1 U438 ( .A(n289), .B(n397), .ZN(n389) );
  XOR2_X1 U439 ( .A(G120GAT), .B(G71GAT), .Z(n426) );
  XNOR2_X1 U440 ( .A(n426), .B(n383), .ZN(n387) );
  XOR2_X1 U441 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n385) );
  XNOR2_X1 U442 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n391), .B(n390), .ZN(n569) );
  NOR2_X1 U445 ( .A1(n564), .A2(n554), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n393), .B(KEYINPUT46), .ZN(n411) );
  XOR2_X1 U447 ( .A(G155GAT), .B(G78GAT), .Z(n395) );
  XNOR2_X1 U448 ( .A(G22GAT), .B(G211GAT), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n410) );
  XOR2_X1 U450 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U451 ( .A1(G231GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U453 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n401) );
  XNOR2_X1 U454 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U456 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U457 ( .A(G15GAT), .B(G127GAT), .Z(n427) );
  XOR2_X1 U458 ( .A(KEYINPUT12), .B(G64GAT), .Z(n405) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(G71GAT), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n427), .B(n406), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U463 ( .A(n410), .B(n409), .Z(n558) );
  INV_X1 U464 ( .A(n558), .ZN(n573) );
  NOR2_X1 U465 ( .A1(n411), .A2(n573), .ZN(n412) );
  NAND2_X1 U466 ( .A1(n412), .A2(n548), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n414), .B(n413), .ZN(n421) );
  XOR2_X1 U468 ( .A(n548), .B(KEYINPUT99), .Z(n415) );
  XNOR2_X1 U469 ( .A(KEYINPUT36), .B(n415), .ZN(n578) );
  NOR2_X1 U470 ( .A1(n558), .A2(n578), .ZN(n417) );
  XNOR2_X1 U471 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n418) );
  NAND2_X1 U473 ( .A1(n564), .A2(n418), .ZN(n419) );
  NOR2_X1 U474 ( .A1(n569), .A2(n419), .ZN(n420) );
  XNOR2_X1 U475 ( .A(KEYINPUT48), .B(n422), .ZN(n522) );
  NOR2_X1 U476 ( .A1(n469), .A2(n522), .ZN(n423) );
  XOR2_X1 U477 ( .A(n423), .B(KEYINPUT54), .Z(n424) );
  NAND2_X1 U478 ( .A1(n455), .A2(n563), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n425), .B(KEYINPUT55), .ZN(n441) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U482 ( .A(KEYINPUT20), .B(G183GAT), .Z(n431) );
  NAND2_X1 U483 ( .A1(G227GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U485 ( .A(n433), .B(n432), .Z(n438) );
  XOR2_X1 U486 ( .A(G176GAT), .B(G190GAT), .Z(n435) );
  XNOR2_X1 U487 ( .A(G43GAT), .B(G99GAT), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n436), .B(KEYINPUT84), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U491 ( .A(n440), .B(n439), .Z(n472) );
  INV_X1 U492 ( .A(n472), .ZN(n526) );
  NAND2_X1 U493 ( .A1(n441), .A2(n526), .ZN(n557) );
  NOR2_X1 U494 ( .A1(n548), .A2(n557), .ZN(n444) );
  NOR2_X1 U495 ( .A1(n564), .A2(n569), .ZN(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT77), .B(n445), .Z(n481) );
  NAND2_X1 U497 ( .A1(n548), .A2(n573), .ZN(n446) );
  XOR2_X1 U498 ( .A(KEYINPUT16), .B(n446), .Z(n463) );
  XOR2_X1 U499 ( .A(n512), .B(KEYINPUT91), .Z(n447) );
  XNOR2_X1 U500 ( .A(n447), .B(KEYINPUT27), .ZN(n457) );
  NAND2_X1 U501 ( .A1(n510), .A2(n457), .ZN(n448) );
  XNOR2_X1 U502 ( .A(KEYINPUT92), .B(n448), .ZN(n523) );
  XOR2_X1 U503 ( .A(n455), .B(KEYINPUT28), .Z(n517) );
  OR2_X1 U504 ( .A1(n523), .A2(n517), .ZN(n449) );
  NOR2_X1 U505 ( .A1(n526), .A2(n449), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n450), .B(KEYINPUT93), .ZN(n462) );
  NOR2_X1 U507 ( .A1(n472), .A2(n469), .ZN(n451) );
  XOR2_X1 U508 ( .A(KEYINPUT94), .B(n451), .Z(n452) );
  NAND2_X1 U509 ( .A1(n452), .A2(n455), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n453), .B(KEYINPUT95), .ZN(n454) );
  XNOR2_X1 U511 ( .A(KEYINPUT25), .B(n454), .ZN(n459) );
  NOR2_X1 U512 ( .A1(n526), .A2(n455), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n456), .B(KEYINPUT26), .ZN(n562) );
  NAND2_X1 U514 ( .A1(n457), .A2(n562), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n465), .A2(n460), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n477) );
  NAND2_X1 U518 ( .A1(n463), .A2(n477), .ZN(n495) );
  INV_X1 U519 ( .A(n495), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n481), .A2(n464), .ZN(n475) );
  NOR2_X1 U521 ( .A1(n465), .A2(n475), .ZN(n467) );
  XNOR2_X1 U522 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U524 ( .A(G1GAT), .B(n468), .Z(G1324GAT) );
  NOR2_X1 U525 ( .A1(n469), .A2(n475), .ZN(n471) );
  XNOR2_X1 U526 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n471), .B(n470), .ZN(G1325GAT) );
  NOR2_X1 U528 ( .A1(n472), .A2(n475), .ZN(n474) );
  XNOR2_X1 U529 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  INV_X1 U531 ( .A(n517), .ZN(n525) );
  NOR2_X1 U532 ( .A1(n525), .A2(n475), .ZN(n476) );
  XOR2_X1 U533 ( .A(G22GAT), .B(n476), .Z(G1327GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT98), .B(KEYINPUT39), .Z(n486) );
  NAND2_X1 U535 ( .A1(n558), .A2(n477), .ZN(n478) );
  NOR2_X1 U536 ( .A1(n578), .A2(n478), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT37), .B(n479), .ZN(n509) );
  INV_X1 U538 ( .A(n509), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n481), .A2(n480), .ZN(n484) );
  XNOR2_X1 U540 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(KEYINPUT38), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n491) );
  NAND2_X1 U543 ( .A1(n491), .A2(n510), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(n487), .ZN(G1328GAT) );
  NAND2_X1 U546 ( .A1(n491), .A2(n512), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G36GAT), .B(n488), .ZN(G1329GAT) );
  NAND2_X1 U548 ( .A1(n526), .A2(n491), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT40), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  XNOR2_X1 U551 ( .A(G50GAT), .B(KEYINPUT102), .ZN(n493) );
  NAND2_X1 U552 ( .A1(n517), .A2(n491), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1331GAT) );
  INV_X1 U554 ( .A(n554), .ZN(n494) );
  NAND2_X1 U555 ( .A1(n564), .A2(n494), .ZN(n508) );
  NOR2_X1 U556 ( .A1(n508), .A2(n495), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT103), .B(n496), .Z(n505) );
  NAND2_X1 U558 ( .A1(n510), .A2(n505), .ZN(n500) );
  XOR2_X1 U559 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n498) );
  XNOR2_X1 U560 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U563 ( .A1(n512), .A2(n505), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(KEYINPUT106), .ZN(n502) );
  XNOR2_X1 U565 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  XOR2_X1 U566 ( .A(G71GAT), .B(KEYINPUT107), .Z(n504) );
  NAND2_X1 U567 ( .A1(n505), .A2(n526), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U570 ( .A1(n505), .A2(n517), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NOR2_X1 U572 ( .A1(n509), .A2(n508), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n518), .A2(n510), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n518), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n513), .B(KEYINPUT108), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G92GAT), .B(n514), .ZN(G1337GAT) );
  XOR2_X1 U578 ( .A(G99GAT), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U579 ( .A1(n518), .A2(n526), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1338GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n520) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U584 ( .A(G106GAT), .B(n521), .Z(G1339GAT) );
  NOR2_X1 U585 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U586 ( .A(KEYINPUT113), .B(n524), .Z(n539) );
  AND2_X1 U587 ( .A1(n525), .A2(n539), .ZN(n527) );
  NAND2_X1 U588 ( .A1(n527), .A2(n526), .ZN(n534) );
  NOR2_X1 U589 ( .A1(n564), .A2(n534), .ZN(n528) );
  XOR2_X1 U590 ( .A(n528), .B(KEYINPUT114), .Z(n529) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  NOR2_X1 U592 ( .A1(n554), .A2(n534), .ZN(n531) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U595 ( .A1(n558), .A2(n534), .ZN(n532) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(n532), .Z(n533) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  NOR2_X1 U598 ( .A1(n534), .A2(n548), .ZN(n538) );
  XOR2_X1 U599 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n536) );
  XNOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U603 ( .A1(n539), .A2(n562), .ZN(n547) );
  NOR2_X1 U604 ( .A1(n564), .A2(n547), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1344GAT) );
  NOR2_X1 U607 ( .A1(n554), .A2(n547), .ZN(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n544), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n558), .A2(n547), .ZN(n545) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(n545), .Z(n546) );
  XNOR2_X1 U613 ( .A(G155GAT), .B(n546), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(G162GAT), .B(n549), .Z(G1347GAT) );
  NOR2_X1 U616 ( .A1(n564), .A2(n557), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n553) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n554), .A2(n557), .ZN(n555) );
  XOR2_X1 U623 ( .A(n556), .B(n555), .Z(G1349GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(G183GAT), .B(n559), .Z(G1350GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n577) );
  NOR2_X1 U630 ( .A1(n564), .A2(n577), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT121), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(n568), .B(n567), .Z(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n571) );
  INV_X1 U635 ( .A(n577), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n574), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n572), .ZN(G1353GAT) );
  XOR2_X1 U639 ( .A(G211GAT), .B(KEYINPUT125), .Z(n576) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G218GAT), .B(n581), .Z(G1355GAT) );
endmodule

