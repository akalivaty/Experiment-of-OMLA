//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  NOR2_X1   g004(.A1(G237), .A2(G953), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n191), .A2(G143), .A3(G214), .ZN(new_n192));
  AOI21_X1  g006(.A(G143), .B1(new_n191), .B2(G214), .ZN(new_n193));
  OAI21_X1  g007(.A(G131), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G237), .ZN(new_n195));
  INV_X1    g009(.A(G953), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G214), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(G143), .A3(G214), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n194), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(G146), .B(new_n206), .C1(new_n210), .C2(new_n204), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n210), .A2(KEYINPUT19), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(KEYINPUT19), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n203), .B(new_n211), .C1(G146), .C2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n200), .B1(new_n199), .B2(new_n201), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT18), .ZN(new_n217));
  NAND2_X1  g031(.A1(KEYINPUT18), .A2(G131), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n199), .A2(new_n201), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G125), .B(G140), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n190), .B1(new_n215), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n194), .A2(new_n225), .A3(new_n202), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n216), .A2(KEYINPUT17), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n206), .B1(new_n210), .B2(new_n204), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n221), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n226), .A2(new_n227), .A3(new_n229), .A4(new_n211), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n190), .A3(new_n223), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n230), .A2(KEYINPUT81), .A3(new_n223), .A4(new_n190), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n224), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(G475), .A2(G902), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n187), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n190), .B1(new_n230), .B2(new_n223), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n233), .B2(new_n234), .ZN(new_n240));
  OAI21_X1  g054(.A(G475), .B1(new_n240), .B2(G902), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  AOI211_X1 g058(.A(KEYINPUT82), .B(new_n224), .C1(new_n233), .C2(new_n234), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT20), .B(new_n236), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT83), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT83), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G116), .B(G122), .ZN(new_n251));
  INV_X1    g065(.A(G107), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n198), .A2(G128), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n198), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT64), .A2(G134), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT13), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n254), .B1(new_n256), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n198), .A2(KEYINPUT13), .A3(G128), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(KEYINPUT84), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(G134), .B1(new_n265), .B2(KEYINPUT84), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n253), .B(new_n263), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT14), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n251), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G122), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G116), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n252), .B1(new_n274), .B2(KEYINPUT14), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n272), .A2(new_n275), .B1(new_n252), .B2(new_n251), .ZN(new_n276));
  INV_X1    g090(.A(new_n263), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n257), .A2(new_n262), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n270), .A2(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT71), .B(G217), .Z(new_n281));
  XOR2_X1   g095(.A(KEYINPUT9), .B(G234), .Z(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n196), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT85), .ZN(new_n285));
  INV_X1    g099(.A(new_n283), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n270), .A2(new_n279), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n280), .A2(KEYINPUT85), .A3(new_n283), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G478), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(KEYINPUT15), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n291), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n196), .A2(G952), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(G234), .B2(G237), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI211_X1 g111(.A(new_n289), .B(new_n196), .C1(G234), .C2(G237), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT21), .B(G898), .Z(new_n300));
  OAI21_X1  g114(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n248), .A2(new_n250), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G137), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n260), .A2(new_n261), .B1(KEYINPUT11), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(KEYINPUT11), .A3(G134), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT11), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G137), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G131), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(KEYINPUT64), .A2(G134), .ZN(new_n312));
  NOR2_X1   g126(.A1(KEYINPUT64), .A2(G134), .ZN(new_n313));
  OAI22_X1  g127(.A1(new_n312), .A2(new_n313), .B1(new_n308), .B2(G137), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n314), .A2(new_n200), .A3(new_n307), .A4(new_n309), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(KEYINPUT65), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n317), .B(G131), .C1(new_n306), .C2(new_n310), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(G104), .A3(new_n252), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n189), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n323));
  OAI22_X1  g137(.A1(new_n189), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n324));
  INV_X1    g138(.A(G101), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n252), .A2(G104), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n189), .A2(G107), .ZN(new_n328));
  OAI21_X1  g142(.A(G101), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G128), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n221), .A3(G143), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n198), .B(G146), .C1(new_n331), .C2(KEYINPUT1), .ZN(new_n333));
  XNOR2_X1  g147(.A(G143), .B(G146), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G128), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n330), .A2(new_n332), .A3(new_n333), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n332), .A3(new_n333), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n326), .A3(new_n329), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n320), .A2(new_n340), .A3(KEYINPUT12), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n320), .A2(new_n340), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT12), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n320), .A2(new_n340), .A3(KEYINPUT78), .A4(KEYINPUT12), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n339), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G101), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT4), .A3(new_n326), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT0), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n334), .B1(new_n354), .B2(new_n331), .ZN(new_n355));
  XOR2_X1   g169(.A(KEYINPUT0), .B(G128), .Z(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n334), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n351), .A2(new_n358), .A3(G101), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n330), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT10), .A3(new_n338), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n350), .A2(new_n360), .A3(new_n319), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n348), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G140), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n196), .A2(G227), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n360), .A2(new_n350), .A3(new_n362), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n320), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n363), .A2(new_n367), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n364), .A2(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G469), .ZN(new_n373));
  NAND2_X1  g187(.A1(G469), .A2(G902), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n348), .A2(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n363), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n368), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G469), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n289), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n373), .A2(new_n374), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n282), .A2(new_n289), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n382), .A2(G221), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(KEYINPUT76), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(G116), .B(G119), .Z(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT2), .B(G113), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n353), .A2(new_n388), .A3(new_n359), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n386), .A2(new_n387), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n391));
  INV_X1    g205(.A(G119), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G116), .ZN(new_n393));
  OAI211_X1 g207(.A(G113), .B(new_n393), .C1(new_n386), .C2(new_n391), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n361), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  XOR2_X1   g210(.A(G110), .B(G122), .Z(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n397), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n389), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(KEYINPUT6), .A3(new_n400), .ZN(new_n401));
  MUX2_X1   g215(.A(new_n338), .B(new_n357), .S(G125), .Z(new_n402));
  NAND2_X1  g216(.A1(new_n196), .A2(G224), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n396), .A2(new_n405), .A3(new_n397), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n402), .B1(KEYINPUT79), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(KEYINPUT79), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n394), .A2(new_n390), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n330), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n395), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n397), .B(KEYINPUT8), .Z(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n402), .A2(KEYINPUT79), .A3(new_n408), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n411), .A2(new_n400), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n407), .A2(new_n289), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(KEYINPUT80), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G214), .B1(G237), .B2(G902), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n304), .A2(new_n385), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(G472), .A2(G902), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n191), .A2(G210), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(new_n325), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n428), .B(new_n429), .Z(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT28), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n316), .A2(new_n318), .A3(new_n357), .ZN(new_n433));
  INV_X1    g247(.A(new_n388), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n260), .A2(new_n305), .A3(new_n261), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n259), .A2(G137), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n435), .A2(KEYINPUT66), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G131), .B1(new_n435), .B2(KEYINPUT66), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n338), .B(new_n315), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT68), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n433), .A2(new_n442), .A3(new_n434), .A4(new_n439), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n433), .A2(new_n439), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n388), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n432), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n440), .A2(new_n432), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT69), .B(new_n431), .C1(new_n447), .C2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT67), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n451), .A3(KEYINPUT30), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(KEYINPUT30), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n433), .A2(new_n439), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n457), .A2(new_n388), .B1(new_n441), .B2(new_n443), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT31), .B1(new_n458), .B2(new_n430), .ZN(new_n459));
  AOI211_X1 g273(.A(KEYINPUT67), .B(new_n453), .C1(new_n433), .C2(new_n439), .ZN(new_n460));
  AND4_X1   g274(.A1(new_n433), .A2(new_n439), .A3(new_n454), .A4(new_n455), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n388), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n462), .A2(KEYINPUT31), .A3(new_n444), .A4(new_n430), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n450), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n441), .A2(new_n443), .B1(new_n388), .B2(new_n445), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n448), .B1(new_n466), .B2(new_n432), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT69), .B1(new_n467), .B2(new_n431), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n426), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT32), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT70), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n447), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT70), .B1(new_n466), .B2(new_n432), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n448), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT29), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(new_n431), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n448), .B(new_n430), .C1(new_n466), .C2(new_n432), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n476), .C1(new_n430), .C2(new_n458), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n289), .ZN(new_n480));
  OAI21_X1  g294(.A(G472), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n431), .B1(new_n447), .B2(new_n449), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n462), .A2(new_n444), .A3(new_n430), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT31), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n463), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n488), .A3(new_n450), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT32), .A3(new_n426), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n471), .A2(new_n481), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n196), .A2(G221), .A3(G234), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT73), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT22), .B(G137), .Z(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT74), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n392), .A2(G128), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n331), .A2(G119), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT24), .B(G110), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n497), .B1(KEYINPUT72), .B2(KEYINPUT23), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n503), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n502), .B1(new_n505), .B2(new_n497), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n501), .B1(new_n506), .B2(G110), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(new_n211), .C1(G146), .C2(new_n210), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n229), .A2(new_n211), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(G110), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n509), .B(new_n510), .C1(new_n499), .C2(new_n500), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n496), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n495), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n289), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT25), .ZN(new_n516));
  INV_X1    g330(.A(new_n281), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(G234), .B2(new_n289), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n513), .A2(new_n519), .A3(new_n289), .A4(new_n514), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n513), .A2(new_n514), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n518), .A2(G902), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(KEYINPUT75), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n513), .A2(new_n514), .A3(new_n524), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n425), .A2(new_n491), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(G101), .ZN(G3));
  INV_X1    g346(.A(new_n469), .ZN(new_n533));
  INV_X1    g347(.A(G472), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n489), .B2(new_n289), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n533), .A2(new_n535), .A3(new_n385), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n248), .A2(new_n250), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n419), .A2(new_n420), .ZN(new_n538));
  INV_X1    g352(.A(new_n420), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n407), .A2(new_n418), .A3(new_n289), .A4(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n538), .A2(new_n423), .A3(new_n301), .A4(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n288), .A2(new_n543), .A3(new_n290), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n284), .A2(KEYINPUT33), .A3(new_n287), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n289), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G478), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n291), .A2(G478), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT86), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT86), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n551), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n537), .A2(new_n542), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n536), .A2(new_n530), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT34), .B(G104), .Z(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(G6));
  OR2_X1    g371(.A1(new_n244), .A2(new_n245), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n187), .B1(new_n559), .B2(new_n237), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n241), .B(KEYINPUT87), .Z(new_n561));
  NAND4_X1  g375(.A1(new_n560), .A2(new_n246), .A3(new_n561), .A4(new_n294), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n541), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n536), .A2(new_n530), .A3(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G107), .Z(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(G9));
  OAI21_X1  g382(.A(new_n289), .B1(new_n465), .B2(new_n468), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G472), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n496), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(new_n512), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n524), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n521), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n570), .A2(new_n469), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n570), .A2(KEYINPUT90), .A3(new_n469), .A4(new_n575), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n425), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT37), .B(G110), .Z(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(G12));
  INV_X1    g396(.A(new_n385), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n538), .A2(new_n423), .A3(new_n540), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AND4_X1   g399(.A1(new_n491), .A2(new_n583), .A3(new_n585), .A4(new_n575), .ZN(new_n586));
  INV_X1    g400(.A(G900), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n296), .B1(new_n298), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n562), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G128), .ZN(G30));
  XNOR2_X1  g405(.A(new_n422), .B(KEYINPUT38), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n592), .A2(new_n423), .ZN(new_n593));
  INV_X1    g407(.A(new_n575), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n242), .A2(new_n246), .A3(new_n249), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n249), .B1(new_n242), .B2(new_n246), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n294), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n485), .B(G472), .C1(new_n466), .C2(new_n430), .ZN(new_n599));
  NAND2_X1  g413(.A1(G472), .A2(G902), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT91), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n471), .A2(new_n603), .A3(new_n490), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n593), .A2(new_n594), .A3(new_n598), .A4(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT92), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n588), .B(KEYINPUT39), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n385), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(KEYINPUT40), .Z(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G143), .ZN(G45));
  NAND2_X1  g425(.A1(new_n537), .A2(new_n553), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n588), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n586), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G146), .ZN(G48));
  AOI22_X1  g429(.A1(new_n348), .A2(new_n371), .B1(new_n376), .B2(new_n368), .ZN(new_n616));
  OAI21_X1  g430(.A(G469), .B1(new_n616), .B2(G902), .ZN(new_n617));
  INV_X1    g431(.A(new_n383), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n380), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n554), .A2(new_n491), .A3(new_n530), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT93), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT41), .B(G113), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G15));
  INV_X1    g437(.A(new_n530), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n489), .A2(KEYINPUT32), .A3(new_n426), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT32), .B1(new_n489), .B2(new_n426), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n624), .B1(new_n627), .B2(new_n481), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n628), .A2(KEYINPUT94), .A3(new_n563), .A4(new_n619), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n563), .A2(new_n491), .A3(new_n530), .A4(new_n619), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT94), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G116), .ZN(G18));
  INV_X1    g448(.A(new_n304), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT95), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n619), .A2(new_n585), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n380), .A2(new_n617), .A3(new_n618), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT95), .B1(new_n638), .B2(new_n584), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n491), .A2(new_n635), .A3(new_n640), .A4(new_n575), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G119), .ZN(G21));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n644));
  AOI211_X1 g458(.A(new_n644), .B(new_n534), .C1(new_n489), .C2(new_n289), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT96), .B1(new_n569), .B2(G472), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT97), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n522), .B2(new_n529), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n521), .A2(KEYINPUT97), .A3(new_n528), .A4(new_n525), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n475), .A2(new_n431), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n488), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(new_n426), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n647), .A2(new_n619), .A3(new_n651), .A4(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n597), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n537), .A2(KEYINPUT98), .A3(new_n294), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n659), .A3(new_n542), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n643), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n570), .A2(new_n644), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n535), .A2(KEYINPUT96), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n651), .A2(new_n662), .A3(new_n655), .A4(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n660), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n664), .A2(KEYINPUT99), .A3(new_n619), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G122), .ZN(G24));
  NOR3_X1   g482(.A1(new_n645), .A2(new_n646), .A3(new_n654), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n575), .A3(new_n613), .A4(new_n640), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G125), .ZN(G27));
  INV_X1    g485(.A(new_n423), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n422), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n612), .A2(new_n588), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n373), .A2(new_n380), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n374), .B(KEYINPUT100), .Z(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n383), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(KEYINPUT101), .A3(new_n628), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n675), .A2(new_n679), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n491), .A2(new_n530), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n681), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n491), .A2(new_n651), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n680), .A2(new_n688), .A3(KEYINPUT42), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G131), .ZN(G33));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n685), .B1(new_n692), .B2(new_n589), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT102), .B1(new_n562), .B2(new_n588), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n694), .A2(new_n679), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n673), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G134), .ZN(G36));
  OR2_X1    g511(.A1(new_n372), .A2(KEYINPUT45), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n372), .A2(KEYINPUT45), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(G469), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(KEYINPUT46), .A3(new_n678), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n380), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT46), .B1(new_n700), .B2(new_n678), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n618), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n704), .A2(new_n607), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n595), .A2(new_n596), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n553), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n707), .A2(KEYINPUT43), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(KEYINPUT43), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n594), .B1(new_n570), .B2(new_n469), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n712), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(KEYINPUT103), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(KEYINPUT103), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n714), .B(new_n673), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G137), .ZN(G39));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n704), .B(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n491), .A2(new_n530), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n675), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G140), .ZN(G42));
  NAND3_X1  g538(.A1(new_n708), .A2(new_n296), .A3(new_n709), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n656), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n592), .A2(new_n423), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n726), .A2(KEYINPUT50), .A3(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n708), .A2(new_n296), .A3(new_n709), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n733), .A2(new_n664), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n380), .A2(new_n617), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n384), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n673), .B(new_n734), .C1(new_n721), .C2(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n739));
  INV_X1    g553(.A(new_n604), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n673), .A2(new_n619), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n624), .A3(new_n297), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n743), .A2(new_n537), .A3(new_n553), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n741), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n733), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n669), .A2(new_n575), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n739), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n745), .B(KEYINPUT109), .C1(new_n747), .C2(new_n748), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n738), .A2(KEYINPUT110), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n732), .A2(new_n737), .A3(new_n752), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n747), .A2(new_n748), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n744), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n757), .B2(KEYINPUT109), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n295), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n732), .A2(new_n757), .A3(new_n737), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n761), .B1(new_n763), .B2(KEYINPUT51), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(KEYINPUT108), .A3(new_n739), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n743), .A2(new_n612), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n760), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n733), .A2(new_n688), .A3(new_n746), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT48), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n734), .A2(new_n640), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n768), .A2(KEYINPUT111), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n696), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n687), .B2(new_n689), .ZN(new_n775));
  INV_X1    g589(.A(new_n294), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n612), .B1(new_n537), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n424), .A2(new_n302), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n536), .A3(new_n530), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n580), .A2(new_n779), .A3(new_n531), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n647), .A2(new_n613), .A3(new_n655), .A4(new_n679), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n560), .A2(new_n246), .A3(new_n561), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n782), .A2(new_n385), .A3(new_n588), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n491), .A3(new_n776), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n594), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n780), .B1(new_n785), .B2(new_n673), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n620), .A2(new_n641), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n629), .B2(new_n632), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n667), .A2(KEYINPUT104), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT104), .B1(new_n667), .B2(new_n788), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n775), .B(new_n786), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n586), .B1(new_n589), .B2(new_n613), .ZN(new_n794));
  INV_X1    g608(.A(new_n588), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n604), .A2(new_n594), .A3(new_n795), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n585), .A2(new_n658), .A3(new_n659), .A4(new_n679), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n670), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT106), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT106), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n794), .A2(KEYINPUT52), .A3(new_n670), .A4(new_n798), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(KEYINPUT105), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(KEYINPUT105), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n802), .B(new_n804), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n792), .A2(new_n793), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n801), .A2(new_n805), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT53), .B1(new_n791), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n809), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT107), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n786), .B2(new_n696), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n781), .A2(new_n784), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n575), .A3(new_n673), .ZN(new_n816));
  INV_X1    g630(.A(new_n780), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n813), .A2(new_n816), .A3(new_n817), .A4(new_n696), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n667), .A2(new_n788), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n793), .B1(new_n687), .B2(new_n689), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n808), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n793), .B1(new_n791), .B2(new_n810), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n812), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n760), .A2(new_n766), .A3(new_n772), .A4(new_n767), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n829), .B2(new_n770), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n773), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n832));
  OR2_X1    g646(.A1(G952), .A2(G953), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n773), .A2(new_n830), .A3(new_n834), .A4(new_n827), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n384), .B1(new_n735), .B2(KEYINPUT49), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n649), .A2(new_n650), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n837), .B(new_n838), .C1(KEYINPUT49), .C2(new_n735), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n604), .A2(new_n592), .A3(new_n707), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n840), .A3(new_n423), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n836), .A2(new_n841), .ZN(G75));
  NOR2_X1   g656(.A1(new_n196), .A2(G952), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n289), .B1(new_n822), .B2(new_n823), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(G210), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n401), .A2(new_n406), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(new_n404), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT55), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n846), .B2(new_n845), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n845), .A2(new_n847), .A3(new_n853), .ZN(new_n855));
  INV_X1    g669(.A(new_n850), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n843), .B1(new_n854), .B2(new_n857), .ZN(G51));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n677), .B(KEYINPUT57), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n822), .A2(new_n823), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT54), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n863), .B2(new_n825), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n859), .B1(new_n864), .B2(new_n616), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n844), .A2(G469), .A3(new_n698), .A4(new_n699), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n824), .B1(new_n822), .B2(new_n823), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n860), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(KEYINPUT115), .A3(new_n378), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n865), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n843), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n871), .A2(KEYINPUT116), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(G54));
  NAND3_X1  g691(.A1(new_n844), .A2(KEYINPUT58), .A3(G475), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n559), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n843), .ZN(G60));
  AND2_X1   g694(.A1(new_n544), .A2(new_n545), .ZN(new_n881));
  NAND2_X1  g695(.A1(G478), .A2(G902), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT59), .Z(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n881), .B(new_n884), .C1(new_n867), .C2(new_n868), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n881), .B1(new_n826), .B2(new_n884), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(KEYINPUT117), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(KEYINPUT117), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n843), .B(new_n886), .C1(new_n888), .C2(new_n889), .ZN(G63));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n891));
  NAND2_X1  g705(.A1(G217), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT118), .Z(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT60), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n822), .B2(new_n823), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n523), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(KEYINPUT119), .A3(new_n872), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n573), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT119), .B1(new_n897), .B2(new_n872), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n891), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n891), .B1(new_n896), .B2(KEYINPUT120), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n872), .A4(new_n899), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(G66));
  AOI21_X1  g720(.A(new_n196), .B1(new_n300), .B2(G224), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n817), .B1(new_n789), .B2(new_n790), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(new_n196), .ZN(new_n909));
  INV_X1    g723(.A(G898), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n848), .B1(new_n910), .B2(G953), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n909), .B(new_n911), .ZN(G69));
  NOR2_X1   g726(.A1(new_n196), .A2(G900), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT123), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n775), .B(KEYINPUT124), .Z(new_n915));
  AND2_X1   g729(.A1(new_n794), .A2(new_n670), .ZN(new_n916));
  INV_X1    g730(.A(new_n705), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n658), .A2(new_n659), .A3(new_n585), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n688), .A3(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n718), .A2(new_n723), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n915), .A2(new_n916), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n914), .B1(new_n921), .B2(new_n196), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n457), .B(new_n214), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n610), .A2(new_n916), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT62), .Z(new_n926));
  NOR2_X1   g740(.A1(new_n608), .A2(new_n674), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n628), .A2(new_n777), .A3(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n718), .A2(new_n723), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT121), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n926), .A2(new_n932), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n196), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n924), .B1(new_n935), .B2(new_n923), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n196), .B1(G227), .B2(G900), .ZN(new_n937));
  INV_X1    g751(.A(new_n924), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n936), .B(new_n940), .ZN(G72));
  NOR2_X1   g755(.A1(new_n458), .A2(new_n431), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n908), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n931), .A2(new_n944), .A3(new_n933), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n600), .B(KEYINPUT63), .Z(new_n946));
  AOI21_X1  g760(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n921), .B2(new_n908), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n458), .A2(new_n431), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n943), .A2(new_n946), .A3(new_n949), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT125), .Z(new_n953));
  NAND3_X1  g767(.A1(new_n809), .A2(new_n811), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n872), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n956));
  OR3_X1    g770(.A1(new_n947), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n947), .B2(new_n955), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(G57));
endmodule


