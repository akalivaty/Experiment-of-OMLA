//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n447, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT66), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT68), .Z(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  XOR2_X1   g033(.A(G325), .B(KEYINPUT69), .Z(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT70), .Z(new_n461));
  NAND2_X1  g036(.A1(new_n457), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(new_n465), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(G160));
  INV_X1    g054(.A(new_n473), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(KEYINPUT71), .A3(G136), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n482), .B1(new_n473), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n472), .B1(new_n469), .B2(new_n470), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n481), .A2(new_n484), .B1(G124), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G100), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n487), .A2(new_n472), .A3(KEYINPUT72), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT72), .B1(new_n487), .B2(new_n472), .ZN(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G112), .B2(new_n472), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  INV_X1    g067(.A(new_n470), .ZN(new_n493));
  NOR2_X1   g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n472), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  XOR2_X1   g070(.A(KEYINPUT73), .B(KEYINPUT4), .Z(new_n496));
  OR2_X1    g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n495), .A2(new_n499), .B1(G102), .B2(new_n466), .ZN(new_n500));
  INV_X1    g075(.A(G126), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n469), .B2(new_n470), .ZN(new_n502));
  AND2_X1   g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  OAI21_X1  g078(.A(G2105), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n497), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  NAND2_X1  g081(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G166));
  XNOR2_X1  g096(.A(KEYINPUT75), .B(G51), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(G89), .A3(new_n515), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n524), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n523), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n531), .A2(KEYINPUT77), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n523), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n524), .A2(new_n529), .A3(new_n526), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n529), .B1(new_n524), .B2(new_n526), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n532), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n533), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT78), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n511), .A2(new_n515), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT6), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n545), .A2(new_n547), .A3(G543), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n544), .A2(G90), .B1(G52), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n543), .A2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n509), .B2(new_n510), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT79), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n510), .ZN(new_n557));
  AOI21_X1  g132(.A(G543), .B1(KEYINPUT74), .B2(KEYINPUT5), .ZN(new_n558));
  OAI21_X1  g133(.A(G56), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(new_n560), .A3(new_n554), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n556), .A2(new_n561), .A3(G651), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n544), .A2(G81), .B1(G43), .B2(new_n548), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n511), .A2(G65), .ZN(new_n572));
  INV_X1    g147(.A(G78), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(new_n508), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(new_n544), .B2(G91), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n548), .A2(KEYINPUT80), .A3(new_n576), .A4(G53), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n545), .A2(new_n547), .A3(KEYINPUT80), .A4(G543), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT9), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n577), .A2(KEYINPUT81), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT81), .B1(new_n577), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n575), .B1(new_n581), .B2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND2_X1  g160(.A1(new_n544), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n548), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n513), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  INV_X1    g167(.A(G48), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n516), .A2(new_n592), .B1(new_n518), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n513), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n516), .A2(new_n599), .B1(new_n518), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT10), .B1(new_n516), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n511), .A2(new_n606), .A3(new_n515), .A4(G92), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n609));
  OAI21_X1  g184(.A(G66), .B1(new_n557), .B2(new_n558), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n513), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g187(.A1(new_n515), .A2(G54), .A3(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n548), .A2(G54), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n615), .B(KEYINPUT82), .C1(new_n616), .C2(new_n513), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n608), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G171), .B2(new_n620), .ZN(G284));
  OAI21_X1  g197(.A(new_n621), .B1(G171), .B2(new_n620), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(G299), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(G868), .B2(new_n625), .ZN(new_n626));
  MUX2_X1   g201(.A(new_n624), .B(new_n626), .S(KEYINPUT83), .Z(G297));
  MUX2_X1   g202(.A(new_n624), .B(new_n626), .S(KEYINPUT83), .Z(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n618), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n618), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n471), .A2(new_n466), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n480), .A2(G135), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n640), .A2(KEYINPUT85), .B1(G123), .B2(new_n485), .ZN(new_n641));
  NOR2_X1   g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(new_n472), .B2(G111), .ZN(new_n643));
  OAI221_X1 g218(.A(new_n641), .B1(KEYINPUT85), .B2(new_n640), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(KEYINPUT86), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(KEYINPUT86), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G2096), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(G2096), .B1(new_n645), .B2(new_n646), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n639), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT87), .Z(G156));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2435), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2438), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT88), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2443), .B(G2446), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1341), .B(G1348), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n665), .A2(G14), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XOR2_X1   g244(.A(G2067), .B(G2678), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n668), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT89), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n667), .A3(new_n668), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  INV_X1    g251(.A(new_n669), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n667), .A3(new_n670), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n648), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2100), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n683), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n687), .A2(KEYINPUT20), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(new_n683), .A3(new_n686), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n690), .B(new_n692), .C1(KEYINPUT20), .C2(new_n687), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(G229));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G35), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G162), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT29), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(G2090), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(G2090), .ZN(new_n706));
  INV_X1    g281(.A(G1341), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n565), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n708), .B2(G19), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n706), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n705), .B(new_n711), .C1(new_n707), .C2(new_n710), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n647), .A2(new_n701), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT100), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n708), .A2(G5), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G171), .B2(new_n708), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT101), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1961), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n712), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT31), .B(G11), .Z(new_n720));
  INV_X1    g295(.A(KEYINPUT30), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n701), .B1(new_n721), .B2(G28), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n721), .B2(G28), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n480), .A2(G141), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n485), .A2(G129), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n466), .A2(G105), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT26), .Z(new_n728));
  NAND4_X1  g303(.A1(new_n724), .A2(new_n725), .A3(new_n726), .A4(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G29), .B2(G32), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n720), .B(new_n723), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G2084), .ZN(new_n735));
  AND2_X1   g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  NOR2_X1   g311(.A1(KEYINPUT24), .A2(G34), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n736), .A2(new_n737), .A3(G29), .ZN(new_n738));
  INV_X1    g313(.A(G160), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G29), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n734), .B1(new_n735), .B2(new_n740), .C1(new_n732), .C2(new_n733), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n701), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n701), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT102), .B(G2078), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n740), .A2(new_n735), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n701), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT28), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n480), .A2(G140), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT96), .ZN(new_n751));
  OR2_X1    g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n485), .A2(G128), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n755), .A2(KEYINPUT97), .A3(G29), .ZN(new_n756));
  AOI21_X1  g331(.A(KEYINPUT97), .B1(new_n755), .B2(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n749), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n708), .A2(G4), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n618), .B2(new_n708), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G1348), .Z(new_n763));
  NAND4_X1  g338(.A1(new_n746), .A2(new_n747), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n708), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n708), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT99), .B(G1966), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n708), .A2(G20), .ZN(new_n769));
  OAI211_X1 g344(.A(KEYINPUT23), .B(new_n769), .C1(new_n625), .C2(new_n708), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(KEYINPUT23), .B2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(G1956), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n719), .A2(new_n764), .A3(new_n768), .A4(new_n773), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT98), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n776), .A2(G2105), .B1(G139), .B2(new_n480), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n466), .A2(G103), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G33), .B(new_n780), .S(G29), .Z(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G2072), .Z(new_n782));
  NOR2_X1   g357(.A1(G16), .A2(G24), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n602), .B(KEYINPUT93), .Z(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1986), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n708), .A2(G23), .ZN(new_n787));
  INV_X1    g362(.A(G288), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n708), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT33), .Z(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G1976), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n708), .A2(G6), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n595), .B2(new_n708), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  INV_X1    g369(.A(G1981), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n708), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n708), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT94), .B(G1971), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n790), .A2(G1976), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n791), .A2(new_n796), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n786), .B1(new_n802), .B2(KEYINPUT34), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n480), .A2(G131), .B1(G119), .B2(new_n485), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n472), .A2(G107), .ZN(new_n805));
  OR3_X1    g380(.A1(KEYINPUT91), .A2(G95), .A3(G2105), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT91), .B1(G95), .B2(G2105), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n806), .A2(G2104), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n804), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G25), .B(new_n809), .S(G29), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT92), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT35), .B(G1991), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n803), .B(new_n813), .C1(KEYINPUT34), .C2(new_n802), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(KEYINPUT95), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n774), .A2(new_n782), .A3(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n548), .A2(G55), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n511), .A2(G93), .A3(new_n515), .ZN(new_n821));
  AND2_X1   g396(.A1(G80), .A2(G543), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n511), .B2(G67), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n820), .B(new_n821), .C1(new_n823), .C2(new_n513), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n618), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT39), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT104), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n824), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n564), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n562), .A2(new_n824), .A3(new_n563), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n831), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n826), .B1(new_n836), .B2(G860), .ZN(G145));
  XNOR2_X1  g412(.A(new_n647), .B(G160), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n809), .B(G164), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n485), .A2(G130), .ZN(new_n843));
  NOR2_X1   g418(.A1(G106), .A2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n845));
  INV_X1    g420(.A(G142), .ZN(new_n846));
  OAI221_X1 g421(.A(new_n843), .B1(new_n844), .B2(new_n845), .C1(new_n846), .C2(new_n473), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(new_n636), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n491), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n840), .A2(new_n849), .A3(new_n841), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n755), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n777), .A2(KEYINPUT106), .A3(new_n779), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  OR3_X1    g432(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT105), .ZN(new_n858));
  OAI21_X1  g433(.A(KEYINPUT105), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(new_n730), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n730), .B1(new_n858), .B2(new_n859), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n853), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n860), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n851), .A2(new_n864), .A3(new_n852), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g443(.A(G166), .B(G288), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n595), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n869), .A2(new_n595), .ZN(new_n872));
  OAI21_X1  g447(.A(G290), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n874), .A2(new_n602), .A3(new_n870), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(KEYINPUT108), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(KEYINPUT108), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n879), .B2(new_n876), .ZN(new_n881));
  AND2_X1   g456(.A1(G299), .A2(new_n618), .ZN(new_n882));
  NOR2_X1   g457(.A1(G299), .A2(new_n618), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT107), .B1(new_n882), .B2(new_n883), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(G299), .B2(new_n618), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n885), .B1(new_n889), .B2(new_n884), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n835), .B(new_n631), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n882), .A2(new_n883), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n894), .B2(new_n891), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n881), .B(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(new_n620), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n832), .A2(G868), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n897), .A2(new_n898), .ZN(G295));
  NAND2_X1  g474(.A1(G295), .A2(KEYINPUT109), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n897), .A2(KEYINPUT109), .A3(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(G331));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n562), .A2(new_n824), .A3(new_n563), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n824), .B1(new_n563), .B2(new_n562), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT77), .B1(new_n531), .B2(new_n532), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n537), .A2(new_n538), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n835), .A2(new_n533), .A3(new_n539), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n909), .A2(G171), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G171), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n894), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n873), .A2(new_n875), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n909), .A2(new_n910), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(G301), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n910), .A3(G171), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n913), .B(new_n914), .C1(new_n890), .C2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n919), .A2(new_n866), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n889), .A2(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n893), .A2(new_n884), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(new_n917), .A3(new_n916), .A4(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(KEYINPUT111), .B(new_n894), .C1(new_n911), .C2(new_n912), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n876), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n920), .A2(new_n928), .A3(KEYINPUT112), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT112), .B1(new_n920), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n913), .B1(new_n890), .B2(new_n918), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n876), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(KEYINPUT110), .A3(new_n866), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT41), .B1(new_n886), .B2(new_n888), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n917), .B(new_n916), .C1(new_n936), .C2(new_n885), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n914), .B1(new_n937), .B2(new_n913), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n938), .B2(G37), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n939), .A3(new_n919), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n903), .B1(new_n931), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n920), .A2(new_n928), .A3(new_n941), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT44), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT113), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n927), .A2(new_n876), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n919), .A2(new_n866), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n920), .A2(new_n928), .A3(KEYINPUT112), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n941), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n940), .A2(new_n941), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT44), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n944), .A2(new_n945), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n903), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n947), .A2(new_n959), .ZN(G397));
  AND2_X1   g535(.A1(G160), .A2(G40), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT114), .B(G1384), .Z(new_n962));
  AOI21_X1  g537(.A(KEYINPUT45), .B1(new_n505), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT115), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n755), .B(new_n759), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n729), .B(G1996), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n809), .A2(new_n812), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n809), .A2(new_n812), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(G290), .A2(G1986), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n965), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(G160), .A2(G40), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n505), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n505), .A2(KEYINPUT50), .A3(new_n978), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n977), .A2(new_n979), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n983), .A2(G1348), .B1(G2067), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT118), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI221_X1 g562(.A(KEYINPUT118), .B1(new_n984), .B2(G2067), .C1(new_n983), .C2(G1348), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT60), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT121), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n618), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n990), .B2(new_n618), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n987), .A2(new_n988), .ZN(new_n995));
  OAI22_X1  g570(.A1(new_n993), .A2(new_n994), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n990), .A2(new_n618), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT121), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n995), .A2(new_n989), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n992), .ZN(new_n1000));
  INV_X1    g575(.A(new_n982), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT50), .B1(new_n505), .B2(new_n978), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n961), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n772), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n577), .A2(new_n580), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n575), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n505), .B2(new_n978), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(new_n977), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT56), .B(G2072), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1004), .A2(new_n1008), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1004), .A2(new_n1013), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n625), .A2(new_n1005), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(new_n1007), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT61), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1020), .A2(KEYINPUT61), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1021), .A2(new_n1022), .B1(new_n1023), .B2(new_n1014), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT58), .B(G1341), .Z(new_n1025));
  NAND2_X1  g600(.A1(new_n984), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n1027), .B2(G1996), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n565), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT120), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1031), .A3(new_n565), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1030), .A2(KEYINPUT59), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT59), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n996), .A2(new_n1000), .A3(new_n1024), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n995), .A2(new_n618), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1037), .A2(KEYINPUT119), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1020), .B1(new_n1037), .B2(KEYINPUT119), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1017), .B(new_n1016), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n984), .A2(G8), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1042), .B(new_n1044), .C1(new_n1043), .C2(G288), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G305), .A2(G1981), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n595), .A2(new_n795), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT49), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(KEYINPUT49), .A3(new_n1047), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1042), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n984), .B(G8), .C1(new_n1043), .C2(G288), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT52), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1045), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1056));
  OAI22_X1  g631(.A1(new_n1056), .A2(G1971), .B1(G2090), .B2(new_n1003), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1059), .B(KEYINPUT55), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1060), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(G8), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1055), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1027), .B2(G2078), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1067), .A2(new_n1009), .A3(new_n977), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1065), .A2(G2078), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1961), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1003), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1066), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1072), .B(KEYINPUT124), .ZN(new_n1075));
  INV_X1    g650(.A(new_n963), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1076), .A2(new_n961), .A3(new_n1069), .A4(new_n1011), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1066), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1074), .B1(new_n1078), .B2(G171), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1064), .B1(new_n1079), .B2(KEYINPUT54), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n735), .B(new_n961), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(G168), .C1(new_n1068), .C2(new_n767), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(G8), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1081), .B1(new_n1068), .B2(new_n767), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(G8), .A3(G286), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1087), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1082), .A2(G8), .A3(new_n1085), .A4(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1088), .A2(KEYINPUT123), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1073), .A2(G171), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1078), .B2(G171), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1080), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1041), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1055), .B(KEYINPUT116), .Z(new_n1104));
  AND2_X1   g679(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1089), .A2(G8), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G168), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1104), .A2(new_n1105), .A3(KEYINPUT63), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1064), .B2(new_n1107), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1052), .A2(new_n1043), .A3(new_n788), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1047), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1109), .A2(new_n1111), .B1(new_n1042), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1063), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1104), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1103), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1095), .A2(new_n1118), .A3(new_n1096), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1098), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1064), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1097), .A2(KEYINPUT62), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1119), .A2(KEYINPUT125), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n976), .B1(new_n1117), .B2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n971), .B(KEYINPUT126), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n969), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(G2067), .B2(new_n755), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(new_n965), .ZN(new_n1132));
  INV_X1    g707(.A(G1996), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n965), .A2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1134), .A2(KEYINPUT46), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n965), .B1(new_n967), .B2(new_n729), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(KEYINPUT46), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT47), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n965), .A2(new_n975), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT48), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n972), .A2(new_n965), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT127), .Z(new_n1143));
  AOI211_X1 g718(.A(new_n1132), .B(new_n1139), .C1(new_n1141), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1128), .A2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g720(.A1(G229), .A2(new_n463), .ZN(new_n1147));
  NOR2_X1   g721(.A1(G401), .A2(G227), .ZN(new_n1148));
  NAND4_X1  g722(.A1(new_n867), .A2(new_n957), .A3(new_n1147), .A4(new_n1148), .ZN(G225));
  INV_X1    g723(.A(G225), .ZN(G308));
endmodule


