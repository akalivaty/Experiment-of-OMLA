//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n450), .B(new_n451), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT67), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n464), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT68), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n473), .A2(new_n476), .A3(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n466), .A2(G2105), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n462), .A2(new_n463), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(new_n482), .B2(G137), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n482), .A2(G136), .ZN(new_n486));
  INV_X1    g061(.A(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n467), .B2(new_n469), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n487), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n487), .C1(new_n462), .C2(new_n463), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n464), .A2(new_n470), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n500), .B2(new_n503), .ZN(G164));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n515), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n510), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT69), .B(G51), .Z(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n517), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n525), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n509), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n518), .A2(new_n535), .B1(new_n523), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n509), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n518), .A2(new_n541), .B1(new_n523), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(KEYINPUT70), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n505), .A2(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G81), .B1(new_n514), .B2(G43), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n546), .B(new_n547), .C1(new_n509), .C2(new_n539), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n528), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n514), .B2(G53), .ZN(new_n564));
  OAI221_X1 g139(.A(new_n559), .B1(new_n560), .B2(new_n518), .C1(new_n562), .C2(new_n564), .ZN(G299));
  NOR2_X1   g140(.A1(G171), .A2(KEYINPUT71), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT71), .ZN(new_n567));
  NOR3_X1   g142(.A1(new_n534), .A2(new_n537), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  OAI221_X1 g145(.A(new_n515), .B1(new_n518), .B2(new_n516), .C1(new_n508), .C2(new_n509), .ZN(G303));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n509), .B1(new_n528), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(G49), .B2(new_n514), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n545), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  OAI21_X1  g151(.A(G61), .B1(new_n526), .B2(new_n527), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT72), .B1(new_n579), .B2(G651), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n581));
  AOI211_X1 g156(.A(new_n581), .B(new_n509), .C1(new_n577), .C2(new_n578), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g158(.A1(KEYINPUT6), .A2(G651), .ZN(new_n584));
  NOR2_X1   g159(.A1(KEYINPUT6), .A2(G651), .ZN(new_n585));
  OAI211_X1 g160(.A(G48), .B(G543), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n517), .A2(KEYINPUT73), .A3(G48), .A4(G543), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n588), .A2(new_n589), .B1(new_n545), .B2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n583), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n509), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n545), .A2(G85), .B1(new_n514), .B2(G47), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G290));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n518), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n528), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n597), .B1(new_n518), .B2(new_n596), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G301), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G284));
  AOI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n559), .B1(new_n560), .B2(new_n518), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n562), .A2(new_n564), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n609), .B1(new_n612), .B2(G868), .ZN(G297));
  OAI21_X1  g188(.A(new_n609), .B1(new_n612), .B2(G868), .ZN(G280));
  INV_X1    g189(.A(G860), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n604), .B1(G559), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT75), .ZN(G148));
  NOR2_X1   g192(.A1(new_n604), .A2(G559), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  OR3_X1    g194(.A1(new_n618), .A2(KEYINPUT76), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(KEYINPUT76), .B1(new_n618), .B2(new_n619), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n620), .B(new_n621), .C1(G868), .C2(new_n550), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g198(.A1(new_n464), .A2(new_n470), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n479), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT77), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT78), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n482), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n488), .A2(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n487), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT79), .ZN(new_n638));
  INV_X1    g213(.A(G2096), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n630), .A2(new_n632), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT80), .Z(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(G401));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n628), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n639), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n672), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT81), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n675), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n685), .A2(new_n687), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n689), .B1(new_n688), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G26), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n482), .A2(G140), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n488), .A2(G128), .ZN(new_n698));
  OR2_X1    g273(.A1(G104), .A2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(G2104), .C1(G116), .C2(new_n487), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n696), .B1(new_n702), .B2(new_n694), .ZN(new_n703));
  INV_X1    g278(.A(G2067), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n694), .A2(G32), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT89), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT26), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n488), .A2(G129), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n479), .ZN(new_n711));
  AND3_X1   g286(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n694), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT27), .B(G1996), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(G164), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G27), .B2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G2078), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n705), .A2(new_n716), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n723), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT93), .ZN(new_n727));
  INV_X1    g302(.A(G1966), .ZN(new_n728));
  AND3_X1   g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n727), .B1(new_n726), .B2(new_n728), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n722), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n694), .A2(G35), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G162), .B2(new_n694), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT29), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(G2090), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(G2090), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n723), .A2(G19), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n549), .B2(G16), .ZN(new_n739));
  INV_X1    g314(.A(G1341), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NOR4_X1   g317(.A1(new_n735), .A2(new_n736), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n723), .A2(G20), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT23), .Z(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G299), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1956), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n728), .B2(new_n726), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n723), .A2(G5), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G171), .B2(new_n723), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT94), .B(G1961), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT31), .B(G11), .Z(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT92), .B(G28), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT30), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n754), .B2(KEYINPUT30), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n752), .B(new_n757), .C1(new_n694), .C2(new_n638), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n723), .A2(G4), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(new_n723), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1348), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n748), .A2(new_n758), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n694), .B1(KEYINPUT24), .B2(G34), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(KEYINPUT24), .B2(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n484), .B2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND4_X1   g343(.A1(new_n731), .A2(new_n743), .A3(new_n763), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n624), .A2(G127), .ZN(new_n771));
  NAND2_X1  g346(.A1(G115), .A2(G2104), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n487), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT87), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(KEYINPUT87), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT86), .B(KEYINPUT25), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n487), .A2(G103), .A3(G2104), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n778), .A2(new_n779), .B1(new_n482), .B2(G139), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n774), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G33), .B(new_n781), .S(G29), .Z(new_n782));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n782), .A2(new_n783), .A3(G2072), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n782), .B2(G2072), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n713), .A2(new_n715), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n787), .B1(new_n767), .B2(new_n766), .C1(new_n782), .C2(G2072), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n770), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n788), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(KEYINPUT90), .C1(new_n785), .C2(new_n784), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n769), .A2(new_n789), .A3(new_n791), .A4(KEYINPUT95), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n791), .A2(new_n769), .A3(new_n789), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n723), .A2(G23), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G288), .B2(G16), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT82), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT33), .B(G1976), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n803), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n800), .A2(new_n805), .A3(new_n801), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n723), .A2(G6), .ZN(new_n808));
  INV_X1    g383(.A(G305), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n723), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT32), .B(G1981), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NOR2_X1   g388(.A1(G16), .A2(G22), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G166), .B2(G16), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT83), .B(G1971), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n807), .A2(new_n812), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n723), .A2(G24), .ZN(new_n820));
  INV_X1    g395(.A(G290), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n723), .ZN(new_n822));
  INV_X1    g397(.A(G1986), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n694), .A2(G25), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n482), .A2(G131), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n488), .A2(G119), .ZN(new_n827));
  OR2_X1    g402(.A1(G95), .A2(G2105), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n828), .B(G2104), .C1(G107), .C2(new_n487), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(new_n694), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT35), .B(G1991), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n824), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n819), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT84), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n818), .A2(new_n837), .A3(KEYINPUT34), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n837), .B1(new_n818), .B2(KEYINPUT34), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(KEYINPUT85), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OAI221_X1 g419(.A(new_n836), .B1(KEYINPUT85), .B2(new_n842), .C1(new_n839), .C2(new_n840), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n792), .A2(new_n795), .B1(new_n844), .B2(new_n845), .ZN(G311));
  NAND2_X1  g421(.A1(new_n795), .A2(new_n792), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(G150));
  AOI22_X1  g424(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(new_n509), .ZN(new_n851));
  INV_X1    g426(.A(G93), .ZN(new_n852));
  INV_X1    g427(.A(G55), .ZN(new_n853));
  OAI22_X1  g428(.A1(new_n518), .A2(new_n852), .B1(new_n523), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n615), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT37), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n851), .A2(new_n854), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(new_n544), .A3(new_n548), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n855), .B1(new_n540), .B2(new_n543), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT97), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n760), .A2(G559), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n859), .A2(new_n864), .A3(new_n860), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n863), .B1(new_n862), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT99), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n873));
  OR3_X1    g448(.A1(new_n870), .A2(new_n873), .A3(KEYINPUT39), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n870), .B2(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n615), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n857), .B1(new_n872), .B2(new_n876), .ZN(G145));
  XNOR2_X1  g452(.A(new_n484), .B(new_n638), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n492), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n781), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n774), .A2(new_n775), .A3(KEYINPUT100), .A4(new_n780), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n503), .A2(new_n500), .ZN(new_n883));
  INV_X1    g458(.A(new_n498), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n712), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G164), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n886), .A2(new_n888), .A3(new_n701), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n701), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n881), .B(new_n882), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n702), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n886), .A2(new_n888), .A3(new_n701), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n893), .A2(new_n880), .A3(new_n781), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n626), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n482), .A2(G142), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n488), .A2(G130), .ZN(new_n899));
  OR2_X1    g474(.A1(G106), .A2(G2105), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n900), .B(G2104), .C1(G118), .C2(new_n487), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n902), .A2(KEYINPUT101), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(KEYINPUT101), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n626), .A2(new_n904), .A3(new_n903), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n906), .A2(new_n831), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n831), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n879), .B1(new_n896), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n910), .B1(new_n896), .B2(KEYINPUT103), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n891), .A2(new_n895), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n913), .B1(new_n912), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT102), .B1(new_n896), .B2(new_n910), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n896), .A2(new_n910), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n908), .A2(new_n909), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n921), .A2(new_n891), .A3(new_n895), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(G37), .B1(new_n924), .B2(new_n879), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n918), .A2(KEYINPUT40), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT40), .B1(new_n918), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(G395));
  AND2_X1   g503(.A1(new_n574), .A2(new_n575), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n821), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G290), .A2(G288), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT107), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n809), .A2(G166), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(G305), .A2(G303), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n933), .A2(new_n935), .A3(new_n937), .A4(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n932), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n941), .B(new_n934), .C1(new_n938), .C2(new_n936), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n943), .B1(KEYINPUT108), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(KEYINPUT108), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n945), .B(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n859), .A2(new_n864), .A3(new_n860), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n864), .B1(new_n859), .B2(new_n860), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n618), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n618), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n862), .A2(new_n951), .A3(new_n865), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n760), .B2(G299), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n612), .A2(KEYINPUT105), .A3(new_n604), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n760), .A2(G299), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT41), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT41), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n955), .A2(new_n956), .A3(new_n960), .A4(new_n957), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OR3_X1    g537(.A1(new_n953), .A2(KEYINPUT106), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n953), .A2(new_n958), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n953), .B2(new_n962), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n963), .B(new_n968), .C1(new_n964), .C2(new_n965), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n947), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n947), .A2(new_n969), .ZN(new_n971));
  OAI21_X1  g546(.A(G868), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n858), .A2(new_n619), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(G295));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n973), .ZN(G331));
  OAI21_X1  g550(.A(G168), .B1(new_n566), .B2(new_n568), .ZN(new_n976));
  INV_X1    g551(.A(G171), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G286), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n976), .B(new_n978), .C1(new_n948), .C2(new_n949), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n978), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n862), .A2(new_n980), .A3(new_n865), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n981), .A3(new_n958), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n979), .A2(new_n981), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(new_n962), .ZN(new_n984));
  AOI21_X1  g559(.A(G37), .B1(new_n984), .B2(new_n943), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n940), .A2(new_n942), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n988), .B(new_n982), .C1(new_n983), .C2(new_n962), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n962), .B1(new_n981), .B2(new_n979), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n979), .A2(new_n981), .A3(new_n958), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n943), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G37), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n993), .A2(new_n989), .A3(new_n987), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n994), .A3(new_n989), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n990), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(KEYINPUT44), .A3(new_n995), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(G397));
  INV_X1    g578(.A(G40), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n1004), .B(new_n480), .C1(new_n482), .C2(G137), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n476), .B1(new_n473), .B2(G2105), .ZN(new_n1006));
  AOI211_X1 g581(.A(KEYINPUT68), .B(new_n487), .C1(new_n471), .C2(new_n472), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G164), .B2(G1384), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n701), .B(G2067), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(G1996), .B2(new_n887), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n712), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1011), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT112), .Z(new_n1017));
  NOR2_X1   g592(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n830), .B(new_n833), .Z(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n823), .A3(new_n821), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(G1986), .A3(G290), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT111), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1384), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n885), .A2(KEYINPUT121), .A3(KEYINPUT45), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(KEYINPUT45), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(G164), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1010), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n728), .B1(new_n1032), .B2(new_n1008), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1005), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n475), .B2(new_n477), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n885), .A2(new_n1027), .A3(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1035), .A2(new_n767), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1033), .A2(G168), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G8), .ZN(new_n1041));
  AOI21_X1  g616(.A(G168), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT51), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1044), .A3(G8), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT62), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1384), .B1(new_n883), .B2(new_n884), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1005), .B(new_n1048), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  INV_X1    g625(.A(new_n578), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n507), .B2(G61), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n581), .B1(new_n1052), .B2(new_n509), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n579), .A2(KEYINPUT72), .A3(G651), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n590), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT115), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n583), .A2(new_n1058), .A3(new_n1054), .A4(new_n590), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n590), .B1(new_n509), .B2(new_n1052), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G1981), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1050), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AND4_X1   g640(.A1(KEYINPUT116), .A2(new_n1060), .A3(KEYINPUT49), .A4(new_n1062), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1057), .A2(new_n1059), .B1(G1981), .B2(new_n1061), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT116), .B1(new_n1067), .B2(KEYINPUT49), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1065), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n929), .A2(G1976), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1049), .A2(G8), .A3(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n929), .A2(G1976), .ZN(new_n1072));
  OR3_X1    g647(.A1(new_n1071), .A2(KEYINPUT52), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(KEYINPUT52), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT114), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1071), .A2(new_n1076), .A3(KEYINPUT52), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1069), .A2(new_n1073), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G2090), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1035), .A2(new_n1080), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1081));
  INV_X1    g656(.A(G1971), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1048), .A2(KEYINPUT45), .B1(G164), .B2(new_n1030), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(new_n1008), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n1086));
  INV_X1    g661(.A(G8), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(G166), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(G8), .A3(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1048), .A2(new_n1037), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1008), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1094), .B1(new_n1048), .B2(new_n1095), .ZN(new_n1096));
  NOR4_X1   g671(.A1(G164), .A2(KEYINPUT120), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n1098), .A3(new_n1080), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1087), .B1(new_n1099), .B2(new_n1084), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1091), .B1(new_n1100), .B2(new_n1090), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1079), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1083), .A2(new_n1008), .A3(G2078), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1083), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(new_n719), .A3(new_n1035), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1105), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(KEYINPUT124), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n719), .A2(KEYINPUT53), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1032), .A2(new_n1008), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1114));
  INV_X1    g689(.A(G1961), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1112), .A2(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(G301), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1043), .A2(new_n1118), .A3(new_n1045), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1047), .A2(new_n1102), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n885), .A2(new_n1095), .A3(new_n1027), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT120), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1048), .A2(new_n1037), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1048), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1035), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1083), .A2(new_n1008), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1126), .A2(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(G299), .B(KEYINPUT57), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1121), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1130), .A2(new_n1121), .A3(new_n1132), .ZN(new_n1135));
  INV_X1    g710(.A(G1348), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1038), .A2(new_n1036), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(new_n1008), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1035), .A2(new_n704), .A3(new_n1048), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1140), .A2(new_n604), .ZN(new_n1141));
  AOI21_X1  g716(.A(G1956), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1107), .A2(new_n1035), .A3(new_n1129), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1131), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1134), .A2(new_n1135), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NOR4_X1   g720(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT122), .A4(new_n1131), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1144), .B1(new_n1146), .B2(new_n1133), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1138), .A2(new_n1139), .A3(KEYINPUT60), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT60), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n604), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n760), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(new_n1132), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1144), .A2(new_n1157), .A3(KEYINPUT61), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1083), .A2(new_n1008), .A3(G1996), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT58), .B(G1341), .Z(new_n1160));
  AND2_X1   g735(.A1(new_n1049), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n550), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT59), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1164), .B(new_n550), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1154), .A2(new_n1158), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1145), .B1(new_n1149), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT54), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1115), .B1(new_n1137), .B2(new_n1008), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n474), .A2(new_n1005), .A3(new_n1112), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1083), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  AOI211_X1 g748(.A(new_n606), .B(new_n1173), .C1(new_n1106), .C2(new_n1110), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1169), .B1(new_n1117), .B2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1104), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT124), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1177));
  OAI211_X1 g752(.A(G301), .B(new_n1116), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1173), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1178), .B(KEYINPUT54), .C1(new_n977), .C2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1175), .A2(new_n1102), .A3(new_n1180), .A4(new_n1046), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1120), .B1(new_n1168), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1078), .A2(new_n1073), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1033), .A2(new_n1039), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1184), .A2(G8), .A3(G168), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1090), .B1(new_n1085), .B2(G8), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1091), .A2(KEYINPUT63), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1183), .A2(new_n1187), .A3(new_n1069), .A4(new_n1188), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1079), .A2(new_n1101), .A3(new_n1185), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(KEYINPUT63), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1050), .B(KEYINPUT117), .Z(new_n1192));
  OR2_X1    g767(.A1(G288), .A2(G1976), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT118), .Z(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT116), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1067), .A2(KEYINPUT116), .A3(KEYINPUT49), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1195), .B1(new_n1199), .B2(new_n1065), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1060), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1192), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1085), .A2(G8), .A3(new_n1090), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1069), .A2(new_n1203), .A3(new_n1078), .A4(new_n1073), .ZN(new_n1204));
  AOI21_X1  g779(.A(KEYINPUT119), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1201), .B1(new_n1069), .B2(new_n1194), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1192), .ZN(new_n1207));
  OAI211_X1 g782(.A(new_n1204), .B(KEYINPUT119), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1191), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1026), .B1(new_n1182), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(KEYINPUT46), .B1(new_n1018), .B2(new_n1014), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  AOI211_X1 g789(.A(new_n887), .B(new_n1012), .C1(KEYINPUT46), .C2(new_n1014), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1214), .B1(new_n1011), .B2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1216), .B(KEYINPUT47), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n831), .A2(new_n833), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT125), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1017), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n702), .A2(new_n704), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1222), .A2(new_n1018), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1021), .A2(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1021), .A2(new_n1224), .ZN(new_n1228));
  OAI211_X1 g803(.A(new_n1217), .B(new_n1223), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1211), .A2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g806(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1233));
  OAI21_X1  g807(.A(new_n1233), .B1(new_n691), .B2(new_n692), .ZN(new_n1234));
  AOI21_X1  g808(.A(new_n1234), .B1(new_n918), .B2(new_n925), .ZN(new_n1235));
  AND2_X1   g809(.A1(new_n1235), .A2(new_n999), .ZN(G308));
  NAND2_X1  g810(.A1(new_n1235), .A2(new_n999), .ZN(G225));
endmodule


