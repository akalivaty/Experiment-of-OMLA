//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n610,
    new_n611, new_n612, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n662, new_n665, new_n667, new_n668,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1243, new_n1244;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT64), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT65), .Z(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n463));
  NAND4_X1  g038(.A1(new_n460), .A2(new_n462), .A3(G137), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n461), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(new_n467), .B2(G112), .ZN(new_n477));
  OR3_X1    g052(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n460), .A2(new_n463), .A3(new_n462), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n481), .B(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n483), .A2(new_n486), .A3(new_n467), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n483), .B2(new_n467), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI211_X1 g064(.A(new_n480), .B(new_n485), .C1(new_n489), .C2(G136), .ZN(G162));
  AND2_X1   g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n460), .A2(new_n462), .A3(new_n497), .A4(new_n463), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT3), .B(G2104), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n500), .A2(new_n497), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n495), .B1(new_n499), .B2(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n508), .B(G543), .C1(new_n510), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  AND4_X1   g090(.A1(new_n507), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(G88), .B1(G50), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n507), .A2(G62), .A3(new_n513), .A4(new_n514), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n519), .A2(new_n523), .A3(KEYINPUT73), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n518), .A2(G50), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n507), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n520), .B2(new_n521), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n525), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n524), .A2(new_n532), .ZN(G166));
  NAND2_X1  g108(.A1(new_n513), .A2(new_n514), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n506), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n508), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(G89), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n518), .A2(G51), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n518), .A2(G52), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT74), .B(G90), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n527), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n537), .A2(new_n508), .B1(KEYINPUT5), .B2(new_n506), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(new_n507), .ZN(new_n557));
  INV_X1    g132(.A(G64), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n548), .B1(new_n554), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n552), .A2(new_n553), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n556), .A2(new_n507), .A3(new_n515), .A4(new_n550), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT75), .B1(new_n563), .B2(new_n549), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n560), .B(new_n548), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n561), .A2(new_n566), .ZN(G301));
  INV_X1    g142(.A(G301), .ZN(G171));
  NAND2_X1  g143(.A1(new_n518), .A2(G43), .ZN(new_n569));
  INV_X1    g144(.A(G81), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n527), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n507), .A2(G56), .A3(new_n513), .A4(new_n514), .ZN(new_n573));
  NAND2_X1  g148(.A1(G68), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n530), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT77), .B1(new_n571), .B2(new_n575), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G860), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT78), .ZN(G153));
  AND3_X1   g157(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G36), .ZN(G176));
  NAND2_X1  g159(.A1(G1), .A2(G3), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT8), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(G188));
  NAND3_X1  g162(.A1(new_n556), .A2(G65), .A3(new_n507), .ZN(new_n588));
  NAND2_X1  g163(.A1(G78), .A2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT9), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT9), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n515), .A2(new_n595), .A3(G53), .A4(G543), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n594), .B1(new_n593), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G91), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n527), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n591), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(KEYINPUT80), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n530), .B1(new_n588), .B2(new_n589), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n601), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n605), .B1(new_n607), .B2(new_n599), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n604), .A2(new_n608), .ZN(G299));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n524), .A2(new_n610), .A3(new_n532), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(new_n524), .B2(new_n532), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(G303));
  INV_X1    g188(.A(G74), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n534), .B2(new_n538), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n615), .A2(G651), .B1(G49), .B2(new_n518), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n516), .B2(G87), .ZN(new_n618));
  INV_X1    g193(.A(G87), .ZN(new_n619));
  NOR3_X1   g194(.A1(new_n527), .A2(KEYINPUT82), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n616), .B1(new_n618), .B2(new_n620), .ZN(G288));
  NAND4_X1  g196(.A1(new_n507), .A2(G61), .A3(new_n513), .A4(new_n514), .ZN(new_n622));
  NAND2_X1  g197(.A1(G73), .A2(G543), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(KEYINPUT83), .B1(new_n624), .B2(G651), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n518), .A2(G48), .ZN(new_n626));
  INV_X1    g201(.A(G86), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n527), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n530), .B1(new_n622), .B2(new_n623), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT83), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n631), .ZN(G305));
  NAND2_X1  g207(.A1(new_n539), .A2(G60), .ZN(new_n633));
  NAND2_X1  g208(.A1(G72), .A2(G543), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n530), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT84), .B(G47), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n518), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G85), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n527), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(G290));
  INV_X1    g216(.A(G868), .ZN(new_n642));
  NOR2_X1   g217(.A1(G301), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g218(.A1(new_n556), .A2(G92), .A3(new_n507), .A4(new_n515), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT10), .ZN(new_n645));
  NAND4_X1  g220(.A1(new_n507), .A2(G66), .A3(new_n513), .A4(new_n514), .ZN(new_n646));
  NAND2_X1  g221(.A1(G79), .A2(G543), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G651), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n518), .A2(G54), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(KEYINPUT85), .B1(new_n645), .B2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT10), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n644), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n655));
  AOI22_X1  g230(.A1(new_n648), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT86), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n643), .B1(new_n659), .B2(new_n642), .ZN(G284));
  AOI21_X1  g235(.A(new_n643), .B1(new_n659), .B2(new_n642), .ZN(G321));
  NAND2_X1  g236(.A1(G299), .A2(new_n642), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n642), .B2(G168), .ZN(G297));
  OAI21_X1  g238(.A(new_n662), .B1(new_n642), .B2(G168), .ZN(G280));
  INV_X1    g239(.A(G559), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n659), .B1(new_n665), .B2(G860), .ZN(G148));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G868), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(G868), .B2(new_n580), .ZN(G323));
  XNOR2_X1  g244(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g245(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT88), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G111), .ZN(new_n674));
  AOI22_X1  g249(.A1(new_n671), .A2(new_n672), .B1(new_n674), .B2(G2105), .ZN(new_n675));
  AOI22_X1  g250(.A1(new_n484), .A2(G123), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n487), .A2(new_n488), .ZN(new_n677));
  INV_X1    g252(.A(G135), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(G2096), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(G2096), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT12), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT13), .ZN(new_n684));
  NAND2_X1  g259(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n684), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(KEYINPUT87), .B2(G2100), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n686), .B1(new_n688), .B2(new_n685), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n680), .A2(new_n681), .A3(new_n689), .ZN(G156));
  XNOR2_X1  g265(.A(G2427), .B(G2438), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2430), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT15), .B(G2435), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(KEYINPUT14), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT90), .ZN(new_n697));
  XOR2_X1   g272(.A(G1341), .B(G1348), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G2451), .B(G2454), .Z(new_n700));
  XNOR2_X1  g275(.A(G2443), .B(G2446), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n706), .A3(G14), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G401));
  XOR2_X1   g283(.A(G2084), .B(G2090), .Z(new_n709));
  XNOR2_X1  g284(.A(G2067), .B(G2678), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(KEYINPUT17), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n709), .A2(new_n710), .ZN(new_n713));
  AOI21_X1  g288(.A(KEYINPUT18), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(G2072), .B(G2078), .Z(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n711), .B2(KEYINPUT18), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(G2096), .B(G2100), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(G227));
  XOR2_X1   g294(.A(G1971), .B(G1976), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT19), .ZN(new_n721));
  XOR2_X1   g296(.A(G1956), .B(G2474), .Z(new_n722));
  XOR2_X1   g297(.A(G1961), .B(G1966), .Z(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT20), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n722), .A2(new_n723), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n721), .A2(new_n724), .A3(new_n727), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n726), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(G1991), .B(G1996), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(G1981), .B(G1986), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(G229));
  INV_X1    g313(.A(G16), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n739), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT102), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G1966), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT103), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n739), .A2(G5), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G171), .B2(new_n739), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(G1961), .ZN(new_n747));
  NOR2_X1   g322(.A1(G27), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2078), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT24), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(G34), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n752), .B1(new_n753), .B2(G34), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n475), .A2(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G2084), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n750), .A2(new_n751), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT30), .B(G28), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n759), .A2(new_n752), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n758), .B(new_n762), .C1(new_n751), .C2(new_n750), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n679), .A2(new_n752), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n752), .A2(G32), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n489), .A2(G141), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT26), .Z(new_n769));
  NAND3_X1  g344(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n484), .B2(G129), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n766), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n765), .B1(new_n774), .B2(new_n775), .C1(new_n742), .C2(G1966), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n744), .A2(new_n747), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n752), .A2(G33), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT25), .ZN(new_n779));
  NAND2_X1  g354(.A1(G103), .A2(G2104), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(G2105), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n500), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  INV_X1    g359(.A(G139), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n783), .B1(new_n467), .B2(new_n784), .C1(new_n677), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n778), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2072), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n756), .A2(new_n757), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n774), .B2(new_n775), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT101), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n746), .A2(G1961), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n788), .A2(new_n790), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT101), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n777), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT104), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n777), .A2(new_n796), .A3(KEYINPUT104), .A4(new_n792), .ZN(new_n800));
  NOR2_X1   g375(.A1(G4), .A2(G16), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n659), .B2(G16), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT96), .B(G1348), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n802), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n752), .A2(G35), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G162), .B2(new_n752), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT29), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(G2090), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n752), .A2(G26), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT28), .ZN(new_n811));
  INV_X1    g386(.A(G140), .ZN(new_n812));
  OR3_X1    g387(.A1(new_n677), .A2(KEYINPUT98), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT98), .B1(new_n677), .B2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n816));
  OR3_X1    g391(.A1(KEYINPUT99), .A2(G104), .A3(G2105), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT99), .B1(G104), .B2(G2105), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n484), .B2(G128), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n811), .B1(new_n821), .B2(new_n752), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT100), .B(G2067), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n739), .A2(G20), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT23), .Z(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G299), .B2(G16), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT105), .B(G1956), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n808), .B2(G2090), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n739), .A2(G19), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT97), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n578), .A2(new_n579), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(G16), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(G1341), .Z(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n829), .B2(new_n827), .ZN(new_n837));
  AND4_X1   g412(.A1(new_n809), .A2(new_n824), .A3(new_n831), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n799), .A2(new_n800), .A3(new_n805), .A4(new_n838), .ZN(new_n839));
  MUX2_X1   g414(.A(G23), .B(G288), .S(G16), .Z(new_n840));
  XOR2_X1   g415(.A(KEYINPUT33), .B(G1976), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT93), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT83), .ZN(new_n844));
  AOI211_X1 g419(.A(new_n844), .B(new_n530), .C1(new_n622), .C2(new_n623), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n625), .A2(new_n845), .A3(new_n628), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G16), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G6), .B2(G16), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT32), .B(G1981), .Z(new_n849));
  OR2_X1    g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n843), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(G16), .A2(G22), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G166), .B2(G16), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(G1971), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT34), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n852), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n752), .A2(G25), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n489), .A2(G131), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n862));
  INV_X1    g437(.A(G107), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(G2105), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n484), .B2(G119), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n860), .B1(new_n866), .B2(G29), .ZN(new_n867));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G1991), .Z(new_n868));
  XOR2_X1   g443(.A(new_n867), .B(new_n868), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n739), .A2(G24), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT92), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n640), .B2(new_n739), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G1986), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT94), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n873), .B1(new_n874), .B2(KEYINPUT36), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n857), .A2(new_n859), .A3(new_n869), .A4(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(KEYINPUT36), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n839), .A2(new_n878), .ZN(G311));
  INV_X1    g454(.A(G311), .ZN(G150));
  NAND2_X1  g455(.A1(new_n518), .A2(G55), .ZN(new_n881));
  INV_X1    g456(.A(G93), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n527), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(G80), .A2(G543), .ZN(new_n884));
  INV_X1    g459(.A(G67), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n557), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n886), .B2(G651), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(KEYINPUT106), .B(G860), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(KEYINPUT107), .B(KEYINPUT37), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n659), .A2(G559), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n887), .B1(new_n578), .B2(new_n579), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n887), .A2(new_n576), .A3(new_n572), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(KEYINPUT38), .Z(new_n897));
  XNOR2_X1  g472(.A(new_n893), .B(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT39), .Z(new_n899));
  OAI21_X1  g474(.A(new_n892), .B1(new_n899), .B2(new_n889), .ZN(G145));
  XNOR2_X1  g475(.A(new_n679), .B(new_n475), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(G162), .Z(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n821), .A2(G164), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n815), .A2(new_n820), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n497), .A2(new_n501), .A3(new_n502), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n500), .A2(new_n906), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n907), .B2(new_n495), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n866), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n484), .A2(G130), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n467), .A2(G118), .ZN(new_n913));
  OAI21_X1  g488(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n915), .B1(G142), .B2(new_n489), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(new_n683), .Z(new_n917));
  XNOR2_X1  g492(.A(new_n773), .B(new_n786), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n904), .A2(new_n866), .A3(new_n908), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n918), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n911), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n911), .A2(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n903), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n911), .A2(new_n920), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n919), .A2(new_n921), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n902), .A3(new_n922), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g507(.A1(new_n654), .A2(new_n656), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n604), .B2(new_n608), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n603), .A2(KEYINPUT80), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n607), .A2(new_n605), .A3(new_n599), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n654), .A4(new_n656), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n937), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n896), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n659), .B2(new_n665), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n659), .A2(new_n665), .A3(new_n945), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n948), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n950), .A2(new_n946), .A3(new_n938), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT42), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(G305), .B(G288), .ZN(new_n953));
  NOR2_X1   g528(.A1(G166), .A2(new_n640), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(G166), .A2(new_n640), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n961));
  INV_X1    g536(.A(new_n938), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n947), .A2(new_n948), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n950), .A2(new_n946), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n961), .B(new_n963), .C1(new_n964), .C2(new_n944), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n952), .A2(new_n960), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n960), .B1(new_n952), .B2(new_n965), .ZN(new_n967));
  OAI21_X1  g542(.A(G868), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n888), .A2(new_n642), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(G295));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n969), .ZN(G331));
  OAI21_X1  g546(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT76), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(G286), .A3(new_n565), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(G286), .B1(new_n973), .B2(new_n565), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n945), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n976), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n896), .B1(new_n978), .B2(new_n974), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n944), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n945), .B1(new_n975), .B2(new_n976), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n896), .A3(new_n974), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n938), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n959), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n926), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n938), .A2(KEYINPUT109), .A3(new_n941), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n934), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT109), .B1(new_n938), .B2(new_n941), .ZN(new_n989));
  OAI22_X1  g564(.A1(new_n988), .A2(new_n989), .B1(new_n977), .B2(new_n979), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n959), .B1(new_n990), .B2(new_n983), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT43), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n980), .A2(new_n983), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n960), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n994), .A2(new_n984), .A3(new_n995), .A4(new_n926), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(KEYINPUT44), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n992), .A2(new_n996), .A3(KEYINPUT110), .A4(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n1002));
  INV_X1    g577(.A(new_n985), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n995), .B1(new_n1003), .B2(new_n994), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n985), .A2(new_n991), .A3(KEYINPUT43), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1001), .A2(new_n1006), .ZN(G397));
  NAND4_X1  g582(.A1(G303), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT73), .B1(new_n519), .B2(new_n523), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n529), .A2(new_n531), .A3(new_n525), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT81), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n524), .A2(new_n610), .A3(new_n532), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1011), .A2(KEYINPUT55), .A3(G8), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(G8), .A3(new_n1012), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1008), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n499), .A2(new_n503), .ZN(new_n1021));
  INV_X1    g596(.A(new_n495), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1384), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n907), .B2(new_n495), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(KEYINPUT50), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  INV_X1    g605(.A(G2090), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT114), .B1(new_n1036), .B2(G2090), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT113), .B(G1971), .Z(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1020), .B1(new_n1023), .B2(KEYINPUT45), .ZN(new_n1040));
  OAI211_X1 g615(.A(KEYINPUT45), .B(new_n1026), .C1(new_n907), .C2(new_n495), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1039), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1032), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1019), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1981), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n629), .B2(new_n631), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT117), .B1(new_n846), .B2(new_n1052), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n516), .A2(G86), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(new_n626), .C1(new_n630), .C2(KEYINPUT83), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  NOR4_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n845), .A4(G1981), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1054), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT49), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1051), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n624), .A2(G651), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n844), .ZN(new_n1064));
  INV_X1    g639(.A(new_n628), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(new_n1052), .A3(new_n631), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1058), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n629), .A2(KEYINPUT117), .A3(new_n1052), .A4(new_n631), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1053), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT49), .ZN(new_n1070));
  INV_X1    g645(.A(G1976), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n616), .B(G1976), .C1(new_n618), .C2(new_n620), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(KEYINPUT116), .A3(new_n1050), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1050), .A3(new_n1073), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1073), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT52), .B1(new_n1076), .B2(new_n1051), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1062), .A2(new_n1070), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1048), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT119), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1050), .B1(new_n1069), .B2(KEYINPUT49), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1061), .B(new_n1053), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OR2_X1    g661(.A1(G288), .A2(G1976), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1050), .B(KEYINPUT118), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT45), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(G164), .B2(G1384), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1092), .A2(new_n751), .A3(new_n1020), .A4(new_n1041), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT124), .B(G1961), .Z(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1092), .A2(new_n1099), .A3(new_n1020), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1094), .A2(G2078), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1041), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1033), .B1(new_n1027), .B2(new_n1091), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n1099), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1098), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n973), .A2(new_n1108), .A3(new_n565), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n973), .B2(new_n565), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n561), .B2(new_n566), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1042), .B1(new_n1040), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1092), .A2(KEYINPUT121), .A3(new_n1020), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n1101), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1036), .A2(new_n1096), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n973), .A2(new_n1108), .A3(new_n565), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1112), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1111), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1966), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1041), .B1(new_n1104), .B2(KEYINPUT121), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1115), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1029), .A2(new_n757), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(G168), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G8), .ZN(new_n1128));
  AOI21_X1  g703(.A(G168), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT51), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1131), .A3(G8), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1121), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT122), .B(G1996), .Z(new_n1134));
  NAND4_X1  g709(.A1(new_n1092), .A2(new_n1020), .A3(new_n1041), .A4(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT58), .B(G1341), .Z(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1027), .B2(new_n1033), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n578), .A2(KEYINPUT123), .A3(new_n579), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT59), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n580), .A2(KEYINPUT123), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT60), .B1(new_n652), .B2(new_n657), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n803), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1145));
  INV_X1    g720(.A(G2067), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1020), .A2(new_n1146), .A3(new_n1023), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1140), .A2(new_n1143), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  AND4_X1   g724(.A1(new_n652), .A2(new_n1145), .A3(new_n657), .A4(new_n1147), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n652), .A2(new_n657), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT60), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT56), .B(G2072), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1104), .A2(new_n1041), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(G1956), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1157), .B1(new_n607), .B2(new_n599), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n593), .A2(new_n596), .ZN(new_n1159));
  NOR4_X1   g734(.A1(new_n606), .A2(new_n601), .A3(KEYINPUT57), .A4(new_n1159), .ZN(new_n1160));
  OAI22_X1  g735(.A1(new_n1155), .A2(new_n1156), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(G1956), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1036), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n603), .A2(KEYINPUT57), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1159), .A2(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n607), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .A4(new_n1154), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1161), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1149), .B(new_n1152), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1161), .B1(new_n658), .B2(new_n1148), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n1167), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1133), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1043), .B1(G2090), .B2(new_n1036), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1043), .B(KEYINPUT120), .C1(G2090), .C2(new_n1036), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(G8), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1180), .A2(new_n1008), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1080), .A2(new_n1047), .A3(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1081), .B(new_n1090), .C1(new_n1175), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n1184));
  AOI211_X1 g759(.A(new_n1049), .B(G286), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1080), .A2(new_n1047), .A3(new_n1181), .A4(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1079), .A2(new_n1074), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1187), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1188), .B1(new_n1019), .B2(new_n1046), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1008), .A2(new_n1045), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1190), .A2(KEYINPUT63), .A3(new_n1185), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1184), .A2(new_n1186), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(KEYINPUT126), .B1(new_n1183), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1186), .A2(new_n1184), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1189), .A2(new_n1181), .A3(new_n1174), .A4(new_n1133), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1088), .A2(new_n1089), .B1(new_n1048), .B2(new_n1080), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1182), .ZN(new_n1204));
  AOI21_X1  g779(.A(G301), .B1(new_n1117), .B2(new_n1116), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1193), .A2(new_n1200), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n905), .B(new_n1146), .ZN(new_n1209));
  INV_X1    g784(.A(G1996), .ZN(new_n1210));
  INV_X1    g785(.A(new_n773), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1092), .A2(new_n1033), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n1210), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1214), .B(KEYINPUT112), .ZN(new_n1215));
  AOI22_X1  g790(.A1(new_n1212), .A2(new_n1213), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1216));
  AND2_X1   g791(.A1(new_n910), .A2(new_n868), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n910), .A2(new_n868), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1213), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1213), .ZN(new_n1221));
  NOR2_X1   g796(.A1(G290), .A2(G1986), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT111), .ZN(new_n1223));
  NAND2_X1  g798(.A1(G290), .A2(G1986), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1221), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1220), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1208), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n821), .A2(new_n1146), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1221), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1223), .A2(new_n1221), .ZN(new_n1231));
  XNOR2_X1  g806(.A(new_n1231), .B(KEYINPUT48), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1220), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1215), .B1(KEYINPUT127), .B2(KEYINPUT46), .ZN(new_n1234));
  NAND2_X1  g809(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1235));
  MUX2_X1   g810(.A(new_n1215), .B(new_n1234), .S(new_n1235), .Z(new_n1236));
  NAND2_X1  g811(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1236), .B1(new_n1237), .B2(new_n1213), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n1238), .B(KEYINPUT47), .ZN(new_n1239));
  NOR3_X1   g814(.A1(new_n1230), .A2(new_n1233), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1227), .A2(new_n1240), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g816(.A(G319), .ZN(new_n1243));
  NOR4_X1   g817(.A1(G401), .A2(new_n1243), .A3(G227), .A4(G229), .ZN(new_n1244));
  OAI211_X1 g818(.A(new_n1244), .B(new_n931), .C1(new_n1004), .C2(new_n1005), .ZN(G225));
  INV_X1    g819(.A(G225), .ZN(G308));
endmodule


