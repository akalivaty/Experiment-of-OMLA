//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028;
  AND2_X1   g000(.A1(KEYINPUT68), .A2(G218gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(KEYINPUT68), .A2(G218gat), .ZN(new_n203));
  OAI21_X1  g002(.A(G211gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G211gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT69), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G211gat), .B(G218gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n206), .A2(new_n207), .A3(new_n212), .A4(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n206), .A2(new_n207), .B1(new_n215), .B2(new_n212), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G226gat), .A2(G233gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT27), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT27), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(G190gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT28), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT27), .B(G183gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(KEYINPUT28), .A3(new_n226), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NOR3_X1   g036(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(KEYINPUT66), .B(new_n233), .C1(new_n237), .C2(new_n238), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n243), .A3(new_n228), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n232), .A2(new_n241), .A3(new_n242), .A4(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246));
  INV_X1    g045(.A(G169gat), .ZN(new_n247));
  INV_X1    g046(.A(G176gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT23), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(G190gat), .A3(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(G190gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT23), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n251), .A2(new_n254), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n250), .B1(G169gat), .B2(G176gat), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT64), .A4(new_n234), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT25), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n226), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n255), .B1(new_n263), .B2(new_n252), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n257), .A2(new_n259), .A3(new_n234), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT25), .A4(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT29), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n221), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n220), .B1(new_n245), .B2(new_n267), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n219), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  INV_X1    g072(.A(new_n219), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT29), .B1(new_n245), .B2(new_n267), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n273), .B(new_n274), .C1(new_n221), .C2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT70), .ZN(new_n278));
  XNOR2_X1  g077(.A(G64gat), .B(G92gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n272), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n272), .A2(new_n276), .A3(KEYINPUT30), .A4(new_n280), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n272), .A2(new_n276), .ZN(new_n285));
  INV_X1    g084(.A(new_n280), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G127gat), .B(G134gat), .Z(new_n290));
  XNOR2_X1  g089(.A(G113gat), .B(G120gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(KEYINPUT1), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G113gat), .B(G120gat), .Z(new_n293));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294));
  XNOR2_X1  g093(.A(G127gat), .B(G134gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n292), .A2(new_n296), .A3(KEYINPUT67), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT67), .B1(new_n292), .B2(new_n296), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n268), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n292), .A2(new_n296), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n292), .A2(new_n296), .A3(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(new_n245), .A3(new_n267), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G227gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT34), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT34), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n307), .A2(new_n314), .A3(new_n311), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n306), .A3(new_n310), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT33), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G15gat), .B(G43gat), .Z(new_n319));
  XNOR2_X1  g118(.A(G71gat), .B(G99gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n313), .B(new_n315), .C1(new_n318), .C2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n316), .A2(KEYINPUT32), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n316), .B2(new_n317), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n314), .B1(new_n307), .B2(new_n311), .ZN(new_n326));
  AOI211_X1 g125(.A(KEYINPUT34), .B(new_n310), .C1(new_n300), .C2(new_n306), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n323), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n324), .B1(new_n323), .B2(new_n328), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G228gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(G148gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT73), .B1(new_n333), .B2(G141gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n335));
  INV_X1    g134(.A(G141gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(G148gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n334), .B(new_n337), .C1(new_n336), .C2(G148gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  INV_X1    g138(.A(G155gat), .ZN(new_n340));
  INV_X1    g139(.A(G162gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n339), .B1(new_n342), .B2(KEYINPUT2), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n342), .A2(new_n339), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT71), .B(KEYINPUT2), .Z(new_n346));
  XNOR2_X1  g145(.A(G141gat), .B(G148gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT72), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n345), .B(new_n350), .C1(new_n346), .C2(new_n347), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n344), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n269), .B1(new_n217), .B2(new_n218), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT3), .B1(new_n353), .B2(KEYINPUT78), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n206), .A2(new_n207), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n215), .A2(new_n212), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n357), .B2(new_n216), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n352), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT29), .B1(new_n352), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n274), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n332), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT3), .B1(new_n353), .B2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n358), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n352), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(G228gat), .B(G233gat), .C1(new_n363), .C2(new_n274), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT80), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n338), .A2(new_n343), .ZN(new_n373));
  INV_X1    g172(.A(new_n351), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT71), .B(KEYINPUT2), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n333), .A2(G141gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n336), .A2(G148gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n350), .B1(new_n378), .B2(new_n345), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n373), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n362), .B1(new_n358), .B2(new_n367), .ZN(new_n381));
  AOI211_X1 g180(.A(KEYINPUT79), .B(KEYINPUT29), .C1(new_n357), .C2(new_n216), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n269), .B1(new_n380), .B2(KEYINPUT3), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n332), .B1(new_n384), .B2(new_n219), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n372), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n365), .B1(new_n371), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT31), .B(G50gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT81), .B(G22gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n390), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(new_n365), .C1(new_n371), .C2(new_n386), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n392), .B1(new_n391), .B2(new_n394), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n289), .B(new_n331), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n380), .A2(new_n301), .ZN(new_n400));
  INV_X1    g199(.A(new_n301), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n352), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n399), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n301), .B1(new_n352), .B2(new_n362), .ZN(new_n404));
  AOI211_X1 g203(.A(KEYINPUT3), .B(new_n344), .C1(new_n349), .C2(new_n351), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n398), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n380), .B2(new_n301), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n352), .A2(KEYINPUT4), .A3(new_n304), .A4(new_n303), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(KEYINPUT5), .B(new_n403), .C1(new_n406), .C2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT4), .B1(new_n299), .B2(new_n352), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n380), .A2(new_n407), .A3(new_n301), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n401), .B1(new_n380), .B2(KEYINPUT3), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n352), .A2(new_n362), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n399), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT75), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n420), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n426), .B1(new_n411), .B2(new_n419), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n426), .A3(new_n419), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n428), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT77), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n432), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(KEYINPUT77), .A3(new_n428), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n431), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT35), .B1(new_n397), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n392), .ZN(new_n440));
  INV_X1    g239(.A(new_n394), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT80), .B1(new_n369), .B2(new_n370), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n383), .A2(new_n372), .A3(new_n385), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n393), .B1(new_n444), .B2(new_n365), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n440), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n432), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(new_n428), .A3(new_n433), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT35), .B1(new_n450), .B2(new_n430), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n448), .A2(new_n451), .A3(new_n289), .A4(new_n331), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n439), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n447), .B(new_n446), .C1(new_n438), .C2(new_n288), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n430), .B(new_n281), .C1(new_n434), .C2(new_n432), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT38), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n280), .B1(new_n285), .B2(KEYINPUT37), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n272), .A2(new_n276), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n285), .A2(KEYINPUT37), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n463), .A2(new_n457), .A3(new_n286), .A4(new_n460), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n458), .A2(KEYINPUT83), .A3(new_n457), .A4(new_n460), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n462), .A2(new_n468), .B1(new_n447), .B2(new_n446), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT39), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n407), .B1(new_n305), .B2(new_n380), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n352), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n404), .A2(new_n405), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n471), .B(new_n399), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n426), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n380), .A2(new_n301), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n352), .A2(new_n401), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n398), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT39), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n472), .B(new_n473), .C1(new_n405), .C2(new_n404), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n482), .B2(new_n399), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n470), .B1(new_n477), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n399), .ZN(new_n485));
  INV_X1    g284(.A(new_n481), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n487), .A2(KEYINPUT40), .A3(new_n426), .A4(new_n476), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n288), .A2(new_n484), .A3(new_n449), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n426), .A3(new_n476), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n432), .B1(new_n491), .B2(new_n470), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT82), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n288), .A4(new_n488), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n454), .A2(new_n455), .B1(new_n469), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n456), .ZN(new_n497));
  INV_X1    g296(.A(new_n461), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n468), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n495), .A2(new_n499), .A3(new_n454), .A4(new_n448), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n331), .B(KEYINPUT36), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n453), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G29gat), .ZN(new_n505));
  INV_X1    g304(.A(G36gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G50gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G43gat), .ZN(new_n515));
  INV_X1    g314(.A(G43gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G50gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n517), .A3(KEYINPUT15), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT87), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n510), .A2(new_n509), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT14), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(new_n505), .A3(new_n506), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n512), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n507), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n510), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n528), .A2(new_n518), .A3(new_n524), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530));
  OR2_X1    g329(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n532));
  AOI21_X1  g331(.A(G50gat), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n514), .B2(G43gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n516), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n530), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n529), .A2(new_n538), .A3(KEYINPUT90), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT90), .B1(new_n529), .B2(new_n538), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n519), .B(new_n527), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n516), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT89), .B1(new_n516), .B2(G50gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n532), .ZN(new_n548));
  NOR2_X1   g347(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n514), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT15), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n528), .A2(new_n518), .A3(new_n524), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n544), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n529), .A2(new_n538), .A3(KEYINPUT90), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n555), .A2(KEYINPUT91), .A3(new_n519), .A4(new_n527), .ZN(new_n556));
  XOR2_X1   g355(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n557));
  NAND3_X1  g356(.A1(new_n543), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n555), .A2(KEYINPUT17), .A3(new_n519), .A4(new_n527), .ZN(new_n559));
  XNOR2_X1  g358(.A(G15gat), .B(G22gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT16), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(G1gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(G1gat), .B2(new_n560), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(G8gat), .Z(new_n564));
  AND2_X1   g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n564), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n543), .A2(new_n556), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT93), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n566), .A2(KEYINPUT93), .A3(new_n567), .A4(new_n569), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT94), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n566), .A2(KEYINPUT18), .A3(new_n567), .A4(new_n569), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n567), .B(KEYINPUT13), .Z(new_n578));
  INV_X1    g377(.A(new_n569), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n568), .B1(new_n543), .B2(new_n556), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT85), .B(G197gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT11), .B(G169gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT12), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT18), .B1(new_n570), .B2(new_n571), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n582), .B1(new_n593), .B2(new_n574), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n593), .B2(new_n574), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n596), .B2(new_n590), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT95), .B1(new_n592), .B2(new_n597), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n559), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G99gat), .B(G106gat), .Z(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n606), .B2(new_n610), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n543), .A2(new_n556), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI211_X1 g417(.A(new_n604), .B(new_n616), .C1(new_n618), .C2(new_n557), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n616), .ZN(new_n620));
  NAND3_X1  g419(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT98), .ZN(new_n624));
  OR3_X1    g423(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n624), .B1(new_n619), .B2(new_n622), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n625), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n625), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G57gat), .B(G64gat), .Z(new_n633));
  INV_X1    g432(.A(KEYINPUT9), .ZN(new_n634));
  INV_X1    g433(.A(G71gat), .ZN(new_n635));
  INV_X1    g434(.A(G78gat), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G71gat), .B(G78gat), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n637), .B(new_n633), .C1(new_n641), .C2(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(KEYINPUT21), .ZN(new_n646));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(G127gat), .Z(new_n649));
  AOI21_X1  g448(.A(new_n568), .B1(KEYINPUT21), .B2(new_n645), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G183gat), .B(G211gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT97), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n340), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n654), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n632), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT100), .ZN(new_n663));
  INV_X1    g462(.A(new_n613), .ZN(new_n664));
  INV_X1    g463(.A(new_n615), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n645), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT10), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n644), .B(new_n643), .C1(new_n613), .C2(new_n615), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n616), .A2(KEYINPUT10), .A3(new_n645), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n663), .B1(new_n671), .B2(KEYINPUT99), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT99), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT101), .ZN(new_n677));
  XNOR2_X1  g476(.A(G176gat), .B(G204gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n666), .A2(new_n668), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(new_n663), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n663), .ZN(new_n683));
  MUX2_X1   g482(.A(new_n680), .B(new_n671), .S(new_n683), .Z(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n679), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n661), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n504), .A2(new_n603), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n438), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n288), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT16), .B(G8gat), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT42), .Z(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(G8gat), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT102), .Z(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1325gat));
  AOI21_X1  g497(.A(G15gat), .B1(new_n689), .B2(new_n331), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT103), .ZN(new_n700));
  INV_X1    g499(.A(new_n501), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(G15gat), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n689), .B2(new_n702), .ZN(G1326gat));
  NOR2_X1   g502(.A1(new_n395), .A2(new_n396), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT43), .B(G22gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  AND3_X1   g506(.A1(new_n495), .A2(new_n499), .A3(new_n448), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n433), .A2(KEYINPUT77), .A3(new_n428), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT77), .B1(new_n433), .B2(new_n428), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n709), .A2(new_n710), .A3(new_n432), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n289), .B1(new_n711), .B2(new_n431), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT84), .B1(new_n712), .B2(new_n704), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n501), .B(new_n500), .C1(new_n708), .C2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n603), .B1(new_n714), .B2(new_n453), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n660), .A2(new_n687), .ZN(new_n716));
  INV_X1    g515(.A(new_n632), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n438), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n719), .A2(G29gat), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT45), .Z(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  INV_X1    g522(.A(new_n598), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n716), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n726));
  AOI211_X1 g525(.A(new_n717), .B(new_n726), .C1(new_n714), .C2(new_n453), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n503), .B2(new_n632), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n725), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT105), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n733), .B(new_n725), .C1(new_n727), .C2(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n723), .B1(new_n735), .B2(new_n720), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G29gat), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n735), .A2(new_n723), .A3(new_n720), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n722), .B1(new_n737), .B2(new_n738), .ZN(G1328gat));
  OAI21_X1  g538(.A(G36gat), .B1(new_n735), .B2(new_n289), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n719), .A2(G36gat), .A3(new_n289), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1329gat));
  INV_X1    g542(.A(new_n331), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n531), .A2(new_n532), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n719), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n731), .B2(new_n501), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT47), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n701), .A3(new_n734), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n746), .B1(new_n750), .B2(new_n745), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n751), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n704), .A3(new_n734), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G50gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n448), .A2(G50gat), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n503), .A2(new_n602), .A3(new_n718), .A4(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n763));
  OAI21_X1  g562(.A(G50gat), .B1(new_n731), .B2(new_n448), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n759), .B1(new_n764), .B2(new_n756), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n760), .B1(new_n753), .B2(G50gat), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT108), .B1(new_n768), .B2(new_n765), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1331gat));
  NAND3_X1  g569(.A1(new_n661), .A2(new_n724), .A3(new_n686), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n504), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n438), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g573(.A(new_n772), .B(KEYINPUT109), .Z(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n288), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT49), .B(G64gat), .Z(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n776), .B2(new_n778), .ZN(G1333gat));
  NAND3_X1  g578(.A1(new_n775), .A2(G71gat), .A3(new_n701), .ZN(new_n780));
  INV_X1    g579(.A(new_n772), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n635), .B1(new_n781), .B2(new_n744), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n780), .A2(KEYINPUT50), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT50), .B1(new_n780), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(G1334gat));
  NAND2_X1  g584(.A1(new_n775), .A2(new_n704), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G78gat), .ZN(G1335gat));
  INV_X1    g586(.A(new_n660), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n598), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT110), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n790), .A2(KEYINPUT51), .A3(new_n503), .A4(new_n632), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT111), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n504), .A2(new_n717), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT51), .A4(new_n790), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n790), .A2(new_n503), .A3(new_n632), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n792), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n799), .A2(new_n608), .A3(new_n438), .A4(new_n686), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n686), .B(new_n790), .C1(new_n727), .C2(new_n730), .ZN(new_n801));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801), .B2(new_n720), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1336gat));
  NAND2_X1  g602(.A1(new_n798), .A2(new_n791), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n687), .A2(new_n289), .A3(G92gat), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT112), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT113), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n804), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  OAI21_X1  g609(.A(G92gat), .B1(new_n801), .B2(new_n289), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT52), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n799), .A2(KEYINPUT114), .A3(new_n805), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT114), .B1(new_n799), .B2(new_n805), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n814), .B(new_n811), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n813), .A2(new_n817), .ZN(G1337gat));
  NOR3_X1   g617(.A1(new_n744), .A2(G99gat), .A3(new_n687), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n799), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G99gat), .B1(new_n801), .B2(new_n501), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1338gat));
  OR2_X1    g621(.A1(new_n801), .A2(new_n448), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  XNOR2_X1  g623(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n448), .A2(G106gat), .A3(new_n687), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n799), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n823), .A2(G106gat), .B1(new_n804), .B2(new_n827), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n826), .A2(new_n828), .B1(new_n829), .B2(new_n830), .ZN(G1339gat));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n688), .A2(new_n598), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n575), .A2(new_n590), .A3(new_n583), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n567), .B1(new_n566), .B2(new_n569), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n579), .A2(new_n580), .A3(new_n578), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n589), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n669), .A2(new_n663), .A3(new_n670), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n672), .B2(new_n674), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n671), .A2(new_n844), .A3(new_n683), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n679), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n842), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n675), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT116), .B1(new_n849), .B2(KEYINPUT55), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  NOR4_X1   g650(.A1(new_n843), .A2(new_n846), .A3(new_n851), .A4(new_n840), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n682), .B(new_n847), .C1(new_n850), .C2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n632), .A2(new_n839), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n594), .A2(new_n596), .A3(new_n590), .ZN(new_n857));
  AOI221_X4 g656(.A(new_n582), .B1(new_n595), .B2(new_n591), .C1(new_n574), .C2(new_n593), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n835), .A2(new_n838), .A3(new_n686), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n632), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(KEYINPUT117), .A3(new_n861), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n856), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n834), .B1(new_n866), .B2(new_n788), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n704), .A2(new_n744), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n867), .A2(KEYINPUT118), .A3(new_n438), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n853), .B1(new_n592), .B2(new_n597), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n863), .B1(new_n870), .B2(new_n860), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n865), .A2(new_n871), .A3(new_n717), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n788), .B1(new_n872), .B2(new_n855), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n438), .B(new_n868), .C1(new_n873), .C2(new_n833), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n288), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877), .B2(new_n598), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n867), .A2(new_n438), .A3(new_n289), .A4(new_n868), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(G113gat), .A3(new_n602), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n832), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n288), .B(new_n724), .C1(new_n869), .C2(new_n876), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT119), .B(new_n881), .C1(new_n884), .C2(G113gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1340gat));
  INV_X1    g685(.A(G120gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n879), .A2(new_n887), .A3(new_n687), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n877), .A2(new_n686), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n887), .ZN(G1341gat));
  AND3_X1   g689(.A1(new_n880), .A2(G127gat), .A3(new_n788), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n288), .B(new_n660), .C1(new_n869), .C2(new_n876), .ZN(new_n892));
  AOI21_X1  g691(.A(G127gat), .B1(new_n892), .B2(KEYINPUT120), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n788), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n891), .B1(new_n893), .B2(new_n896), .ZN(G1342gat));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n879), .B2(new_n717), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n717), .A2(G134gat), .A3(new_n288), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n869), .B2(new_n876), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT56), .B(new_n901), .C1(new_n869), .C2(new_n876), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n898), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n874), .A2(new_n875), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n874), .A2(new_n875), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n900), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n902), .A2(new_n903), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n910), .A2(KEYINPUT121), .A3(new_n911), .A4(new_n899), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n906), .A2(new_n912), .ZN(G1343gat));
  INV_X1    g712(.A(KEYINPUT57), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n867), .A2(new_n914), .A3(new_n704), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n701), .A2(new_n720), .A3(new_n288), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n917));
  INV_X1    g716(.A(new_n601), .ZN(new_n918));
  INV_X1    g717(.A(new_n682), .ZN(new_n919));
  INV_X1    g718(.A(new_n846), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n671), .A2(KEYINPUT99), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(new_n683), .A3(new_n674), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n920), .B(KEYINPUT55), .C1(new_n922), .C2(new_n842), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n851), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n849), .A2(KEYINPUT116), .A3(KEYINPUT55), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n849), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT122), .B1(new_n843), .B2(new_n846), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n929), .A3(new_n840), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n926), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n632), .B1(new_n935), .B2(new_n861), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n660), .B1(new_n936), .B2(new_n856), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n448), .B1(new_n937), .B2(new_n834), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n915), .B(new_n916), .C1(new_n938), .C2(new_n914), .ZN(new_n939));
  OAI21_X1  g738(.A(G141gat), .B1(new_n939), .B2(new_n603), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n873), .A2(new_n833), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(new_n720), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n701), .A2(new_n288), .A3(new_n448), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n603), .A2(G141gat), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT58), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n944), .A2(G141gat), .A3(new_n603), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n950), .A2(new_n600), .A3(new_n601), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n717), .B1(new_n951), .B2(new_n860), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n788), .B1(new_n952), .B2(new_n855), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n704), .B1(new_n953), .B2(new_n833), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT57), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n955), .A2(new_n598), .A3(new_n915), .A4(new_n916), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n949), .B1(new_n956), .B2(G141gat), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT58), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n948), .B1(new_n957), .B2(new_n958), .ZN(G1344gat));
  NAND3_X1  g758(.A1(new_n945), .A2(new_n333), .A3(new_n686), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT59), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G148gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n939), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n686), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n688), .A2(new_n602), .A3(KEYINPUT124), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT124), .B1(new_n688), .B2(new_n602), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n914), .B(new_n704), .C1(new_n953), .C2(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(KEYINPUT57), .B1(new_n941), .B2(new_n448), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n968), .A2(new_n686), .A3(new_n916), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n961), .B1(new_n970), .B2(G148gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n960), .B1(new_n964), .B2(new_n971), .ZN(G1345gat));
  OAI21_X1  g771(.A(G155gat), .B1(new_n939), .B2(new_n660), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n945), .A2(new_n340), .A3(new_n788), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1346gat));
  OAI21_X1  g774(.A(G162gat), .B1(new_n939), .B2(new_n717), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n945), .A2(new_n341), .A3(new_n632), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1347gat));
  NOR2_X1   g777(.A1(new_n438), .A2(new_n289), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n868), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n941), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(G169gat), .B1(new_n981), .B2(new_n598), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n603), .A2(new_n247), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n981), .B2(new_n983), .ZN(G1348gat));
  NAND2_X1  g783(.A1(new_n981), .A2(new_n686), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g785(.A1(new_n981), .A2(new_n788), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n987), .A2(new_n230), .ZN(new_n988));
  NAND2_X1  g787(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n222), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n989), .B1(new_n988), .B2(new_n990), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(G1350gat));
  NOR2_X1   g792(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n994), .B1(new_n981), .B2(new_n632), .ZN(new_n995));
  NAND2_X1  g794(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n996));
  XOR2_X1   g795(.A(new_n995), .B(new_n996), .Z(G1351gat));
  NOR2_X1   g796(.A1(new_n941), .A2(new_n448), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n501), .A2(new_n979), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(G197gat), .B1(new_n1001), .B2(new_n598), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n968), .A2(new_n969), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n1003), .A2(new_n999), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n602), .A2(G197gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(G1352gat));
  OR2_X1    g805(.A1(new_n687), .A2(G204gat), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT62), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1003), .A2(new_n686), .A3(new_n999), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(G204gat), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1353gat));
  NAND4_X1  g811(.A1(new_n968), .A2(new_n788), .A3(new_n969), .A4(new_n999), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(G211gat), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1014), .A2(KEYINPUT63), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT63), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1013), .A2(new_n1016), .A3(G211gat), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n788), .A2(new_n208), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n1000), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n1019), .A2(KEYINPUT126), .ZN(new_n1020));
  AND2_X1   g819(.A1(new_n1019), .A2(KEYINPUT126), .ZN(new_n1021));
  OAI211_X1 g820(.A(new_n1015), .B(new_n1017), .C1(new_n1020), .C2(new_n1021), .ZN(G1354gat));
  NOR2_X1   g821(.A1(new_n202), .A2(new_n203), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n717), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n210), .B1(new_n1000), .B2(new_n717), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1025), .A2(KEYINPUT127), .ZN(new_n1026));
  INV_X1    g825(.A(KEYINPUT127), .ZN(new_n1027));
  OAI211_X1 g826(.A(new_n1027), .B(new_n210), .C1(new_n1000), .C2(new_n717), .ZN(new_n1028));
  AOI22_X1  g827(.A1(new_n1004), .A2(new_n1024), .B1(new_n1026), .B2(new_n1028), .ZN(G1355gat));
endmodule


