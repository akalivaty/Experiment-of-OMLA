

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590;

  XNOR2_X1 U322 ( .A(n410), .B(KEYINPUT48), .ZN(n411) );
  XNOR2_X1 U323 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U324 ( .A(n414), .B(KEYINPUT121), .ZN(n415) );
  XNOR2_X1 U325 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U326 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U327 ( .A(n402), .B(KEYINPUT107), .ZN(n403) );
  XNOR2_X1 U328 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U329 ( .A(G22GAT), .B(G155GAT), .Z(n427) );
  XNOR2_X1 U330 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n384) );
  XNOR2_X1 U331 ( .A(n447), .B(n384), .ZN(n385) );
  XNOR2_X1 U332 ( .A(n412), .B(n411), .ZN(n537) );
  INV_X1 U333 ( .A(KEYINPUT72), .ZN(n362) );
  INV_X1 U334 ( .A(KEYINPUT33), .ZN(n390) );
  XNOR2_X1 U335 ( .A(n363), .B(n362), .ZN(n364) );
  NOR2_X1 U336 ( .A1(n525), .A2(n417), .ZN(n577) );
  XNOR2_X1 U337 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U338 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U339 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n291) );
  XNOR2_X1 U341 ( .A(KEYINPUT87), .B(KEYINPUT4), .ZN(n290) );
  XNOR2_X1 U342 ( .A(n291), .B(n290), .ZN(n310) );
  XOR2_X1 U343 ( .A(G85GAT), .B(G155GAT), .Z(n293) );
  XNOR2_X1 U344 ( .A(G120GAT), .B(G148GAT), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U346 ( .A(KEYINPUT5), .B(KEYINPUT85), .Z(n295) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(G57GAT), .ZN(n294) );
  XNOR2_X1 U348 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U349 ( .A(n297), .B(n296), .Z(n303) );
  XNOR2_X1 U350 ( .A(G134GAT), .B(G127GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n298), .B(KEYINPUT0), .ZN(n445) );
  XOR2_X1 U352 ( .A(G162GAT), .B(n445), .Z(n300) );
  NAND2_X1 U353 ( .A1(G225GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U355 ( .A(G29GAT), .B(n301), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U357 ( .A(n304), .B(KEYINPUT86), .Z(n308) );
  XOR2_X1 U358 ( .A(KEYINPUT82), .B(KEYINPUT3), .Z(n306) );
  XNOR2_X1 U359 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n419) );
  XNOR2_X1 U361 ( .A(G1GAT), .B(n419), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n497) );
  INV_X1 U364 ( .A(n497), .ZN(n525) );
  XOR2_X1 U365 ( .A(G183GAT), .B(KEYINPUT19), .Z(n312) );
  XNOR2_X1 U366 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n446) );
  XOR2_X1 U368 ( .A(n446), .B(KEYINPUT88), .Z(n314) );
  NAND2_X1 U369 ( .A1(G226GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U371 ( .A(G36GAT), .B(G190GAT), .Z(n330) );
  XOR2_X1 U372 ( .A(n315), .B(n330), .Z(n319) );
  XOR2_X1 U373 ( .A(G169GAT), .B(G8GAT), .Z(n379) );
  XOR2_X1 U374 ( .A(G64GAT), .B(G92GAT), .Z(n317) );
  XNOR2_X1 U375 ( .A(G176GAT), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n317), .B(n316), .ZN(n383) );
  XNOR2_X1 U377 ( .A(n379), .B(n383), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n325) );
  XNOR2_X1 U379 ( .A(G211GAT), .B(KEYINPUT80), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n320), .B(KEYINPUT21), .ZN(n321) );
  XOR2_X1 U381 ( .A(n321), .B(KEYINPUT81), .Z(n323) );
  XNOR2_X1 U382 ( .A(G197GAT), .B(G218GAT), .ZN(n322) );
  XOR2_X1 U383 ( .A(n323), .B(n322), .Z(n423) );
  INV_X1 U384 ( .A(n423), .ZN(n324) );
  XOR2_X1 U385 ( .A(n325), .B(n324), .Z(n500) );
  INV_X1 U386 ( .A(n500), .ZN(n527) );
  XOR2_X1 U387 ( .A(KEYINPUT119), .B(n527), .Z(n413) );
  XOR2_X1 U388 ( .A(G29GAT), .B(G43GAT), .Z(n327) );
  XNOR2_X1 U389 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n326) );
  XNOR2_X1 U390 ( .A(n327), .B(n326), .ZN(n368) );
  XNOR2_X1 U391 ( .A(n368), .B(KEYINPUT9), .ZN(n346) );
  XOR2_X1 U392 ( .A(KEYINPUT10), .B(G92GAT), .Z(n329) );
  XNOR2_X1 U393 ( .A(G134GAT), .B(G106GAT), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n334) );
  XOR2_X1 U395 ( .A(G99GAT), .B(G85GAT), .Z(n386) );
  XNOR2_X1 U396 ( .A(n386), .B(n330), .ZN(n332) );
  AND2_X1 U397 ( .A1(G232GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U398 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U399 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U400 ( .A(G50GAT), .B(G162GAT), .Z(n418) );
  XOR2_X1 U401 ( .A(KEYINPUT70), .B(KEYINPUT64), .Z(n336) );
  XNOR2_X1 U402 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n418), .B(n337), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n341) );
  INV_X1 U406 ( .A(KEYINPUT69), .ZN(n340) );
  NAND2_X1 U407 ( .A1(n341), .A2(n340), .ZN(n344) );
  INV_X1 U408 ( .A(n341), .ZN(n342) );
  NAND2_X1 U409 ( .A1(n342), .A2(KEYINPUT69), .ZN(n343) );
  NAND2_X1 U410 ( .A1(n344), .A2(n343), .ZN(n345) );
  XOR2_X1 U411 ( .A(n346), .B(n345), .Z(n401) );
  INV_X1 U412 ( .A(n401), .ZN(n454) );
  XOR2_X1 U413 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n348) );
  XNOR2_X1 U414 ( .A(G8GAT), .B(G64GAT), .ZN(n347) );
  XNOR2_X1 U415 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U416 ( .A(G183GAT), .B(G127GAT), .Z(n350) );
  XNOR2_X1 U417 ( .A(G15GAT), .B(G71GAT), .ZN(n349) );
  XNOR2_X1 U418 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U419 ( .A(n352), .B(n351), .ZN(n367) );
  XOR2_X1 U420 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n354) );
  XNOR2_X1 U421 ( .A(KEYINPUT71), .B(KEYINPUT15), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U423 ( .A(n427), .B(G78GAT), .Z(n356) );
  XOR2_X1 U424 ( .A(G1GAT), .B(KEYINPUT66), .Z(n371) );
  XNOR2_X1 U425 ( .A(n371), .B(G211GAT), .ZN(n355) );
  XNOR2_X1 U426 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U427 ( .A(n358), .B(n357), .Z(n360) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n365) );
  XNOR2_X1 U430 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n361), .B(KEYINPUT67), .ZN(n382) );
  XNOR2_X1 U432 ( .A(n382), .B(KEYINPUT73), .ZN(n363) );
  XOR2_X1 U433 ( .A(n367), .B(n366), .Z(n585) );
  INV_X1 U434 ( .A(n585), .ZN(n571) );
  XOR2_X1 U435 ( .A(n368), .B(KEYINPUT29), .Z(n370) );
  NAND2_X1 U436 ( .A1(G229GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n372) );
  XOR2_X1 U438 ( .A(n372), .B(n371), .Z(n374) );
  XNOR2_X1 U439 ( .A(G50GAT), .B(G36GAT), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U441 ( .A(KEYINPUT30), .B(G141GAT), .Z(n376) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(G22GAT), .ZN(n375) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n381) );
  XOR2_X1 U445 ( .A(G113GAT), .B(G15GAT), .Z(n448) );
  XOR2_X1 U446 ( .A(n448), .B(n379), .Z(n380) );
  XNOR2_X1 U447 ( .A(n381), .B(n380), .ZN(n568) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n395) );
  XOR2_X1 U449 ( .A(G120GAT), .B(G71GAT), .Z(n447) );
  XOR2_X1 U450 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U451 ( .A1(G230GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n388), .B(n387), .ZN(n393) );
  XNOR2_X1 U453 ( .A(G106GAT), .B(G78GAT), .ZN(n389) );
  XNOR2_X1 U454 ( .A(n389), .B(G148GAT), .ZN(n431) );
  XNOR2_X1 U455 ( .A(n431), .B(KEYINPUT68), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n582) );
  XNOR2_X1 U457 ( .A(n582), .B(KEYINPUT41), .ZN(n556) );
  NOR2_X1 U458 ( .A1(n568), .A2(n556), .ZN(n397) );
  XOR2_X1 U459 ( .A(KEYINPUT46), .B(KEYINPUT106), .Z(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n398) );
  NAND2_X1 U461 ( .A1(n571), .A2(n398), .ZN(n399) );
  NOR2_X1 U462 ( .A1(n454), .A2(n399), .ZN(n400) );
  XNOR2_X1 U463 ( .A(KEYINPUT47), .B(n400), .ZN(n409) );
  XOR2_X1 U464 ( .A(KEYINPUT36), .B(n401), .Z(n588) );
  NAND2_X1 U465 ( .A1(n585), .A2(n588), .ZN(n404) );
  INV_X1 U466 ( .A(KEYINPUT45), .ZN(n402) );
  NOR2_X1 U467 ( .A1(n582), .A2(n405), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n406), .B(KEYINPUT108), .ZN(n407) );
  NAND2_X1 U469 ( .A1(n407), .A2(n568), .ZN(n408) );
  NAND2_X1 U470 ( .A1(n409), .A2(n408), .ZN(n412) );
  INV_X1 U471 ( .A(KEYINPUT109), .ZN(n410) );
  NAND2_X1 U472 ( .A1(n413), .A2(n537), .ZN(n416) );
  XOR2_X1 U473 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n414) );
  XOR2_X1 U474 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U477 ( .A(n423), .B(n422), .Z(n435) );
  XOR2_X1 U478 ( .A(KEYINPUT22), .B(KEYINPUT83), .Z(n425) );
  XNOR2_X1 U479 ( .A(KEYINPUT24), .B(KEYINPUT84), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U481 ( .A(n426), .B(G204GAT), .Z(n429) );
  XNOR2_X1 U482 ( .A(n427), .B(KEYINPUT78), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U484 ( .A(n430), .B(KEYINPUT79), .Z(n433) );
  XNOR2_X1 U485 ( .A(n431), .B(KEYINPUT23), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n471) );
  NAND2_X1 U488 ( .A1(n577), .A2(n471), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n436), .B(KEYINPUT55), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n437), .B(KEYINPUT122), .ZN(n453) );
  INV_X1 U491 ( .A(G190GAT), .ZN(n455) );
  XOR2_X1 U492 ( .A(G176GAT), .B(G190GAT), .Z(n439) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(G99GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n442) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n440), .B(KEYINPUT77), .ZN(n441) );
  XOR2_X1 U497 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n452) );
  XOR2_X1 U500 ( .A(n446), .B(n445), .Z(n450) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U503 ( .A(n452), .B(n451), .Z(n502) );
  INV_X1 U504 ( .A(n502), .ZN(n536) );
  NAND2_X1 U505 ( .A1(n453), .A2(n536), .ZN(n570) );
  INV_X1 U506 ( .A(n454), .ZN(n564) );
  NOR2_X1 U507 ( .A1(n570), .A2(n564), .ZN(n458) );
  XNOR2_X1 U508 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n456) );
  XNOR2_X1 U509 ( .A(KEYINPUT98), .B(n556), .ZN(n544) );
  NOR2_X1 U510 ( .A1(n544), .A2(n570), .ZN(n462) );
  XOR2_X1 U511 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n460) );
  XNOR2_X1 U512 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n462), .B(n461), .ZN(G1349GAT) );
  NAND2_X1 U515 ( .A1(n536), .A2(n527), .ZN(n463) );
  NAND2_X1 U516 ( .A1(n471), .A2(n463), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n464), .B(KEYINPUT25), .ZN(n467) );
  XOR2_X1 U518 ( .A(n527), .B(KEYINPUT27), .Z(n470) );
  NOR2_X1 U519 ( .A1(n536), .A2(n471), .ZN(n465) );
  XOR2_X1 U520 ( .A(n465), .B(KEYINPUT26), .Z(n575) );
  NOR2_X1 U521 ( .A1(n470), .A2(n575), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n525), .A2(n468), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT89), .B(n469), .Z(n475) );
  NOR2_X1 U525 ( .A1(n497), .A2(n470), .ZN(n538) );
  XOR2_X1 U526 ( .A(n471), .B(KEYINPUT65), .Z(n472) );
  XOR2_X1 U527 ( .A(KEYINPUT28), .B(n472), .Z(n531) );
  INV_X1 U528 ( .A(n531), .ZN(n535) );
  NAND2_X1 U529 ( .A1(n538), .A2(n535), .ZN(n473) );
  NOR2_X1 U530 ( .A1(n536), .A2(n473), .ZN(n474) );
  NOR2_X1 U531 ( .A1(n475), .A2(n474), .ZN(n491) );
  NAND2_X1 U532 ( .A1(n585), .A2(n564), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(KEYINPUT16), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n477), .B(KEYINPUT76), .ZN(n478) );
  NOR2_X1 U535 ( .A1(n491), .A2(n478), .ZN(n479) );
  XNOR2_X1 U536 ( .A(KEYINPUT90), .B(n479), .ZN(n509) );
  NOR2_X1 U537 ( .A1(n568), .A2(n582), .ZN(n494) );
  NAND2_X1 U538 ( .A1(n509), .A2(n494), .ZN(n480) );
  XOR2_X1 U539 ( .A(KEYINPUT91), .B(n480), .Z(n489) );
  NOR2_X1 U540 ( .A1(n497), .A2(n489), .ZN(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U543 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  NOR2_X1 U544 ( .A1(n500), .A2(n489), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G8GAT), .B(KEYINPUT93), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  NOR2_X1 U547 ( .A1(n502), .A2(n489), .ZN(n487) );
  XNOR2_X1 U548 ( .A(KEYINPUT35), .B(KEYINPUT94), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n535), .A2(n489), .ZN(n490) );
  XOR2_X1 U552 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(KEYINPUT95), .Z(n496) );
  NOR2_X1 U554 ( .A1(n491), .A2(n585), .ZN(n492) );
  NAND2_X1 U555 ( .A1(n588), .A2(n492), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n493), .B(KEYINPUT37), .ZN(n522) );
  NAND2_X1 U557 ( .A1(n522), .A2(n494), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n506) );
  NOR2_X1 U559 ( .A1(n506), .A2(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n500), .A2(n506), .ZN(n501) );
  XOR2_X1 U563 ( .A(G36GAT), .B(n501), .Z(G1329GAT) );
  XNOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT96), .ZN(n504) );
  NOR2_X1 U565 ( .A1(n502), .A2(n506), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U567 ( .A(G43GAT), .B(n505), .Z(G1330GAT) );
  NOR2_X1 U568 ( .A1(n506), .A2(n535), .ZN(n508) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(KEYINPUT97), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(G1331GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT100), .B(KEYINPUT42), .Z(n512) );
  INV_X1 U572 ( .A(n568), .ZN(n579) );
  NOR2_X1 U573 ( .A1(n544), .A2(n579), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n509), .A2(n523), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(KEYINPUT99), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n519), .A2(n525), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n515) );
  NAND2_X1 U580 ( .A1(n519), .A2(n527), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  XOR2_X1 U583 ( .A(G71GAT), .B(KEYINPUT103), .Z(n518) );
  NAND2_X1 U584 ( .A1(n519), .A2(n536), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U587 ( .A1(n519), .A2(n531), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U590 ( .A(KEYINPUT104), .B(n524), .Z(n532) );
  NAND2_X1 U591 ( .A1(n525), .A2(n532), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n532), .A2(n527), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U595 ( .A(G99GAT), .B(KEYINPUT105), .Z(n530) );
  NAND2_X1 U596 ( .A1(n532), .A2(n536), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(KEYINPUT110), .ZN(n553) );
  NOR2_X1 U604 ( .A1(n540), .A2(n553), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n541), .B(KEYINPUT111), .ZN(n550) );
  NOR2_X1 U606 ( .A1(n568), .A2(n550), .ZN(n542) );
  XOR2_X1 U607 ( .A(KEYINPUT112), .B(n542), .Z(n543) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  NOR2_X1 U609 ( .A1(n544), .A2(n550), .ZN(n546) );
  XNOR2_X1 U610 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U612 ( .A(G120GAT), .B(n547), .Z(G1341GAT) );
  NOR2_X1 U613 ( .A1(n571), .A2(n550), .ZN(n548) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(n548), .Z(n549) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  NOR2_X1 U616 ( .A1(n564), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NOR2_X1 U619 ( .A1(n575), .A2(n553), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT114), .B(n554), .Z(n565) );
  NOR2_X1 U621 ( .A1(n568), .A2(n565), .ZN(n555) );
  XOR2_X1 U622 ( .A(G141GAT), .B(n555), .Z(G1344GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n565), .ZN(n560) );
  XOR2_X1 U624 ( .A(KEYINPUT52), .B(KEYINPUT115), .Z(n558) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  XNOR2_X1 U628 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n571), .A2(n565), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(G155GAT), .B(n563), .ZN(G1346GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT118), .B(n566), .Z(n567) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n570), .ZN(n569) );
  XOR2_X1 U636 ( .A(G169GAT), .B(n569), .Z(G1348GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(G183GAT), .B(n572), .Z(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n581) );
  INV_X1 U642 ( .A(n575), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT125), .B(n578), .ZN(n587) );
  AND2_X1 U645 ( .A1(n579), .A2(n587), .ZN(n580) );
  XOR2_X1 U646 ( .A(n581), .B(n580), .Z(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(KEYINPUT62), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

