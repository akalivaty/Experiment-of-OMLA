

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598;

  NOR2_X1 U322 ( .A1(n475), .A2(n579), .ZN(n439) );
  XNOR2_X1 U323 ( .A(n319), .B(n318), .ZN(n320) );
  INV_X1 U324 ( .A(n574), .ZN(n547) );
  XNOR2_X1 U325 ( .A(n380), .B(KEYINPUT111), .ZN(n381) );
  XNOR2_X1 U326 ( .A(n382), .B(n381), .ZN(n402) );
  XOR2_X1 U327 ( .A(G106GAT), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U328 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U329 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U330 ( .A(n373), .B(n372), .ZN(n377) );
  INV_X1 U331 ( .A(KEYINPUT102), .ZN(n482) );
  XNOR2_X1 U332 ( .A(n482), .B(KEYINPUT37), .ZN(n483) );
  XNOR2_X1 U333 ( .A(n587), .B(KEYINPUT41), .ZN(n574) );
  XNOR2_X1 U334 ( .A(n484), .B(n483), .ZN(n526) );
  INV_X1 U335 ( .A(G190GAT), .ZN(n463) );
  INV_X1 U336 ( .A(G183GAT), .ZN(n460) );
  INV_X1 U337 ( .A(n513), .ZN(n537) );
  XOR2_X1 U338 ( .A(KEYINPUT38), .B(n485), .Z(n514) );
  XNOR2_X1 U339 ( .A(n463), .B(KEYINPUT58), .ZN(n464) );
  XNOR2_X1 U340 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U341 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n490), .B(n489), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(G78GAT), .B(G1GAT), .Z(n291) );
  XNOR2_X1 U344 ( .A(G57GAT), .B(G127GAT), .ZN(n290) );
  XNOR2_X1 U345 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U346 ( .A(n292), .B(G211GAT), .Z(n294) );
  XOR2_X1 U347 ( .A(G15GAT), .B(G22GAT), .Z(n340) );
  XNOR2_X1 U348 ( .A(G155GAT), .B(n340), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n299) );
  XNOR2_X1 U350 ( .A(G71GAT), .B(KEYINPUT67), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n295), .B(KEYINPUT13), .ZN(n375) );
  XOR2_X1 U352 ( .A(G183GAT), .B(G8GAT), .Z(n326) );
  XOR2_X1 U353 ( .A(n375), .B(n326), .Z(n297) );
  NAND2_X1 U354 ( .A1(G231GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U356 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U357 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n301) );
  XNOR2_X1 U358 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U360 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n303) );
  XNOR2_X1 U361 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U363 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U364 ( .A(n307), .B(n306), .Z(n566) );
  XOR2_X1 U365 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n309) );
  XNOR2_X1 U366 ( .A(G141GAT), .B(G155GAT), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U368 ( .A(G162GAT), .B(KEYINPUT83), .Z(n310) );
  XOR2_X1 U369 ( .A(n311), .B(n310), .Z(n434) );
  XOR2_X1 U370 ( .A(KEYINPUT23), .B(n363), .Z(n313) );
  XOR2_X1 U371 ( .A(KEYINPUT73), .B(G50GAT), .Z(n387) );
  XNOR2_X1 U372 ( .A(G148GAT), .B(n387), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n319) );
  XOR2_X1 U374 ( .A(KEYINPUT84), .B(KEYINPUT22), .Z(n315) );
  XNOR2_X1 U375 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n314) );
  XOR2_X1 U376 ( .A(n315), .B(n314), .Z(n317) );
  NAND2_X1 U377 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n434), .B(n320), .ZN(n325) );
  XOR2_X1 U379 ( .A(G197GAT), .B(KEYINPUT82), .Z(n322) );
  XNOR2_X1 U380 ( .A(G211GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U382 ( .A(G218GAT), .B(KEYINPUT21), .Z(n323) );
  XOR2_X1 U383 ( .A(n324), .B(n323), .Z(n335) );
  XOR2_X1 U384 ( .A(n325), .B(n335), .Z(n475) );
  XOR2_X1 U385 ( .A(G190GAT), .B(G36GAT), .Z(n388) );
  XNOR2_X1 U386 ( .A(n326), .B(KEYINPUT92), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n327), .B(KEYINPUT91), .ZN(n328) );
  XOR2_X1 U388 ( .A(n388), .B(n328), .Z(n330) );
  NAND2_X1 U389 ( .A1(G226GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n330), .B(n329), .ZN(n332) );
  XNOR2_X1 U391 ( .A(G92GAT), .B(G64GAT), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n331), .B(G176GAT), .ZN(n374) );
  XNOR2_X1 U393 ( .A(n332), .B(n374), .ZN(n337) );
  XOR2_X1 U394 ( .A(G169GAT), .B(KEYINPUT19), .Z(n334) );
  XNOR2_X1 U395 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n333) );
  XNOR2_X1 U396 ( .A(n334), .B(n333), .ZN(n444) );
  XNOR2_X1 U397 ( .A(n444), .B(n335), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n510) );
  INV_X1 U399 ( .A(n510), .ZN(n531) );
  XOR2_X1 U400 ( .A(KEYINPUT29), .B(G197GAT), .Z(n339) );
  XNOR2_X1 U401 ( .A(G141GAT), .B(G8GAT), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U403 ( .A(n341), .B(n340), .Z(n344) );
  XOR2_X1 U404 ( .A(G113GAT), .B(G1GAT), .Z(n416) );
  XNOR2_X1 U405 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n342), .B(KEYINPUT7), .ZN(n392) );
  XNOR2_X1 U407 ( .A(n416), .B(n392), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U409 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n346) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U411 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U412 ( .A(n348), .B(n347), .Z(n353) );
  XOR2_X1 U413 ( .A(G169GAT), .B(G50GAT), .Z(n350) );
  XNOR2_X1 U414 ( .A(G29GAT), .B(G36GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n351), .B(KEYINPUT65), .ZN(n352) );
  XOR2_X1 U417 ( .A(n353), .B(n352), .Z(n582) );
  INV_X1 U418 ( .A(n582), .ZN(n572) );
  XNOR2_X1 U419 ( .A(G120GAT), .B(G148GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n354), .B(G57GAT), .ZN(n425) );
  XNOR2_X1 U421 ( .A(G85GAT), .B(KEYINPUT71), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n355), .B(G99GAT), .ZN(n386) );
  XNOR2_X1 U423 ( .A(n425), .B(n386), .ZN(n379) );
  INV_X1 U424 ( .A(KEYINPUT68), .ZN(n356) );
  NAND2_X1 U425 ( .A1(KEYINPUT70), .A2(n356), .ZN(n359) );
  INV_X1 U426 ( .A(KEYINPUT70), .ZN(n357) );
  NAND2_X1 U427 ( .A1(n357), .A2(KEYINPUT68), .ZN(n358) );
  NAND2_X1 U428 ( .A1(n359), .A2(n358), .ZN(n361) );
  XNOR2_X1 U429 ( .A(G204GAT), .B(KEYINPUT72), .ZN(n360) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n364) );
  INV_X1 U431 ( .A(n364), .ZN(n362) );
  NAND2_X1 U432 ( .A1(n363), .A2(n362), .ZN(n367) );
  INV_X1 U433 ( .A(n363), .ZN(n365) );
  NAND2_X1 U434 ( .A1(n365), .A2(n364), .ZN(n366) );
  NAND2_X1 U435 ( .A1(n367), .A2(n366), .ZN(n373) );
  XOR2_X1 U436 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n369) );
  XNOR2_X1 U437 ( .A(KEYINPUT69), .B(KEYINPUT33), .ZN(n368) );
  XNOR2_X1 U438 ( .A(n369), .B(n368), .ZN(n371) );
  NAND2_X1 U439 ( .A1(G230GAT), .A2(G233GAT), .ZN(n370) );
  XOR2_X1 U440 ( .A(n375), .B(n374), .Z(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n587) );
  NOR2_X1 U443 ( .A1(n572), .A2(n574), .ZN(n382) );
  XNOR2_X1 U444 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n380) );
  XOR2_X1 U445 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n384) );
  XNOR2_X1 U446 ( .A(G162GAT), .B(KEYINPUT74), .ZN(n383) );
  XOR2_X1 U447 ( .A(n384), .B(n383), .Z(n401) );
  XNOR2_X1 U448 ( .A(G29GAT), .B(KEYINPUT75), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n385), .B(G134GAT), .ZN(n426) );
  XNOR2_X1 U450 ( .A(n426), .B(n386), .ZN(n399) );
  XOR2_X1 U451 ( .A(G106GAT), .B(KEYINPUT11), .Z(n390) );
  XNOR2_X1 U452 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U454 ( .A(n391), .B(G92GAT), .Z(n397) );
  XOR2_X1 U455 ( .A(n392), .B(KEYINPUT10), .Z(n394) );
  NAND2_X1 U456 ( .A1(G232GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n395), .B(G218GAT), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n555) );
  INV_X1 U462 ( .A(n555), .ZN(n569) );
  AND2_X1 U463 ( .A1(n402), .A2(n569), .ZN(n403) );
  AND2_X1 U464 ( .A1(n566), .A2(n403), .ZN(n405) );
  XNOR2_X1 U465 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n411) );
  XOR2_X1 U467 ( .A(KEYINPUT36), .B(n555), .Z(n596) );
  NOR2_X1 U468 ( .A1(n596), .A2(n566), .ZN(n406) );
  XNOR2_X1 U469 ( .A(KEYINPUT45), .B(n406), .ZN(n407) );
  NAND2_X1 U470 ( .A1(n407), .A2(n572), .ZN(n408) );
  NOR2_X1 U471 ( .A1(n587), .A2(n408), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n409), .B(KEYINPUT114), .ZN(n410) );
  NOR2_X1 U473 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U474 ( .A(KEYINPUT48), .B(n412), .ZN(n559) );
  NOR2_X1 U475 ( .A1(n531), .A2(n559), .ZN(n415) );
  XOR2_X1 U476 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n413) );
  XNOR2_X1 U477 ( .A(KEYINPUT54), .B(n413), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n435) );
  XOR2_X1 U479 ( .A(KEYINPUT88), .B(G85GAT), .Z(n418) );
  XOR2_X1 U480 ( .A(KEYINPUT0), .B(G127GAT), .Z(n445) );
  XNOR2_X1 U481 ( .A(n445), .B(n416), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n430) );
  XOR2_X1 U483 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n420) );
  XNOR2_X1 U484 ( .A(KEYINPUT6), .B(KEYINPUT86), .ZN(n419) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U486 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n422) );
  XNOR2_X1 U487 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n421) );
  XNOR2_X1 U488 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U489 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U492 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U493 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n473) );
  XOR2_X1 U496 ( .A(KEYINPUT90), .B(n473), .Z(n507) );
  INV_X1 U497 ( .A(n507), .ZN(n528) );
  NAND2_X1 U498 ( .A1(n435), .A2(n528), .ZN(n579) );
  INV_X1 U499 ( .A(n439), .ZN(n437) );
  XNOR2_X1 U500 ( .A(KEYINPUT55), .B(KEYINPUT123), .ZN(n438) );
  INV_X1 U501 ( .A(n438), .ZN(n436) );
  NAND2_X1 U502 ( .A1(n437), .A2(n436), .ZN(n441) );
  NAND2_X1 U503 ( .A1(n439), .A2(n438), .ZN(n440) );
  NAND2_X1 U504 ( .A1(n441), .A2(n440), .ZN(n459) );
  XOR2_X1 U505 ( .A(KEYINPUT81), .B(KEYINPUT64), .Z(n443) );
  XNOR2_X1 U506 ( .A(G134GAT), .B(G190GAT), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n443), .B(n442), .ZN(n458) );
  XOR2_X1 U508 ( .A(n444), .B(G43GAT), .Z(n447) );
  XNOR2_X1 U509 ( .A(n445), .B(G99GAT), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U511 ( .A(G71GAT), .B(KEYINPUT20), .Z(n449) );
  NAND2_X1 U512 ( .A1(G227GAT), .A2(G233GAT), .ZN(n448) );
  XOR2_X1 U513 ( .A(n449), .B(n448), .Z(n450) );
  XNOR2_X1 U514 ( .A(n451), .B(n450), .ZN(n456) );
  XOR2_X1 U515 ( .A(G176GAT), .B(G15GAT), .Z(n453) );
  XNOR2_X1 U516 ( .A(G113GAT), .B(G183GAT), .ZN(n452) );
  XNOR2_X1 U517 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U518 ( .A(G120GAT), .B(n454), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U520 ( .A(n458), .B(n457), .Z(n486) );
  NAND2_X1 U521 ( .A1(n459), .A2(n486), .ZN(n575) );
  NOR2_X1 U522 ( .A1(n566), .A2(n575), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n460), .B(KEYINPUT124), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n462), .B(n461), .ZN(G1350GAT) );
  NOR2_X1 U525 ( .A1(n569), .A2(n575), .ZN(n465) );
  INV_X1 U526 ( .A(n566), .ZN(n591) );
  INV_X1 U527 ( .A(n486), .ZN(n541) );
  NOR2_X1 U528 ( .A1(n531), .A2(n541), .ZN(n466) );
  NOR2_X1 U529 ( .A1(n475), .A2(n466), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n467), .B(KEYINPUT25), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT27), .B(n531), .Z(n476) );
  NAND2_X1 U532 ( .A1(n541), .A2(n475), .ZN(n469) );
  XNOR2_X1 U533 ( .A(KEYINPUT26), .B(KEYINPUT93), .ZN(n468) );
  XNOR2_X1 U534 ( .A(n469), .B(n468), .ZN(n581) );
  NAND2_X1 U535 ( .A1(n476), .A2(n581), .ZN(n470) );
  NAND2_X1 U536 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U537 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n474), .B(KEYINPUT94), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n475), .B(KEYINPUT28), .ZN(n513) );
  NAND2_X1 U540 ( .A1(n476), .A2(n507), .ZN(n560) );
  NOR2_X1 U541 ( .A1(n513), .A2(n560), .ZN(n542) );
  NAND2_X1 U542 ( .A1(n542), .A2(n541), .ZN(n477) );
  NAND2_X1 U543 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U544 ( .A(n479), .B(KEYINPUT95), .ZN(n493) );
  NOR2_X1 U545 ( .A1(n591), .A2(n493), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n480), .B(KEYINPUT101), .ZN(n481) );
  NOR2_X1 U547 ( .A1(n596), .A2(n481), .ZN(n484) );
  NOR2_X1 U548 ( .A1(n572), .A2(n587), .ZN(n494) );
  NAND2_X1 U549 ( .A1(n526), .A2(n494), .ZN(n485) );
  NAND2_X1 U550 ( .A1(n486), .A2(n514), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n488) );
  INV_X1 U552 ( .A(G43GAT), .ZN(n487) );
  NOR2_X1 U553 ( .A1(n555), .A2(n566), .ZN(n491) );
  XOR2_X1 U554 ( .A(KEYINPUT16), .B(n491), .Z(n492) );
  NOR2_X1 U555 ( .A1(n493), .A2(n492), .ZN(n516) );
  NAND2_X1 U556 ( .A1(n494), .A2(n516), .ZN(n504) );
  NOR2_X1 U557 ( .A1(n528), .A2(n504), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U560 ( .A(G1GAT), .B(n497), .Z(G1324GAT) );
  NOR2_X1 U561 ( .A1(n531), .A2(n504), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(G1325GAT) );
  NOR2_X1 U564 ( .A1(n504), .A2(n541), .ZN(n503) );
  XOR2_X1 U565 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n501) );
  XNOR2_X1 U566 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  NOR2_X1 U569 ( .A1(n537), .A2(n504), .ZN(n505) );
  XOR2_X1 U570 ( .A(KEYINPUT100), .B(n505), .Z(n506) );
  XNOR2_X1 U571 ( .A(G22GAT), .B(n506), .ZN(G1327GAT) );
  XOR2_X1 U572 ( .A(G29GAT), .B(KEYINPUT39), .Z(n509) );
  NAND2_X1 U573 ( .A1(n514), .A2(n507), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  XOR2_X1 U575 ( .A(G36GAT), .B(KEYINPUT103), .Z(n512) );
  NAND2_X1 U576 ( .A1(n514), .A2(n510), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1329GAT) );
  NAND2_X1 U578 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U580 ( .A1(n582), .A2(n574), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n527), .A2(n516), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n528), .A2(n523), .ZN(n518) );
  XNOR2_X1 U583 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NOR2_X1 U586 ( .A1(n531), .A2(n523), .ZN(n520) );
  XOR2_X1 U587 ( .A(KEYINPUT106), .B(n520), .Z(n521) );
  XNOR2_X1 U588 ( .A(G64GAT), .B(n521), .ZN(G1333GAT) );
  NOR2_X1 U589 ( .A1(n541), .A2(n523), .ZN(n522) );
  XOR2_X1 U590 ( .A(G71GAT), .B(n522), .Z(G1334GAT) );
  NOR2_X1 U591 ( .A1(n537), .A2(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n536) );
  NOR2_X1 U595 ( .A1(n528), .A2(n536), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(G1336GAT) );
  NOR2_X1 U598 ( .A1(n531), .A2(n536), .ZN(n533) );
  XNOR2_X1 U599 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G92GAT), .B(n534), .ZN(G1337GAT) );
  NOR2_X1 U602 ( .A1(n541), .A2(n536), .ZN(n535) );
  XOR2_X1 U603 ( .A(G99GAT), .B(n535), .Z(G1338GAT) );
  NOR2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n539) );
  XNOR2_X1 U605 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U607 ( .A(G106GAT), .B(n540), .Z(G1339GAT) );
  NOR2_X1 U608 ( .A1(n541), .A2(n559), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n544), .B(KEYINPUT115), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n582), .A2(n556), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(KEYINPUT116), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G113GAT), .B(n546), .ZN(G1340GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U615 ( .A1(n556), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U617 ( .A(G120GAT), .B(n550), .Z(G1341GAT) );
  NAND2_X1 U618 ( .A1(n556), .A2(n591), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(KEYINPUT50), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n554) );
  XNOR2_X1 U622 ( .A(G134GAT), .B(KEYINPUT119), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U625 ( .A(n558), .B(n557), .Z(G1343GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n561), .A2(n581), .ZN(n568) );
  NOR2_X1 U628 ( .A1(n572), .A2(n568), .ZN(n562) );
  XOR2_X1 U629 ( .A(G141GAT), .B(n562), .Z(G1344GAT) );
  NOR2_X1 U630 ( .A1(n574), .A2(n568), .ZN(n564) );
  XNOR2_X1 U631 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(G148GAT), .B(n565), .ZN(G1345GAT) );
  NOR2_X1 U634 ( .A1(n566), .A2(n568), .ZN(n567) );
  XOR2_X1 U635 ( .A(G155GAT), .B(n567), .Z(G1346GAT) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT120), .B(n570), .Z(n571) );
  XNOR2_X1 U638 ( .A(G162GAT), .B(n571), .ZN(G1347GAT) );
  NOR2_X1 U639 ( .A1(n572), .A2(n575), .ZN(n573) );
  XOR2_X1 U640 ( .A(G169GAT), .B(n573), .Z(G1348GAT) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U642 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G176GAT), .B(n578), .ZN(G1349GAT) );
  XOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT60), .Z(n584) );
  INV_X1 U646 ( .A(n579), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n595) );
  INV_X1 U648 ( .A(n595), .ZN(n592) );
  NAND2_X1 U649 ( .A1(n592), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n586) );
  XOR2_X1 U651 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n589) );
  NAND2_X1 U654 ( .A1(n592), .A2(n587), .ZN(n588) );
  XNOR2_X1 U655 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U656 ( .A(G204GAT), .B(n590), .ZN(G1353GAT) );
  XOR2_X1 U657 ( .A(G211GAT), .B(KEYINPUT127), .Z(n594) );
  NAND2_X1 U658 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n594), .B(n593), .ZN(G1354GAT) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U661 ( .A(KEYINPUT62), .B(n597), .Z(n598) );
  XNOR2_X1 U662 ( .A(G218GAT), .B(n598), .ZN(G1355GAT) );
endmodule

