//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n577, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT66), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT70), .ZN(new_n465));
  AND3_X1   g040(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT3), .B1(KEYINPUT69), .B2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT68), .Z(new_n476));
  AOI21_X1  g051(.A(new_n472), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n468), .A2(new_n472), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n469), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(new_n472), .B2(G112), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n480), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT71), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n466), .B2(new_n467), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(KEYINPUT72), .B(new_n487), .C1(new_n466), .C2(new_n467), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT73), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n490), .A2(new_n494), .A3(KEYINPUT4), .A4(new_n491), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n473), .A2(new_n496), .A3(new_n487), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n468), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G2105), .B1(G102), .B2(new_n463), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT74), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT74), .A2(G651), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT6), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(G50), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n506), .A2(new_n507), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G75), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n505), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n508), .A2(G88), .A3(new_n510), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n512), .A2(G62), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n514), .A2(new_n521), .ZN(G166));
  NAND2_X1  g097(.A1(new_n508), .A2(new_n510), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n518), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n523), .A2(new_n505), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n518), .A2(KEYINPUT75), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT5), .B(G543), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n535), .A2(G63), .A3(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n530), .A2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n535), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(new_n512), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n508), .A2(new_n510), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n532), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n541), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n540), .A2(new_n546), .ZN(G171));
  AOI22_X1  g122(.A1(new_n535), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n539), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT76), .ZN(new_n550));
  AOI22_X1  g125(.A1(G43), .A2(new_n526), .B1(new_n524), .B2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT77), .Z(new_n561));
  NAND2_X1  g136(.A1(new_n532), .A2(G65), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n563), .A2(KEYINPUT78), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(KEYINPUT78), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n564), .A2(new_n565), .A3(new_n509), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n543), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n524), .A2(G91), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n526), .A2(KEYINPUT9), .A3(G53), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(new_n514), .ZN(new_n577));
  INV_X1    g152(.A(new_n521), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT79), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n514), .B2(new_n521), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G303));
  NAND4_X1  g157(.A1(new_n508), .A2(G49), .A3(G543), .A4(new_n510), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n508), .A2(G87), .A3(new_n510), .A4(new_n532), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  NAND4_X1  g163(.A1(new_n508), .A2(G48), .A3(G543), .A4(new_n510), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n508), .A2(G86), .A3(new_n510), .A4(new_n532), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n532), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n539), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n518), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n597), .A2(KEYINPUT80), .A3(new_n512), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n591), .A2(new_n594), .A3(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n539), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n602), .A2(new_n543), .B1(new_n544), .B2(new_n603), .ZN(new_n604));
  OR3_X1    g179(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT81), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT81), .B1(new_n601), .B2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n524), .A2(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n518), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n526), .A2(G54), .B1(G651), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n608), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n608), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n573), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n573), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n623), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT82), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(KEYINPUT83), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(KEYINPUT83), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n628), .B(new_n629), .C1(G868), .C2(new_n553), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n479), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n469), .A2(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(new_n472), .B2(G111), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  AND2_X1   g216(.A1(new_n473), .A2(new_n463), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2435), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2438), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2451), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1341), .B(G1348), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n660), .A2(G14), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT87), .ZN(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n663), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT88), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n665), .B(KEYINPUT17), .Z(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(new_n670), .B2(new_n666), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n666), .A3(new_n662), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n665), .A2(new_n667), .A3(new_n662), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(G2100), .Z(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT89), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT19), .Z(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  AOI22_X1  g261(.A1(new_n684), .A2(new_n685), .B1(new_n680), .B2(new_n686), .ZN(new_n687));
  OR3_X1    g262(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(new_n688), .C1(new_n685), .C2(new_n684), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT90), .B(G1986), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G16), .B2(G23), .ZN(new_n700));
  OR3_X1    g275(.A1(new_n699), .A2(G16), .A3(G23), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n700), .B(new_n701), .C1(G288), .C2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT33), .B(G1976), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(KEYINPUT92), .B1(new_n706), .B2(G16), .ZN(new_n707));
  OR3_X1    g282(.A1(new_n706), .A2(KEYINPUT92), .A3(G16), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n707), .B(new_n708), .C1(G166), .C2(new_n702), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G6), .B(G305), .S(G16), .Z(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT32), .B(G1981), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n698), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(KEYINPUT93), .B(KEYINPUT34), .C1(new_n712), .C2(new_n715), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(new_n717), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G24), .B(G290), .S(G16), .Z(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G1986), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n479), .A2(G119), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n469), .A2(G131), .ZN(new_n726));
  NOR2_X1   g301(.A1(G95), .A2(G2105), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(new_n472), .B2(G107), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n725), .B(new_n726), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G25), .B(new_n729), .S(G29), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT35), .B(G1991), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n722), .A2(new_n724), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(KEYINPUT94), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(KEYINPUT94), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n734), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n722), .A2(new_n736), .A3(new_n724), .A4(new_n733), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT26), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n479), .B2(G129), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n463), .A2(G105), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n469), .A2(G141), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G29), .B2(G32), .ZN(new_n749));
  MUX2_X1   g324(.A(new_n748), .B(new_n749), .S(KEYINPUT101), .Z(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n498), .B2(new_n502), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n753), .A2(G27), .ZN(new_n755));
  OAI21_X1  g330(.A(KEYINPUT102), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT102), .B2(new_n755), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2078), .ZN(new_n758));
  NAND2_X1  g333(.A1(G168), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G16), .B2(G21), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n753), .A2(G33), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n473), .A2(G127), .ZN(new_n763));
  INV_X1    g338(.A(G115), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n462), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n765), .A2(G2105), .B1(new_n469), .B2(G139), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT100), .B(KEYINPUT25), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n463), .A2(G103), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n762), .B1(new_n770), .B2(new_n753), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n760), .A2(new_n761), .B1(G2072), .B2(new_n771), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n753), .A2(new_n640), .B1(new_n771), .B2(G2072), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT24), .A2(G34), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n776), .A2(new_n753), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G160), .B2(new_n753), .ZN(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(G28), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(G28), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n783), .A2(new_n784), .A3(new_n753), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n772), .A2(new_n775), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n752), .A2(new_n758), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n702), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n702), .ZN(new_n789));
  INV_X1    g364(.A(G1961), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n787), .B(new_n791), .C1(new_n761), .C2(new_n760), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT103), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n702), .A2(KEYINPUT23), .A3(G20), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT23), .ZN(new_n796));
  INV_X1    g371(.A(G20), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G16), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n795), .B(new_n798), .C1(new_n573), .C2(new_n702), .ZN(new_n799));
  INV_X1    g374(.A(G1956), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  OR3_X1    g376(.A1(KEYINPUT96), .A2(G104), .A3(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G116), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n462), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  OAI21_X1  g379(.A(KEYINPUT96), .B1(G104), .B2(G2105), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n479), .A2(G128), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n469), .A2(G140), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT98), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G29), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT99), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n753), .A2(G26), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT28), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n813), .A2(G2067), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(G2067), .B1(new_n813), .B2(new_n815), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n801), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n792), .B2(new_n793), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n739), .A2(new_n740), .A3(new_n794), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n702), .A2(G19), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n553), .B2(new_n702), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1341), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n702), .A2(G4), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n617), .B2(new_n702), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT95), .B(G1348), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(G29), .A2(G35), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G162), .B2(G29), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT29), .ZN(new_n830));
  INV_X1    g405(.A(G2090), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NOR4_X1   g408(.A1(new_n820), .A2(new_n823), .A3(new_n827), .A4(new_n833), .ZN(G311));
  INV_X1    g409(.A(new_n820), .ZN(new_n835));
  INV_X1    g410(.A(new_n823), .ZN(new_n836));
  INV_X1    g411(.A(new_n827), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n832), .ZN(G150));
  NAND2_X1  g413(.A1(new_n535), .A2(G67), .ZN(new_n839));
  INV_X1    g414(.A(G80), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n505), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n841), .A2(new_n512), .ZN(new_n842));
  INV_X1    g417(.A(G55), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n843), .A2(new_n543), .B1(new_n544), .B2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n550), .A3(new_n551), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n846), .B1(new_n550), .B2(new_n551), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n617), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n849), .B1(new_n857), .B2(G860), .ZN(G145));
  INV_X1    g433(.A(KEYINPUT108), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n770), .A2(KEYINPUT106), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n644), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n811), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n503), .B(new_n729), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n479), .A2(G130), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n469), .A2(G142), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n472), .A2(G118), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT107), .Z(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n865), .B(new_n866), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n746), .B(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n864), .A2(new_n871), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n863), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n875), .A3(new_n862), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n640), .B(G160), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G162), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n859), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  AOI211_X1 g460(.A(KEYINPUT108), .B(new_n885), .C1(new_n878), .C2(new_n880), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n881), .A2(new_n883), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n888), .A2(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g466(.A1(new_n846), .A2(G868), .ZN(new_n892));
  NAND2_X1  g467(.A1(G290), .A2(G288), .ZN(new_n893));
  INV_X1    g468(.A(G288), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n605), .A2(new_n894), .A3(new_n606), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(KEYINPUT109), .A3(new_n895), .ZN(new_n899));
  XOR2_X1   g474(.A(G305), .B(G166), .Z(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n903), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n626), .B(new_n853), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n617), .A2(new_n573), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n616), .B1(new_n572), .B2(new_n566), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n914), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n911), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n910), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n906), .B1(new_n905), .B2(new_n909), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n892), .B1(new_n924), .B2(G868), .ZN(G295));
  AOI21_X1  g500(.A(new_n892), .B1(new_n924), .B2(G868), .ZN(G331));
  OAI21_X1  g501(.A(G286), .B1(KEYINPUT111), .B2(G171), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n842), .A2(new_n845), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n552), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G171), .A2(KEYINPUT111), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n929), .A2(new_n850), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n929), .B2(new_n850), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(KEYINPUT111), .B(G171), .C1(new_n851), .C2(new_n852), .ZN(new_n934));
  INV_X1    g509(.A(new_n927), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n929), .A2(new_n850), .A3(new_n930), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n917), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n933), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n919), .B1(new_n933), .B2(new_n937), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n907), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n931), .A2(new_n932), .A3(new_n927), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n920), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n933), .A2(new_n937), .A3(new_n938), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n904), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G37), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n919), .A2(KEYINPUT112), .A3(KEYINPUT41), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n917), .B2(KEYINPUT112), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n952), .A2(new_n937), .A3(new_n933), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n907), .B1(new_n953), .B2(new_n940), .ZN(new_n954));
  AND4_X1   g529(.A1(KEYINPUT43), .A2(new_n954), .A3(new_n947), .A4(new_n946), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n954), .A2(new_n949), .A3(new_n947), .A4(new_n946), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n961), .ZN(G397));
  XNOR2_X1  g537(.A(KEYINPUT113), .B(G1384), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n503), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G40), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n471), .A2(new_n968), .A3(new_n477), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(G1996), .A3(new_n746), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(KEYINPUT114), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n972), .A2(KEYINPUT114), .ZN(new_n974));
  INV_X1    g549(.A(G2067), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n811), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G1996), .B2(new_n746), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n973), .B(new_n974), .C1(new_n971), .C2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n971), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n729), .B(new_n732), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(G290), .B(G1986), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n971), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n503), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n498), .B2(new_n502), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n986), .A2(new_n780), .A3(new_n969), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT118), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n969), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n761), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n970), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n780), .A4(new_n989), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n991), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G8), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G168), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT124), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(G8), .B(new_n1005), .C1(new_n999), .C2(G286), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n999), .A2(G8), .A3(G286), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G305), .A2(G1981), .ZN(new_n1012));
  INV_X1    g587(.A(G1981), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n591), .A2(new_n1013), .A3(new_n594), .A4(new_n598), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT49), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n503), .A2(new_n984), .A3(new_n969), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(KEYINPUT49), .A3(new_n1014), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(G8), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(G288), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G288), .A2(new_n1021), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1018), .A2(new_n1022), .A3(G8), .A4(new_n1024), .ZN(new_n1025));
  AOI211_X1 g600(.A(new_n1001), .B(new_n1023), .C1(new_n987), .C2(new_n969), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1020), .B(new_n1025), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1018), .A2(G8), .A3(new_n1024), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT52), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(KEYINPUT117), .A3(new_n1020), .A4(new_n1025), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n966), .B(new_n963), .C1(new_n498), .C2(new_n502), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n710), .B1(new_n994), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n986), .A2(new_n831), .A3(new_n969), .A4(new_n989), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(G303), .B2(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1039), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n1001), .B(new_n1041), .C1(new_n579), .C2(new_n581), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(KEYINPUT116), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1038), .A2(G8), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1001), .B(new_n1047), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1034), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n970), .B1(new_n985), .B2(new_n966), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(G2078), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n992), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n969), .B1(new_n987), .B2(new_n988), .ZN(new_n1055));
  AOI211_X1 g630(.A(KEYINPUT50), .B(G1384), .C1(new_n498), .C2(new_n502), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n790), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n994), .A2(G2078), .A3(new_n1035), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1054), .B(new_n1057), .C1(new_n1058), .C2(KEYINPUT53), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G171), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT62), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1007), .A2(new_n1062), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1011), .A2(new_n1050), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n999), .A2(G8), .A3(G168), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n999), .A2(KEYINPUT119), .A3(G8), .A4(G168), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1038), .A2(G8), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1028), .B1(new_n1070), .B2(new_n1043), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1043), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1069), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1049), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(KEYINPUT63), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1018), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1020), .A2(new_n1021), .A3(new_n894), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1001), .B(new_n1078), .C1(new_n1079), .C2(new_n1014), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1028), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1072), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1064), .A2(new_n1077), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n476), .A2(new_n474), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1084), .A2(KEYINPUT125), .ZN(new_n1085));
  OAI21_X1  g660(.A(G2105), .B1(new_n1084), .B2(KEYINPUT125), .ZN(new_n1086));
  OAI21_X1  g661(.A(G40), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n963), .B1(new_n498), .B2(new_n502), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(KEYINPUT45), .ZN(new_n1089));
  INV_X1    g664(.A(new_n471), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n967), .A2(new_n1089), .A3(new_n1090), .A4(new_n1053), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1057), .B(new_n1091), .C1(new_n1058), .C2(KEYINPUT53), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G171), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1088), .A2(KEYINPUT45), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(new_n969), .C1(KEYINPUT45), .C2(new_n987), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1052), .B1(new_n1095), .B2(G2078), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1096), .A2(G301), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1093), .A2(KEYINPUT54), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n1049), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1096), .A2(G301), .A3(new_n1057), .A4(new_n1091), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT54), .B1(new_n1060), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(KEYINPUT126), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT126), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n1103), .B(KEYINPUT54), .C1(new_n1060), .C2(new_n1100), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1099), .B(new_n1010), .C1(new_n1102), .C2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT56), .B(G2072), .Z(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1095), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n800), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1107), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1051), .A2(KEYINPUT121), .A3(new_n1094), .A4(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n569), .A2(KEYINPUT120), .A3(new_n571), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(new_n573), .B(new_n1115), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1348), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1078), .A2(new_n975), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1117), .B1(new_n616), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1116), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(new_n1108), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT61), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1119), .A2(new_n616), .A3(new_n1120), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n616), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT60), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1121), .A2(new_n1130), .A3(new_n617), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1126), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1117), .A2(KEYINPUT61), .A3(new_n1124), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1117), .A2(KEYINPUT123), .A3(KEYINPUT61), .A4(new_n1124), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT58), .B(G1341), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1018), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT122), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1095), .A2(G1996), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n553), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT59), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1133), .A2(new_n1136), .A3(new_n1137), .A4(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1105), .B1(new_n1125), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n983), .B1(new_n1083), .B2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n979), .A2(G290), .A3(G1986), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1148));
  XNOR2_X1  g723(.A(new_n1147), .B(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n981), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n729), .A2(new_n731), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n978), .A2(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n811), .A2(G2067), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n979), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n979), .B1(new_n976), .B2(new_n747), .ZN(new_n1155));
  OR3_X1    g730(.A1(new_n979), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT46), .B1(new_n979), .B2(G1996), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT47), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1150), .A2(new_n1154), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1146), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g736(.A1(G401), .A2(G227), .ZN(new_n1163));
  AOI21_X1  g737(.A(new_n1163), .B1(new_n887), .B2(new_n889), .ZN(new_n1164));
  AND4_X1   g738(.A1(G319), .A2(new_n1164), .A3(new_n959), .A4(new_n696), .ZN(G308));
  NAND4_X1  g739(.A1(new_n1164), .A2(new_n959), .A3(G319), .A4(new_n696), .ZN(G225));
endmodule


