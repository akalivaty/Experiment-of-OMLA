

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593;

  XOR2_X2 U326 ( .A(KEYINPUT38), .B(n493), .Z(n504) );
  XOR2_X1 U327 ( .A(n439), .B(n438), .Z(n520) );
  XNOR2_X1 U328 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U329 ( .A(n413), .B(KEYINPUT111), .ZN(n414) );
  XOR2_X1 U330 ( .A(n435), .B(KEYINPUT97), .Z(n294) );
  XOR2_X1 U331 ( .A(G92GAT), .B(G218GAT), .Z(n295) );
  XOR2_X1 U332 ( .A(KEYINPUT25), .B(n467), .Z(n296) );
  INV_X1 U333 ( .A(KEYINPUT46), .ZN(n413) );
  XNOR2_X1 U334 ( .A(n371), .B(KEYINPUT75), .ZN(n372) );
  XNOR2_X1 U335 ( .A(n373), .B(n372), .ZN(n374) );
  NOR2_X1 U336 ( .A1(n591), .A2(n489), .ZN(n490) );
  NOR2_X1 U337 ( .A1(n545), .A2(n442), .ZN(n575) );
  XNOR2_X1 U338 ( .A(n443), .B(KEYINPUT55), .ZN(n570) );
  XNOR2_X1 U339 ( .A(n461), .B(KEYINPUT122), .ZN(n462) );
  XNOR2_X1 U340 ( .A(n463), .B(n462), .ZN(G1350GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n298) );
  XNOR2_X1 U342 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U344 ( .A(G197GAT), .B(n299), .Z(n431) );
  XOR2_X1 U345 ( .A(G50GAT), .B(G162GAT), .Z(n364) );
  XNOR2_X1 U346 ( .A(G78GAT), .B(KEYINPUT73), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n300), .B(G148GAT), .ZN(n385) );
  XOR2_X1 U348 ( .A(n364), .B(n385), .Z(n302) );
  NAND2_X1 U349 ( .A1(G228GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n431), .B(n303), .ZN(n315) );
  XOR2_X1 U352 ( .A(G204GAT), .B(KEYINPUT24), .Z(n305) );
  XNOR2_X1 U353 ( .A(KEYINPUT23), .B(KEYINPUT93), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U355 ( .A(n306), .B(G106GAT), .Z(n308) );
  XOR2_X1 U356 ( .A(G22GAT), .B(G155GAT), .Z(n346) );
  XNOR2_X1 U357 ( .A(n346), .B(G218GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U359 ( .A(n309), .B(KEYINPUT22), .Z(n313) );
  XOR2_X1 U360 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n311) );
  XNOR2_X1 U361 ( .A(G141GAT), .B(KEYINPUT92), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n330) );
  XNOR2_X1 U363 ( .A(n330), .B(KEYINPUT89), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n470) );
  XOR2_X1 U366 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n317) );
  XNOR2_X1 U367 ( .A(KEYINPUT4), .B(KEYINPUT94), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n336) );
  XOR2_X1 U369 ( .A(KEYINPUT5), .B(G57GAT), .Z(n319) );
  XNOR2_X1 U370 ( .A(G1GAT), .B(G127GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U372 ( .A(KEYINPUT77), .B(G155GAT), .Z(n321) );
  XNOR2_X1 U373 ( .A(G120GAT), .B(G148GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n334) );
  XOR2_X1 U376 ( .A(G113GAT), .B(KEYINPUT0), .Z(n448) );
  XOR2_X1 U377 ( .A(G85GAT), .B(G162GAT), .Z(n325) );
  XNOR2_X1 U378 ( .A(G29GAT), .B(G134GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U380 ( .A(n448), .B(n326), .Z(n328) );
  NAND2_X1 U381 ( .A1(G225GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U383 ( .A(n329), .B(KEYINPUT95), .Z(n332) );
  XNOR2_X1 U384 ( .A(n330), .B(KEYINPUT96), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U387 ( .A(n336), .B(n335), .Z(n518) );
  INV_X1 U388 ( .A(n518), .ZN(n545) );
  XOR2_X1 U389 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n338) );
  XNOR2_X1 U390 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n354) );
  XOR2_X1 U392 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n340) );
  NAND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U395 ( .A(n341), .B(KEYINPUT82), .Z(n345) );
  XNOR2_X1 U396 ( .A(G8GAT), .B(G1GAT), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n342), .B(KEYINPUT67), .ZN(n397) );
  XNOR2_X1 U398 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n343), .B(KEYINPUT13), .ZN(n384) );
  XNOR2_X1 U400 ( .A(n397), .B(n384), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n350) );
  XOR2_X1 U402 ( .A(n346), .B(G78GAT), .Z(n348) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G127GAT), .Z(n454) );
  XNOR2_X1 U404 ( .A(n454), .B(G211GAT), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U406 ( .A(n350), .B(n349), .Z(n352) );
  XNOR2_X1 U407 ( .A(G183GAT), .B(G71GAT), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n552) );
  XOR2_X1 U410 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n356) );
  XNOR2_X1 U411 ( .A(KEYINPUT76), .B(KEYINPUT9), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n370) );
  XOR2_X1 U413 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n358) );
  NAND2_X1 U414 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n360) );
  XNOR2_X1 U416 ( .A(G36GAT), .B(G190GAT), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n295), .B(n359), .ZN(n432) );
  XOR2_X1 U418 ( .A(n360), .B(n432), .Z(n363) );
  XNOR2_X1 U419 ( .A(G99GAT), .B(G106GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n361), .B(G85GAT), .ZN(n373) );
  XNOR2_X1 U421 ( .A(KEYINPUT77), .B(n373), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U423 ( .A(n365), .B(n364), .Z(n368) );
  XNOR2_X1 U424 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n366), .B(KEYINPUT8), .ZN(n408) );
  XOR2_X1 U426 ( .A(G43GAT), .B(G134GAT), .Z(n446) );
  XNOR2_X1 U427 ( .A(n408), .B(n446), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n555) );
  NAND2_X1 U430 ( .A1(n552), .A2(n555), .ZN(n417) );
  AND2_X1 U431 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U432 ( .A(G176GAT), .B(n374), .ZN(n378) );
  XOR2_X1 U433 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n376) );
  XNOR2_X1 U434 ( .A(KEYINPUT32), .B(KEYINPUT71), .ZN(n375) );
  XOR2_X1 U435 ( .A(n376), .B(n375), .Z(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n383) );
  XOR2_X1 U437 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n380) );
  XOR2_X1 U438 ( .A(G120GAT), .B(G71GAT), .Z(n449) );
  XOR2_X1 U439 ( .A(G204GAT), .B(G64GAT), .Z(n436) );
  XNOR2_X1 U440 ( .A(n449), .B(n436), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U442 ( .A(n381), .B(G92GAT), .Z(n382) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n582) );
  XNOR2_X1 U446 ( .A(n582), .B(KEYINPUT41), .ZN(n561) );
  XOR2_X1 U447 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n389) );
  XNOR2_X1 U448 ( .A(KEYINPUT64), .B(KEYINPUT66), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n412) );
  XOR2_X1 U450 ( .A(G197GAT), .B(G22GAT), .Z(n391) );
  XNOR2_X1 U451 ( .A(G43GAT), .B(G141GAT), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U453 ( .A(KEYINPUT69), .B(G15GAT), .Z(n393) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(G113GAT), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U456 ( .A(n395), .B(n394), .Z(n405) );
  INV_X1 U457 ( .A(G50GAT), .ZN(n396) );
  NAND2_X1 U458 ( .A1(n396), .A2(n397), .ZN(n400) );
  INV_X1 U459 ( .A(n397), .ZN(n398) );
  NAND2_X1 U460 ( .A1(G50GAT), .A2(n398), .ZN(n399) );
  NAND2_X1 U461 ( .A1(n400), .A2(n399), .ZN(n402) );
  NAND2_X1 U462 ( .A1(G229GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n403), .B(G36GAT), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n407) );
  INV_X1 U466 ( .A(KEYINPUT29), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n408), .B(KEYINPUT68), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n506) );
  INV_X1 U471 ( .A(n506), .ZN(n576) );
  NOR2_X1 U472 ( .A1(n561), .A2(n576), .ZN(n415) );
  OR2_X1 U473 ( .A1(n417), .A2(n416), .ZN(n418) );
  XNOR2_X1 U474 ( .A(KEYINPUT47), .B(n418), .ZN(n424) );
  XNOR2_X1 U475 ( .A(KEYINPUT80), .B(n555), .ZN(n568) );
  XNOR2_X1 U476 ( .A(KEYINPUT36), .B(n568), .ZN(n591) );
  NOR2_X1 U477 ( .A1(n591), .A2(n552), .ZN(n420) );
  XNOR2_X1 U478 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  NAND2_X1 U480 ( .A1(n421), .A2(n576), .ZN(n422) );
  NOR2_X1 U481 ( .A1(n582), .A2(n422), .ZN(n423) );
  NOR2_X1 U482 ( .A1(n424), .A2(n423), .ZN(n425) );
  XNOR2_X1 U483 ( .A(KEYINPUT48), .B(n425), .ZN(n544) );
  XOR2_X1 U484 ( .A(KEYINPUT86), .B(KEYINPUT18), .Z(n427) );
  XNOR2_X1 U485 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U487 ( .A(n428), .B(G183GAT), .Z(n430) );
  XNOR2_X1 U488 ( .A(G169GAT), .B(G176GAT), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n459) );
  XNOR2_X1 U490 ( .A(n459), .B(n431), .ZN(n439) );
  XOR2_X1 U491 ( .A(n432), .B(KEYINPUT98), .Z(n434) );
  NAND2_X1 U492 ( .A1(G226GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U494 ( .A(G8GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n294), .B(n437), .ZN(n438) );
  XNOR2_X1 U496 ( .A(KEYINPUT118), .B(n520), .ZN(n440) );
  NOR2_X1 U497 ( .A1(n544), .A2(n440), .ZN(n441) );
  XOR2_X1 U498 ( .A(KEYINPUT54), .B(n441), .Z(n442) );
  NAND2_X1 U499 ( .A1(n470), .A2(n575), .ZN(n443) );
  XOR2_X1 U500 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n445) );
  XNOR2_X1 U501 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n453) );
  XOR2_X1 U504 ( .A(n449), .B(n448), .Z(n451) );
  NAND2_X1 U505 ( .A1(G227GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n455) );
  XOR2_X1 U508 ( .A(n455), .B(n454), .Z(n457) );
  XNOR2_X1 U509 ( .A(G190GAT), .B(G99GAT), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X2 U511 ( .A(n459), .B(n458), .Z(n567) );
  NOR2_X1 U512 ( .A1(n552), .A2(n567), .ZN(n460) );
  AND2_X1 U513 ( .A1(n570), .A2(n460), .ZN(n463) );
  INV_X1 U514 ( .A(G183GAT), .ZN(n461) );
  INV_X1 U515 ( .A(n552), .ZN(n586) );
  NAND2_X1 U516 ( .A1(n568), .A2(n586), .ZN(n464) );
  XOR2_X1 U517 ( .A(KEYINPUT16), .B(n464), .Z(n477) );
  INV_X1 U518 ( .A(n520), .ZN(n497) );
  INV_X1 U519 ( .A(n567), .ZN(n557) );
  NAND2_X1 U520 ( .A1(n497), .A2(n557), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n465), .A2(n470), .ZN(n466) );
  XNOR2_X1 U522 ( .A(n466), .B(KEYINPUT100), .ZN(n467) );
  NOR2_X1 U523 ( .A1(n557), .A2(n470), .ZN(n468) );
  XNOR2_X1 U524 ( .A(n468), .B(KEYINPUT26), .ZN(n574) );
  XOR2_X1 U525 ( .A(n520), .B(KEYINPUT27), .Z(n471) );
  NAND2_X1 U526 ( .A1(n574), .A2(n471), .ZN(n543) );
  NAND2_X1 U527 ( .A1(n296), .A2(n543), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n469), .A2(n518), .ZN(n476) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT28), .ZN(n526) );
  AND2_X1 U530 ( .A1(n471), .A2(n526), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n472), .A2(n545), .ZN(n529) );
  XOR2_X1 U532 ( .A(KEYINPUT88), .B(n567), .Z(n473) );
  NOR2_X1 U533 ( .A1(n529), .A2(n473), .ZN(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT99), .B(n474), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n488) );
  NAND2_X1 U536 ( .A1(n477), .A2(n488), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT101), .B(n478), .ZN(n507) );
  NOR2_X1 U538 ( .A1(n576), .A2(n582), .ZN(n492) );
  NAND2_X1 U539 ( .A1(n507), .A2(n492), .ZN(n479) );
  XOR2_X1 U540 ( .A(KEYINPUT102), .B(n479), .Z(n485) );
  NAND2_X1 U541 ( .A1(n545), .A2(n485), .ZN(n480) );
  XNOR2_X1 U542 ( .A(KEYINPUT34), .B(n480), .ZN(n481) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NAND2_X1 U544 ( .A1(n485), .A2(n497), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n482), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U547 ( .A1(n485), .A2(n557), .ZN(n483) );
  XNOR2_X1 U548 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  XOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT103), .Z(n487) );
  INV_X1 U550 ( .A(n526), .ZN(n503) );
  NAND2_X1 U551 ( .A1(n503), .A2(n485), .ZN(n486) );
  XNOR2_X1 U552 ( .A(n487), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n495) );
  NAND2_X1 U554 ( .A1(n552), .A2(n488), .ZN(n489) );
  XOR2_X1 U555 ( .A(KEYINPUT104), .B(n490), .Z(n491) );
  XNOR2_X1 U556 ( .A(KEYINPUT37), .B(n491), .ZN(n516) );
  NAND2_X1 U557 ( .A1(n516), .A2(n492), .ZN(n493) );
  NAND2_X1 U558 ( .A1(n504), .A2(n545), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U560 ( .A(G29GAT), .B(n496), .Z(G1328GAT) );
  NAND2_X1 U561 ( .A1(n504), .A2(n497), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n498), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n502) );
  XOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n500) );
  NAND2_X1 U565 ( .A1(n504), .A2(n557), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U570 ( .A1(n506), .A2(n561), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n507), .A2(n517), .ZN(n512) );
  NOR2_X1 U572 ( .A1(n518), .A2(n512), .ZN(n508) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n508), .Z(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n520), .A2(n512), .ZN(n510) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n567), .A2(n512), .ZN(n511) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n511), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n526), .A2(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n525) );
  NOR2_X1 U584 ( .A1(n518), .A2(n525), .ZN(n519) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n519), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n520), .A2(n525), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1337GAT) );
  NOR2_X1 U589 ( .A1(n567), .A2(n525), .ZN(n523) );
  XOR2_X1 U590 ( .A(KEYINPUT110), .B(n523), .Z(n524) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n524), .ZN(G1338GAT) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n527), .Z(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n544), .A2(n529), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n530), .A2(n557), .ZN(n538) );
  NOR2_X1 U597 ( .A1(n576), .A2(n538), .ZN(n531) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n531), .Z(G1340GAT) );
  NOR2_X1 U599 ( .A1(n561), .A2(n538), .ZN(n533) );
  XNOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  NOR2_X1 U603 ( .A1(n552), .A2(n538), .ZN(n536) );
  XNOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n537), .Z(G1342GAT) );
  NOR2_X1 U607 ( .A1(n538), .A2(n568), .ZN(n542) );
  XOR2_X1 U608 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n540) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n539) );
  XNOR2_X1 U610 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n546) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n554) );
  NOR2_X1 U614 ( .A1(n576), .A2(n554), .ZN(n547) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  NOR2_X1 U616 ( .A1(n554), .A2(n561), .ZN(n551) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n548) );
  XNOR2_X1 U619 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n552), .A2(n554), .ZN(n553) );
  XOR2_X1 U622 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n556), .Z(G1347GAT) );
  XNOR2_X1 U625 ( .A(KEYINPUT119), .B(G169GAT), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n570), .A2(n557), .ZN(n560) );
  NOR2_X1 U627 ( .A1(n560), .A2(n576), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  NOR2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n566) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n563) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n562) );
  XNOR2_X1 U632 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(n564), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n590) );
  NOR2_X1 U641 ( .A1(n576), .A2(n590), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(KEYINPUT124), .B(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n584) );
  INV_X1 U648 ( .A(n590), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(n585), .ZN(G1353GAT) );
  XOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT127), .Z(n589) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

