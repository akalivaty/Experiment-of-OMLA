//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  OAI21_X1  g0007(.A(G50), .B1(G58), .B2(G68), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n217), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G68), .ZN(new_n244));
  INV_X1    g0044(.A(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n243), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(new_n211), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(new_n220), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT23), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(new_n211), .B2(G107), .ZN(new_n254));
  INV_X1    g0054(.A(G107), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(KEYINPUT23), .A3(G20), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT22), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n258), .B1(new_n262), .B2(G87), .ZN(new_n263));
  INV_X1    g0063(.A(G87), .ZN(new_n264));
  NOR4_X1   g0064(.A1(new_n261), .A2(KEYINPUT22), .A3(G20), .A4(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n257), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT24), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT69), .B1(new_n269), .B2(new_n210), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n210), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n266), .B2(new_n267), .ZN(new_n274));
  INV_X1    g0074(.A(new_n272), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(new_n270), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  INV_X1    g0077(.A(G1), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT68), .A2(G1), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n279), .A2(G13), .A3(G20), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G33), .A3(new_n280), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n276), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G107), .ZN(new_n285));
  OR3_X1    g0085(.A1(new_n281), .A2(KEYINPUT25), .A3(G107), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT25), .B1(new_n281), .B2(G107), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n285), .A2(KEYINPUT85), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n281), .B(new_n282), .C1(new_n275), .C2(new_n270), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n286), .B(new_n287), .C1(new_n289), .C2(new_n255), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT85), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n268), .A2(new_n274), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n279), .A2(G45), .A3(new_n280), .ZN(new_n294));
  AND2_X1   g0094(.A1(KEYINPUT5), .A2(G41), .ZN(new_n295));
  NOR2_X1   g0095(.A1(KEYINPUT5), .A2(G41), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT67), .ZN(new_n299));
  AND2_X1   g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n210), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G41), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n302), .A2(KEYINPUT67), .A3(G1), .A4(G13), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n298), .A2(G274), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(G257), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n305));
  INV_X1    g0105(.A(G1698), .ZN(new_n306));
  OAI211_X1 g0106(.A(G250), .B(new_n306), .C1(new_n259), .C2(new_n260), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G294), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n300), .A2(new_n210), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT68), .A2(G1), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT68), .A2(G1), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT5), .B(G41), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(G45), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n316), .A2(G264), .A3(new_n301), .A4(new_n303), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n304), .A2(new_n311), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT86), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT86), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n304), .A2(new_n311), .A3(new_n317), .A4(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(G169), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n293), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G200), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT87), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT87), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n318), .A2(new_n329), .A3(new_n326), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(G190), .B1(new_n319), .B2(new_n321), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n293), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT88), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT88), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n293), .B(new_n335), .C1(new_n331), .C2(new_n332), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n325), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n281), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n202), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n314), .A2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n273), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT8), .B(G58), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G20), .A2(G33), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n342), .A2(new_n251), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(G20), .B2(new_n203), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n339), .B1(new_n341), .B2(new_n202), .C1(new_n347), .C2(new_n273), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT9), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT3), .ZN(new_n351));
  INV_X1    g0151(.A(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(KEYINPUT3), .A2(G33), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n306), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(G223), .B1(new_n261), .B2(G77), .ZN(new_n356));
  INV_X1    g0156(.A(G222), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n306), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n356), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n310), .ZN(new_n361));
  INV_X1    g0161(.A(G41), .ZN(new_n362));
  INV_X1    g0162(.A(G45), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n279), .A2(new_n364), .A3(new_n280), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(new_n301), .A3(new_n303), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n366), .A2(new_n219), .ZN(new_n367));
  AOI21_X1  g0167(.A(G1), .B1(new_n362), .B2(new_n363), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n301), .A2(G274), .A3(new_n303), .A4(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n361), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G200), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n348), .A2(new_n349), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n350), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n361), .A2(G190), .A3(new_n367), .A4(new_n369), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT73), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT74), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT10), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(KEYINPUT10), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n377), .A2(KEYINPUT10), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n379), .B(new_n380), .C1(new_n373), .C2(new_n375), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n370), .A2(G179), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n370), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n348), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n344), .A2(G50), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT76), .ZN(new_n388));
  INV_X1    g0188(.A(G77), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n251), .A2(new_n389), .B1(new_n211), .B2(G68), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n276), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n391), .B(KEYINPUT11), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n273), .A2(G68), .A3(new_n340), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT77), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n338), .A2(new_n245), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT12), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n392), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  XOR2_X1   g0198(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n310), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n261), .A2(G1698), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n358), .A2(G232), .A3(G1698), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G238), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n369), .B1(new_n366), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n400), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n404), .B(new_n409), .C1(new_n359), .C2(new_n219), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n310), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n366), .A2(new_n406), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n369), .A3(new_n399), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(G169), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n405), .A2(new_n407), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  OAI211_X1 g0218(.A(G179), .B(new_n413), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n415), .B1(new_n414), .B2(G169), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n398), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(G200), .ZN(new_n423));
  OAI211_X1 g0223(.A(G190), .B(new_n413), .C1(new_n417), .C2(new_n418), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n397), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g0227(.A(KEYINPUT8), .B(G58), .Z(new_n428));
  INV_X1    g0228(.A(KEYINPUT72), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(new_n344), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n429), .B2(new_n344), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n432), .A2(new_n251), .B1(new_n211), .B2(new_n389), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n276), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n273), .A2(G77), .A3(new_n340), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n338), .A2(new_n389), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n365), .A2(new_n301), .A3(G244), .A4(new_n303), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n369), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT70), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n355), .A2(G238), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n358), .A2(G232), .A3(new_n306), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n261), .A2(G107), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n310), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT70), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n438), .A2(new_n369), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT71), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n440), .A2(new_n445), .A3(KEYINPUT71), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n437), .B1(new_n452), .B2(new_n323), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n383), .A3(new_n451), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n439), .A2(KEYINPUT70), .B1(new_n444), .B2(new_n310), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT71), .B1(new_n456), .B2(new_n447), .ZN(new_n457));
  INV_X1    g0257(.A(new_n451), .ZN(new_n458));
  OAI21_X1  g0258(.A(G190), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n450), .A2(G200), .A3(new_n451), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n437), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT17), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n352), .A2(new_n264), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n355), .B2(G226), .ZN(new_n465));
  OAI211_X1 g0265(.A(G223), .B(new_n306), .C1(new_n259), .C2(new_n260), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n401), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n365), .A2(new_n301), .A3(G232), .A4(new_n303), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n369), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  NOR4_X1   g0270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .A4(G190), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n326), .B1(new_n467), .B2(new_n469), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT80), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n468), .A2(new_n369), .ZN(new_n474));
  INV_X1    g0274(.A(G190), .ZN(new_n475));
  OAI211_X1 g0275(.A(G226), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n476));
  INV_X1    g0276(.A(new_n464), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n466), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n310), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n471), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n341), .A2(new_n428), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n281), .A2(new_n342), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n353), .A2(new_n211), .A3(new_n354), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT7), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n353), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n354), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(KEYINPUT79), .A3(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n490), .A2(KEYINPUT79), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(G68), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G58), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n245), .ZN(new_n495));
  OAI21_X1  g0295(.A(G20), .B1(new_n495), .B2(new_n201), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n344), .A2(G159), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n486), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT7), .B1(new_n261), .B2(new_n211), .ZN(new_n501));
  INV_X1    g0301(.A(new_n490), .ZN(new_n502));
  OAI21_X1  g0302(.A(G68), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(KEYINPUT16), .A3(new_n499), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n276), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n484), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n463), .B1(new_n481), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n482), .A2(new_n483), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n493), .A2(new_n499), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n485), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n489), .A2(new_n490), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n498), .B1(new_n511), .B2(G68), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n273), .B1(new_n512), .B2(KEYINPUT16), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n508), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n479), .A2(new_n369), .A3(new_n468), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G169), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n474), .A2(G179), .A3(new_n479), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT18), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n474), .A2(KEYINPUT80), .A3(new_n475), .A4(new_n479), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n470), .B1(new_n515), .B2(new_n326), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n515), .A2(G190), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n514), .A2(new_n523), .A3(KEYINPUT17), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT18), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n516), .A2(new_n517), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n506), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n507), .A2(new_n519), .A3(new_n524), .A4(new_n527), .ZN(new_n528));
  NOR4_X1   g0328(.A1(new_n386), .A2(new_n427), .A3(new_n462), .A4(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT21), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT83), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n301), .B(new_n303), .C1(new_n294), .C2(new_n297), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n301), .A2(G274), .A3(new_n303), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n532), .A2(new_n221), .B1(new_n533), .B2(new_n316), .ZN(new_n534));
  OAI211_X1 g0334(.A(G264), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n535));
  OAI211_X1 g0335(.A(G257), .B(new_n306), .C1(new_n259), .C2(new_n260), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n353), .A2(G303), .A3(new_n354), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n538), .A2(new_n310), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n531), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n310), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n316), .A2(G270), .A3(new_n301), .A4(new_n303), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n304), .A2(new_n541), .A3(new_n542), .A4(KEYINPUT83), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n281), .A2(G116), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G283), .ZN(new_n547));
  INV_X1    g0347(.A(G97), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n211), .C1(G33), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n269), .A2(new_n210), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n220), .A2(G20), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT20), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT20), .A4(new_n551), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n546), .B(new_n556), .C1(new_n220), .C2(new_n289), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G169), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n530), .B1(new_n544), .B2(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n534), .A2(new_n539), .A3(new_n323), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n557), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n545), .B1(new_n284), .B2(G116), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n383), .B1(new_n562), .B2(new_n556), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(KEYINPUT21), .A3(new_n540), .A4(new_n543), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n557), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n567), .C1(new_n544), .C2(new_n326), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n544), .A2(G190), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n566), .B1(new_n544), .B2(new_n326), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT84), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n565), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n491), .A2(G107), .A3(new_n492), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n255), .A2(KEYINPUT6), .A3(G97), .ZN(new_n575));
  XOR2_X1   g0375(.A(G97), .B(G107), .Z(new_n576));
  OAI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(KEYINPUT6), .ZN(new_n577));
  OR3_X1    g0377(.A1(new_n345), .A2(KEYINPUT81), .A3(new_n389), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT81), .B1(new_n345), .B2(new_n389), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n577), .A2(G20), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n276), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n281), .A2(G97), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n289), .B2(new_n548), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(KEYINPUT82), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT82), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n273), .B1(new_n574), .B2(new_n580), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(new_n585), .ZN(new_n590));
  OAI211_X1 g0390(.A(G244), .B(new_n306), .C1(new_n259), .C2(new_n260), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT4), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n358), .A2(KEYINPUT4), .A3(G244), .A4(new_n306), .ZN(new_n594));
  OAI211_X1 g0394(.A(G250), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n547), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n310), .ZN(new_n597));
  INV_X1    g0397(.A(G257), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n532), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n304), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G169), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n597), .A2(G179), .A3(new_n304), .A4(new_n599), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n587), .A2(new_n590), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n589), .A2(new_n585), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(G200), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n532), .A2(new_n598), .B1(new_n533), .B2(new_n316), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n310), .B2(new_n596), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G190), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n358), .A2(new_n211), .A3(G68), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT19), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n211), .B1(new_n409), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(G87), .B2(new_n206), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n251), .B2(new_n548), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n276), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n273), .A2(G87), .A3(new_n281), .A4(new_n282), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n338), .A2(new_n432), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(G238), .B(new_n306), .C1(new_n259), .C2(new_n260), .ZN(new_n621));
  OAI211_X1 g0421(.A(G244), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n622));
  NAND2_X1  g0422(.A1(G33), .A2(G116), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n310), .ZN(new_n625));
  INV_X1    g0425(.A(G250), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n294), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G274), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n279), .A2(G45), .A3(new_n628), .A4(new_n280), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n627), .A2(new_n301), .A3(new_n303), .A4(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n326), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n625), .A2(new_n630), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n620), .B(new_n632), .C1(new_n475), .C2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n616), .B(new_n618), .C1(new_n289), .C2(new_n432), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n383), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n635), .B(new_n636), .C1(G179), .C2(new_n633), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n603), .A2(new_n609), .A3(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n337), .A2(new_n529), .A3(new_n573), .A4(new_n639), .ZN(G372));
  NAND2_X1  g0440(.A1(new_n632), .A2(KEYINPUT89), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n625), .A2(G190), .A3(new_n630), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT89), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n631), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n641), .A2(new_n642), .A3(new_n620), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n637), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n647));
  INV_X1    g0447(.A(new_n293), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n322), .A2(new_n324), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n646), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n334), .A2(new_n336), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n603), .A2(new_n609), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT90), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n601), .A2(new_n602), .ZN(new_n656));
  INV_X1    g0456(.A(new_n604), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n645), .A2(new_n656), .A3(new_n637), .A4(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n637), .B1(new_n658), .B2(KEYINPUT26), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n634), .A2(new_n637), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n603), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n655), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT82), .B1(new_n582), .B2(new_n586), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n589), .A2(new_n588), .A3(new_n585), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n656), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT26), .B1(new_n666), .B2(new_n638), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n604), .B1(new_n601), .B2(new_n602), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(new_n660), .A3(new_n637), .A4(new_n645), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n667), .A2(KEYINPUT90), .A3(new_n637), .A4(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n654), .A2(new_n663), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n529), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n385), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n519), .A2(new_n527), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n422), .A2(new_n455), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n426), .A2(new_n507), .A3(new_n524), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n378), .A2(new_n381), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(G369));
  AND2_X1   g0480(.A1(new_n211), .A2(G13), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n314), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n566), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n572), .A2(new_n569), .A3(new_n568), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n647), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT91), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n692), .B2(new_n691), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n647), .A2(new_n689), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G330), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n337), .B1(new_n293), .B2(new_n688), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n325), .A2(new_n687), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n650), .A2(new_n687), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n647), .A2(new_n687), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n337), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n215), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n209), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n709), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n337), .A2(new_n573), .A3(new_n639), .A4(new_n688), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n540), .A2(new_n543), .ZN(new_n717));
  AOI21_X1  g0517(.A(G179), .B1(new_n625), .B2(new_n630), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n318), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n607), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n720), .A3(KEYINPUT92), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n591), .A2(new_n592), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n595), .A2(new_n547), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n401), .B1(new_n725), .B2(new_n593), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n318), .B(new_n718), .C1(new_n726), .C2(new_n606), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n722), .B1(new_n544), .B2(new_n727), .ZN(new_n728));
  AND4_X1   g0528(.A1(new_n317), .A2(new_n311), .A3(new_n625), .A4(new_n630), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n560), .A2(new_n607), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n560), .A2(new_n607), .A3(new_n729), .A4(KEYINPUT30), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n721), .A2(new_n728), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n734), .B2(new_n687), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n687), .A2(KEYINPUT31), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n732), .A2(new_n733), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n717), .A2(new_n720), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n715), .B1(new_n716), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n671), .A2(new_n688), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT93), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n671), .A2(KEYINPUT93), .A3(new_n688), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT94), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n603), .B2(new_n609), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n666), .A2(KEYINPUT94), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n651), .A2(new_n652), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n658), .A2(KEYINPUT26), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n661), .A2(new_n603), .A3(new_n660), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n753), .A2(new_n754), .A3(new_n637), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n687), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT29), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n741), .B1(new_n747), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n714), .B1(new_n758), .B2(G1), .ZN(G364));
  AOI21_X1  g0559(.A(new_n278), .B1(new_n681), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n708), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n707), .A2(new_n261), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n764), .A2(G355), .B1(new_n220), .B2(new_n707), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n707), .A2(new_n358), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n712), .B2(G45), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n249), .A2(new_n363), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n210), .B1(G20), .B2(new_n383), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n763), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n773), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n211), .A2(new_n326), .A3(G179), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n475), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT97), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT97), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G107), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(G20), .A3(new_n323), .ZN(new_n785));
  INV_X1    g0585(.A(G159), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT32), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OR3_X1    g0587(.A1(new_n785), .A2(KEYINPUT32), .A3(new_n786), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n211), .A2(new_n323), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n475), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G50), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n783), .A2(new_n787), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n777), .A2(G190), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n358), .B1(new_n794), .B2(new_n264), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n790), .A2(G190), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n475), .A2(G200), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n211), .B1(new_n798), .B2(new_n323), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n797), .A2(new_n245), .B1(new_n548), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT96), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n789), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n798), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n784), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n494), .A2(new_n803), .B1(new_n804), .B2(new_n389), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n793), .A2(new_n795), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n785), .B(KEYINPUT98), .Z(new_n807));
  AOI22_X1  g0607(.A1(new_n782), .A2(G283), .B1(new_n807), .B2(G329), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT99), .ZN(new_n809));
  NOR2_X1   g0609(.A1(KEYINPUT33), .A2(G317), .ZN(new_n810));
  AND2_X1   g0610(.A1(KEYINPUT33), .A2(G317), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n796), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n791), .A2(G326), .ZN(new_n813));
  INV_X1    g0613(.A(G294), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n799), .ZN(new_n815));
  INV_X1    g0615(.A(G303), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n261), .B1(new_n816), .B2(new_n794), .C1(new_n804), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n803), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n815), .B(new_n818), .C1(G322), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n806), .B1(new_n809), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n694), .A2(new_n695), .ZN(new_n822));
  INV_X1    g0622(.A(new_n772), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n775), .B1(new_n776), .B2(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(G330), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT95), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n696), .A2(new_n763), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(G396));
  INV_X1    g0628(.A(G283), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n804), .A2(new_n220), .B1(new_n829), .B2(new_n797), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT100), .Z(new_n831));
  INV_X1    g0631(.A(new_n807), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n832), .A2(new_n817), .B1(new_n803), .B2(new_n814), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n261), .B1(new_n799), .B2(new_n548), .ZN(new_n834));
  INV_X1    g0634(.A(new_n791), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n835), .A2(new_n816), .B1(new_n255), .B2(new_n794), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n831), .B(new_n837), .C1(new_n264), .C2(new_n781), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G137), .A2(new_n791), .B1(new_n796), .B2(G150), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT101), .ZN(new_n840));
  INV_X1    g0640(.A(G143), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n841), .B2(new_n803), .C1(new_n786), .C2(new_n804), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT34), .Z(new_n843));
  OAI221_X1 g0643(.A(new_n358), .B1(new_n799), .B2(new_n494), .C1(new_n794), .C2(new_n202), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G132), .B2(new_n807), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n245), .B2(new_n781), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n838), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n773), .A2(new_n770), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n847), .A2(new_n773), .B1(new_n389), .B2(new_n848), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n437), .A2(new_n688), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n461), .A2(new_n850), .B1(new_n453), .B2(new_n454), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n453), .A2(new_n454), .A3(new_n688), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT102), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n460), .A2(new_n437), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n475), .B1(new_n450), .B2(new_n451), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n850), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n455), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT102), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n852), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n849), .B1(new_n861), .B2(new_n771), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n762), .ZN(new_n863));
  INV_X1    g0663(.A(new_n861), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n744), .A2(new_n746), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n741), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n671), .A2(new_n861), .A3(new_n688), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n763), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n863), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT103), .ZN(G384));
  XNOR2_X1  g0672(.A(new_n577), .B(KEYINPUT104), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT35), .ZN(new_n874));
  OAI211_X1 g0674(.A(G116), .B(new_n212), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n874), .B2(new_n873), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT36), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n209), .B(G77), .C1(new_n494), .C2(new_n245), .ZN(new_n878));
  AOI211_X1 g0678(.A(G13), .B(new_n314), .C1(new_n878), .C2(new_n244), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT40), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n514), .A2(new_n685), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n528), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n514), .A2(new_n523), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n506), .A2(new_n526), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT106), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n885), .A2(KEYINPUT106), .A3(new_n886), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n685), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT37), .B1(new_n506), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n885), .A3(new_n886), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT107), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT107), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n893), .A2(new_n885), .A3(new_n896), .A4(new_n886), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n883), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n504), .B(new_n276), .C1(new_n512), .C2(new_n486), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n685), .B1(new_n902), .B2(new_n484), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n528), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n512), .A2(new_n486), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n505), .A2(new_n905), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n906), .A2(new_n508), .B1(new_n526), .B2(new_n892), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n884), .B1(new_n885), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT105), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n894), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI211_X1 g0710(.A(KEYINPUT105), .B(new_n884), .C1(new_n885), .C2(new_n907), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n904), .B(KEYINPUT38), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n881), .B1(new_n901), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n398), .A2(new_n687), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n422), .A2(new_n426), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n414), .A2(G169), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT14), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n419), .A3(new_n416), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n398), .B(new_n687), .C1(new_n918), .C2(new_n425), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n854), .A2(new_n860), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n735), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n716), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n481), .A2(new_n506), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n518), .A2(new_n685), .B1(new_n484), .B2(new_n902), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT37), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT105), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n908), .A2(new_n909), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n929), .A3(new_n894), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n930), .B2(new_n904), .ZN(new_n931));
  INV_X1    g0731(.A(new_n912), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n923), .B(new_n920), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n913), .A2(new_n924), .B1(new_n933), .B2(new_n881), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n934), .A2(new_n529), .A3(new_n923), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n529), .B2(new_n923), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n935), .A2(new_n936), .A3(new_n715), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n747), .A2(new_n529), .A3(new_n757), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n679), .ZN(new_n939));
  XOR2_X1   g0739(.A(KEYINPUT108), .B(KEYINPUT39), .Z(new_n940));
  AND2_X1   g0740(.A1(new_n528), .A2(new_n882), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n514), .A2(new_n518), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n888), .B1(new_n925), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n882), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n944), .A3(new_n890), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT37), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n895), .A2(new_n897), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n941), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n912), .B(new_n940), .C1(new_n948), .C2(KEYINPUT38), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT39), .B1(new_n931), .B2(new_n932), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n422), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n688), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n915), .A2(new_n919), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n867), .B2(new_n852), .ZN(new_n958));
  INV_X1    g0758(.A(new_n931), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n912), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n674), .A2(new_n892), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n955), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n939), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n937), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n314), .B2(new_n681), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n937), .A2(new_n965), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n880), .B1(new_n967), .B2(new_n968), .ZN(G367));
  INV_X1    g0769(.A(new_n766), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n774), .B1(new_n215), .B2(new_n432), .C1(new_n238), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n762), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n797), .A2(new_n786), .B1(new_n245), .B2(new_n799), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G143), .B2(new_n791), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n782), .A2(G77), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n819), .A2(G150), .ZN(new_n976));
  INV_X1    g0776(.A(G137), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n358), .B1(new_n977), .B2(new_n785), .C1(new_n794), .C2(new_n494), .ZN(new_n978));
  INV_X1    g0778(.A(new_n804), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(new_n979), .B2(G50), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n781), .A2(new_n548), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(G283), .ZN(new_n984));
  INV_X1    g0784(.A(new_n794), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(G116), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT46), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n261), .B1(new_n988), .B2(new_n785), .C1(new_n799), .C2(new_n255), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G294), .B2(new_n796), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n983), .A2(new_n984), .A3(new_n987), .A4(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n803), .A2(new_n816), .B1(new_n817), .B2(new_n835), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT113), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n981), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT47), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n972), .B1(new_n995), .B2(new_n773), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n688), .A2(new_n620), .ZN(new_n997));
  MUX2_X1   g0797(.A(new_n646), .B(new_n637), .S(new_n997), .Z(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n772), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT110), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n652), .A2(new_n704), .A3(new_n650), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n703), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n657), .A2(new_n687), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n749), .A2(new_n751), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n668), .A2(new_n687), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1002), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n705), .A2(new_n1011), .A3(KEYINPUT110), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1001), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n705), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1005), .A2(new_n1009), .A3(new_n1002), .ZN(new_n1018));
  OAI21_X1  g0818(.A(KEYINPUT110), .B1(new_n705), .B2(new_n1011), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n1019), .A3(KEYINPUT44), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n702), .A2(new_n1013), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1003), .B1(new_n699), .B2(new_n704), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(new_n696), .Z(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1023), .A3(new_n758), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1020), .A2(new_n1017), .ZN(new_n1026));
  AOI21_X1  g0826(.A(KEYINPUT44), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT111), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT111), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1013), .A2(new_n1029), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1030));
  AND4_X1   g0830(.A1(KEYINPUT112), .A2(new_n1028), .A3(new_n701), .A4(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1013), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n702), .B1(new_n1032), .B2(KEYINPUT111), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT112), .B1(new_n1033), .B2(new_n1030), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1025), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n758), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n708), .B(KEYINPUT41), .Z(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n761), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1011), .A2(new_n337), .A3(new_n704), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT42), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT43), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n666), .B1(new_n1009), .B2(new_n650), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n688), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n998), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT109), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n998), .B(KEYINPUT43), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n702), .A2(new_n1009), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1048), .A2(new_n1053), .A3(new_n1051), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1000), .B1(new_n1039), .B2(new_n1057), .ZN(G387));
  INV_X1    g0858(.A(new_n774), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n764), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1060), .A2(new_n710), .B1(G107), .B2(new_n215), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n235), .A2(new_n363), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n710), .ZN(new_n1063));
  AOI211_X1 g0863(.A(G45), .B(new_n1063), .C1(G68), .C2(G77), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n342), .A2(G50), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n970), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1061), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n358), .B1(new_n785), .B2(new_n343), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n791), .B2(G159), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n804), .B2(new_n245), .C1(new_n202), .C2(new_n803), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n799), .A2(new_n432), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n985), .A2(G77), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n797), .B2(new_n342), .ZN(new_n1075));
  NOR4_X1   g0875(.A1(new_n1072), .A2(new_n982), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G311), .A2(new_n796), .B1(new_n791), .B2(G322), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n804), .B2(new_n816), .C1(new_n988), .C2(new_n803), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT48), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n799), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n985), .A2(G294), .B1(new_n1082), .B2(G283), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT49), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n785), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n358), .B1(new_n1087), .B2(G326), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n781), .B2(new_n220), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT115), .Z(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1076), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n762), .B1(new_n1059), .B2(new_n1069), .C1(new_n1092), .C2(new_n776), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n700), .B2(new_n772), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1023), .B2(new_n761), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1023), .A2(new_n758), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n708), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1023), .A2(new_n758), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(G393));
  OAI221_X1 g0899(.A(new_n774), .B1(new_n548), .B2(new_n215), .C1(new_n242), .C2(new_n970), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n762), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n803), .A2(new_n786), .B1(new_n343), .B2(new_n835), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n794), .A2(new_n245), .B1(new_n841), .B2(new_n785), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G87), .C2(new_n782), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n979), .A2(new_n428), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n799), .A2(new_n389), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n261), .B(new_n1109), .C1(G50), .C2(new_n796), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1103), .A2(new_n1107), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n358), .B1(new_n1087), .B2(G322), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n783), .B(new_n1112), .C1(new_n829), .C2(new_n794), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT117), .Z(new_n1114));
  OAI22_X1  g0914(.A1(new_n803), .A2(new_n817), .B1(new_n988), .B2(new_n835), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT52), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n796), .A2(G303), .B1(new_n1082), .B2(G116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n814), .C2(new_n804), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1111), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1101), .B1(new_n1119), .B2(new_n773), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1011), .B2(new_n823), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1032), .A2(new_n701), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1021), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1028), .A2(new_n701), .A3(new_n1030), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT112), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1033), .A2(KEYINPUT112), .A3(new_n1030), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1024), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1123), .A2(new_n1096), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n708), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1121), .B1(new_n760), .B2(new_n1123), .C1(new_n1128), .C2(new_n1130), .ZN(G390));
  OAI21_X1  g0931(.A(new_n912), .B1(new_n948), .B2(KEYINPUT38), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n853), .B1(new_n756), .B2(new_n861), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n953), .B(new_n1132), .C1(new_n1133), .C2(new_n957), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n741), .A2(new_n956), .A3(new_n861), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n867), .A2(new_n852), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n954), .B1(new_n1136), .B2(new_n956), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1134), .B(new_n1135), .C1(new_n1137), .C2(new_n951), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n920), .A2(new_n923), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(new_n715), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n950), .B(new_n949), .C1(new_n958), .C2(new_n954), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n1134), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n956), .B1(new_n741), .B2(new_n861), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1136), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n923), .A2(G330), .A3(new_n861), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1133), .B(new_n1135), .C1(new_n1148), .C2(new_n956), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n529), .A2(G330), .A3(new_n923), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n938), .A2(new_n1152), .A3(new_n679), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1145), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1153), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1150), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1134), .B1(new_n1137), .B2(new_n951), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1141), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1138), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1155), .A2(new_n1161), .A3(new_n708), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1145), .A2(new_n761), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n848), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n762), .B1(new_n428), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n797), .A2(new_n255), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1109), .B(new_n1166), .C1(G283), .C2(new_n791), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n261), .B1(new_n794), .B2(new_n264), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT118), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(new_n245), .C2(new_n781), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n819), .A2(G116), .B1(G294), .B2(new_n807), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n548), .B2(new_n804), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n819), .A2(G132), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n985), .A2(G150), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT54), .B(G143), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1173), .B1(KEYINPUT53), .B2(new_n1174), .C1(new_n804), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n782), .A2(G50), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n261), .B1(new_n796), .B2(G137), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n791), .A2(G128), .B1(new_n1082), .B2(G159), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n807), .A2(G125), .B1(new_n1174), .B2(KEYINPUT53), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1170), .A2(new_n1172), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1165), .B1(new_n1182), .B2(new_n773), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT119), .Z(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n951), .B2(new_n771), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1162), .A2(new_n1163), .A3(new_n1185), .ZN(G378));
  INV_X1    g0986(.A(KEYINPUT122), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n358), .A2(G41), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n245), .B2(new_n799), .C1(new_n804), .C2(new_n432), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n832), .A2(new_n829), .B1(new_n803), .B2(new_n255), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1074), .B1(new_n797), .B2(new_n548), .C1(new_n220), .C2(new_n835), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n781), .A2(new_n494), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT120), .Z(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(G33), .A2(G41), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1188), .A2(G50), .A3(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G128), .A2(new_n819), .B1(new_n979), .B2(G137), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n791), .A2(G125), .B1(new_n1082), .B2(G150), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1175), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n985), .A2(new_n1202), .B1(new_n796), .B2(G132), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1087), .A2(G124), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1198), .B(new_n1206), .C1(new_n781), .C2(new_n786), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1204), .B2(KEYINPUT59), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1199), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1196), .A2(new_n1197), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n773), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n763), .B1(new_n202), .B2(new_n848), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n386), .A2(new_n348), .A3(new_n892), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n348), .A2(new_n892), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n378), .A2(new_n381), .A3(new_n385), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1213), .A2(new_n1215), .A3(new_n1217), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1211), .B(new_n1212), .C1(new_n1221), .C2(new_n771), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n934), .B2(G330), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n924), .A2(new_n1132), .A3(KEYINPUT40), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n931), .A2(new_n932), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n881), .B1(new_n1225), .B2(new_n1140), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1224), .A2(new_n1226), .A3(new_n1221), .A4(G330), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1136), .A2(new_n960), .A3(new_n956), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n953), .B1(new_n949), .B2(new_n950), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n962), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1223), .A2(new_n1228), .B1(new_n1231), .B2(KEYINPUT121), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1224), .A2(new_n1226), .A3(G330), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1221), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT121), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1235), .A2(new_n964), .A3(new_n1236), .A4(new_n1227), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1222), .B1(new_n1238), .B2(new_n760), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT57), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1153), .B1(new_n1145), .B2(new_n1154), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(new_n1241), .B2(new_n1238), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n964), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1231), .A2(new_n1235), .A3(new_n1227), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1240), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1156), .B1(new_n1160), .B2(new_n1151), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n709), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1187), .B(new_n1239), .C1(new_n1242), .C2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1242), .A2(new_n1247), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1239), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT122), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1248), .A2(new_n1251), .ZN(G375));
  OAI21_X1  g1052(.A(new_n762), .B1(G68), .B2(new_n1164), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n358), .B(new_n1073), .C1(new_n819), .C2(G283), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n255), .B2(new_n804), .C1(new_n816), .C2(new_n832), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G97), .A2(new_n985), .B1(new_n796), .B2(G116), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n975), .B(new_n1256), .C1(new_n814), .C2(new_n835), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G132), .A2(new_n791), .B1(new_n796), .B2(new_n1202), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n803), .B2(new_n977), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT123), .Z(new_n1260));
  AND2_X1   g1060(.A1(new_n807), .A2(G128), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n804), .A2(new_n343), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n358), .B1(new_n799), .B2(new_n202), .C1(new_n794), .C2(new_n786), .ZN(new_n1263));
  OR4_X1    g1063(.A1(new_n1192), .A2(new_n1261), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1255), .A2(new_n1257), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1253), .B1(new_n1265), .B2(new_n773), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n956), .B2(new_n771), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1151), .B2(new_n760), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1154), .A2(new_n1037), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(G381));
  INV_X1    g1072(.A(G384), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1271), .A3(new_n1274), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(G387), .A2(G390), .A3(G378), .A4(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1251), .B2(new_n1248), .ZN(G407));
  INV_X1    g1077(.A(new_n1244), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1231), .B1(new_n1227), .B2(new_n1235), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT57), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n708), .B1(new_n1280), .B2(new_n1241), .ZN(new_n1281));
  AND4_X1   g1081(.A1(new_n1236), .A2(new_n1235), .A3(new_n964), .A4(new_n1227), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1235), .A2(new_n1227), .B1(new_n964), .B2(new_n1236), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT57), .B1(new_n1284), .B2(new_n1246), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1250), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1187), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1239), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT122), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G378), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n686), .A2(G213), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(G407), .A2(G213), .A3(new_n1293), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1294), .B(KEYINPUT124), .ZN(G409));
  INV_X1    g1095(.A(G390), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n758), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1038), .B1(new_n1128), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1057), .B1(new_n1298), .B2(new_n760), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1000), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1296), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1000), .B(G390), .C1(new_n1039), .C2(new_n1057), .ZN(new_n1302));
  XOR2_X1   g1102(.A(G393), .B(G396), .Z(new_n1303));
  AND3_X1   g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1305));
  OR2_X1    g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(KEYINPUT61), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1284), .A2(new_n1038), .A3(new_n1246), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1308), .B(new_n1222), .C1(new_n760), .C2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(G378), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1288), .A2(G378), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(KEYINPUT125), .B1(new_n1314), .B2(new_n1292), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1151), .A2(new_n1153), .A3(KEYINPUT60), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n708), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1157), .A2(KEYINPUT60), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1318), .B2(new_n1270), .ZN(new_n1319));
  OR3_X1    g1119(.A1(new_n1319), .A2(G384), .A3(new_n1268), .ZN(new_n1320));
  OAI21_X1  g1120(.A(G384), .B1(new_n1319), .B2(new_n1268), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(G2897), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1322), .B1(new_n1323), .B2(new_n1291), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1320), .A2(G2897), .A3(new_n1292), .A4(new_n1321), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT125), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n1328), .A3(new_n1291), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1315), .A2(new_n1326), .A3(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1327), .A2(new_n1291), .A3(new_n1322), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  OR2_X1    g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1307), .A2(new_n1330), .A3(new_n1333), .A4(new_n1334), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1324), .B(new_n1325), .C1(new_n1314), .C2(new_n1292), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1331), .A2(KEYINPUT62), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1327), .A2(new_n1339), .A3(new_n1291), .A4(new_n1322), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1336), .A2(new_n1337), .A3(new_n1338), .A4(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1306), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1335), .A2(new_n1342), .ZN(G405));
  AND2_X1   g1143(.A1(new_n1322), .A2(KEYINPUT126), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1288), .A2(new_n1311), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1344), .B1(new_n1290), .B2(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1311), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1322), .A2(KEYINPUT126), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1345), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1348), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1346), .A2(new_n1347), .A3(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT127), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1346), .A2(new_n1351), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1306), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1346), .A2(new_n1347), .A3(new_n1351), .A4(KEYINPUT127), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1354), .A2(new_n1356), .A3(new_n1357), .ZN(G402));
endmodule


