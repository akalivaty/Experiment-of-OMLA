//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  OR2_X1    g002(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT81), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n206));
  NAND4_X1  g005(.A1(new_n204), .A2(new_n205), .A3(G148gat), .A4(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(new_n211), .B2(KEYINPUT2), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT80), .A2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(G148gat), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT81), .B1(new_n217), .B2(G148gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n207), .B(new_n212), .C1(new_n216), .C2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G141gat), .B(G148gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n208), .B(new_n211), .C1(new_n220), .C2(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223));
  INV_X1    g022(.A(G218gat), .ZN(new_n224));
  OR2_X1    g023(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT76), .B(KEYINPUT22), .Z(new_n228));
  OAI21_X1  g027(.A(new_n223), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G211gat), .B(G218gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n230), .B(new_n223), .C1(new_n227), .C2(new_n228), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT29), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n222), .B1(new_n234), .B2(KEYINPUT3), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n236));
  INV_X1    g035(.A(new_n233), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n238));
  AND2_X1   g037(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(KEYINPUT77), .A2(G211gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n238), .B1(new_n241), .B2(new_n224), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n230), .B1(new_n242), .B2(new_n223), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n236), .B1(new_n237), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n219), .A2(new_n245), .A3(new_n221), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n232), .A2(KEYINPUT78), .A3(new_n233), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G228gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G22gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT87), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n247), .B1(new_n243), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n232), .A2(KEYINPUT87), .A3(new_n233), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT3), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n222), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n251), .B(new_n253), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT86), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n256), .B1(new_n255), .B2(new_n262), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT88), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G78gat), .B(G106gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n255), .A2(new_n262), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G22gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT88), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n264), .A3(new_n272), .A4(new_n263), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n267), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n269), .B1(new_n267), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n203), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n251), .A2(new_n253), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n258), .A2(new_n259), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n222), .B1(new_n278), .B2(KEYINPUT3), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n277), .A2(new_n279), .B1(new_n252), .B2(new_n254), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT86), .B1(new_n280), .B2(new_n256), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n272), .B1(new_n281), .B2(new_n271), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n265), .A2(KEYINPUT88), .A3(new_n266), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n268), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n267), .A2(new_n269), .A3(new_n273), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n202), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(KEYINPUT24), .A3(new_n293), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n293), .A2(KEYINPUT24), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n291), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT25), .B1(new_n298), .B2(KEYINPUT66), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n299), .B1(KEYINPUT66), .B2(new_n298), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n291), .A2(new_n297), .A3(new_n294), .A4(new_n295), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n302));
  AOI22_X1  g101(.A1(new_n296), .A2(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G183gat), .ZN(new_n304));
  AOI21_X1  g103(.A(G190gat), .B1(new_n304), .B2(KEYINPUT27), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n305), .B(KEYINPUT28), .C1(KEYINPUT27), .C2(new_n304), .ZN(new_n306));
  AND2_X1   g105(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n308));
  OAI21_X1  g107(.A(G183gat), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT68), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n311), .B(G183gat), .C1(new_n307), .C2(new_n308), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n310), .A2(KEYINPUT69), .A3(new_n305), .A4(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n305), .ZN(new_n316));
  OR2_X1    g115(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n304), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(new_n319), .B2(new_n311), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT69), .B1(new_n320), .B2(new_n310), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n306), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n323), .A2(KEYINPUT71), .ZN(new_n324));
  AOI211_X1 g123(.A(G169gat), .B(G176gat), .C1(new_n323), .C2(KEYINPUT71), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n297), .B1(new_n289), .B2(new_n323), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n324), .A2(new_n325), .B1(new_n326), .B2(KEYINPUT70), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(KEYINPUT70), .B2(new_n326), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n328), .A2(new_n293), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n303), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n288), .B1(new_n330), .B2(KEYINPUT29), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n293), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n333));
  INV_X1    g132(.A(new_n310), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n312), .A2(new_n305), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(new_n314), .A3(new_n313), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n332), .B1(new_n337), .B2(new_n306), .ZN(new_n338));
  OAI211_X1 g137(.A(G226gat), .B(G233gat), .C1(new_n338), .C2(new_n303), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n244), .A2(new_n250), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n331), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n288), .B1(new_n330), .B2(new_n247), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n342), .B2(new_n339), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  AOI21_X1  g146(.A(KEYINPUT30), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n347), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n341), .B2(new_n343), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n339), .A3(new_n340), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n322), .A2(new_n329), .ZN(new_n354));
  INV_X1    g153(.A(new_n303), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n288), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n248), .B1(new_n338), .B2(new_n303), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(new_n288), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n351), .B(new_n353), .C1(new_n358), .C2(new_n340), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT89), .B1(new_n348), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n339), .ZN(new_n362));
  INV_X1    g161(.A(new_n340), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n347), .A3(new_n351), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n352), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n350), .A4(new_n359), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G134gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G127gat), .ZN(new_n372));
  INV_X1    g171(.A(G127gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G134gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT1), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT72), .ZN(new_n377));
  INV_X1    g176(.A(G120gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(G113gat), .ZN(new_n379));
  INV_X1    g178(.A(G113gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n379), .B(new_n381), .C1(new_n380), .C2(G120gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT1), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n380), .A2(G120gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n378), .A2(G113gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n376), .A2(new_n382), .B1(new_n386), .B2(new_n375), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n338), .B2(new_n303), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n376), .A2(new_n382), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n375), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n330), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n393), .B(KEYINPUT64), .Z(new_n394));
  NAND3_X1  g193(.A1(new_n388), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT32), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(G15gat), .B(G43gat), .Z(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G71gat), .B(G99gat), .Z(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n396), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n403), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n395), .B(KEYINPUT32), .C1(new_n397), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n392), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n393), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT34), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n394), .A2(KEYINPUT34), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n407), .A2(new_n413), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n287), .A2(new_n370), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT0), .ZN(new_n421));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT4), .B1(new_n222), .B2(new_n391), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n387), .A2(new_n427), .A3(new_n219), .A4(new_n221), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n222), .A2(KEYINPUT3), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n391), .A3(new_n246), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n387), .A2(new_n219), .A3(new_n221), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n429), .A2(new_n430), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n222), .A2(new_n391), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n433), .ZN(new_n437));
  INV_X1    g236(.A(new_n430), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT83), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n440), .B(new_n430), .C1(new_n436), .C2(new_n433), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n435), .B(KEYINPUT5), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n425), .A2(KEYINPUT84), .A3(new_n428), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n261), .A2(new_n444), .A3(new_n427), .A4(new_n387), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT5), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n447), .A3(new_n430), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n419), .B(new_n424), .C1(new_n442), .C2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n423), .B1(new_n446), .B2(new_n449), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n442), .A2(new_n452), .A3(KEYINPUT85), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT85), .B1(new_n442), .B2(new_n452), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT5), .B1(new_n439), .B2(new_n441), .ZN(new_n456));
  AND4_X1   g255(.A1(new_n430), .A2(new_n429), .A3(new_n432), .A4(new_n434), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n450), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT6), .B1(new_n458), .B2(new_n423), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n451), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(KEYINPUT92), .B(KEYINPUT35), .Z(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n460), .A2(new_n348), .A3(new_n360), .ZN(new_n465));
  INV_X1    g264(.A(new_n416), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(new_n414), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n465), .A2(new_n467), .A3(new_n286), .A4(new_n276), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n418), .A2(new_n464), .B1(KEYINPUT35), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT90), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n456), .A2(new_n457), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n443), .A2(new_n445), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n424), .B1(new_n473), .B2(new_n448), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n423), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n442), .A2(new_n452), .A3(KEYINPUT85), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n419), .A4(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n451), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n365), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n349), .A2(KEYINPUT37), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n351), .B1(new_n358), .B2(new_n340), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n482), .B2(new_n349), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT38), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n331), .A2(new_n339), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT37), .B1(new_n485), .B2(new_n340), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n363), .B1(new_n342), .B2(new_n339), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n470), .B1(new_n480), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n362), .A2(new_n340), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n491), .B(KEYINPUT37), .C1(new_n340), .C2(new_n485), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n347), .B1(new_n364), .B2(new_n351), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n492), .B(new_n484), .C1(new_n493), .C2(new_n481), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n460), .A2(KEYINPUT90), .A3(new_n494), .A4(new_n365), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n482), .A2(KEYINPUT37), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT38), .B1(new_n496), .B2(new_n483), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n490), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n274), .A2(new_n275), .A3(new_n203), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n202), .B1(new_n284), .B2(new_n285), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n443), .A2(new_n445), .A3(new_n432), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n438), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n436), .A2(new_n433), .A3(new_n430), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(KEYINPUT39), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n424), .B1(new_n504), .B2(KEYINPUT39), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n504), .A2(KEYINPUT39), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n510), .A2(KEYINPUT40), .A3(new_n424), .A4(new_n506), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n509), .A2(new_n511), .A3(new_n476), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n361), .A2(new_n368), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n501), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT91), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n513), .A2(new_n286), .A3(new_n276), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n498), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  OR3_X1    g318(.A1(new_n460), .A2(new_n348), .A3(new_n360), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n287), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n415), .A2(new_n416), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n467), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n469), .B1(new_n519), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT100), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OR3_X1    g332(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n535), .B2(new_n534), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT95), .B(G36gat), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G29gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G43gat), .B(G50gat), .Z(new_n541));
  INV_X1    g340(.A(KEYINPUT15), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT96), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n534), .B2(new_n532), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n542), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n539), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT16), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(new_n553), .B2(G1gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(G1gat), .B2(new_n552), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G8gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n545), .A2(KEYINPUT17), .A3(new_n548), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n551), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n549), .A2(new_n556), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G113gat), .B(G141gat), .Z(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT93), .B(G197gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT11), .B(G169gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT12), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT98), .B1(new_n549), .B2(new_n556), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n545), .A2(new_n574), .A3(new_n548), .A4(new_n557), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n575), .A3(new_n561), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n560), .B(KEYINPUT13), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n559), .A2(KEYINPUT18), .A3(new_n560), .A4(new_n561), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT99), .B1(new_n572), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n578), .A2(new_n579), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n571), .A4(new_n564), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n564), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n562), .A2(KEYINPUT97), .A3(new_n563), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(new_n582), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n570), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n531), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n585), .A2(new_n531), .A3(new_n590), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n530), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G99gat), .B(G106gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  NAND3_X1  g403(.A1(new_n551), .A2(new_n558), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  AND2_X1   g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n549), .A2(new_n606), .B1(KEYINPUT41), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n607), .A2(KEYINPUT41), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT101), .ZN(new_n613));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n611), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G57gat), .B(G64gat), .Z(new_n617));
  INV_X1    g416(.A(KEYINPUT9), .ZN(new_n618));
  INV_X1    g417(.A(G71gat), .ZN(new_n619));
  INV_X1    g418(.A(G78gat), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G71gat), .B(G78gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G127gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n557), .B1(new_n625), .B2(new_n624), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n209), .ZN(new_n633));
  XOR2_X1   g432(.A(G183gat), .B(G211gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n631), .B(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n616), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n604), .A2(new_n624), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n604), .A2(new_n624), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(G230gat), .A3(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n643), .A3(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT102), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n638), .A2(new_n643), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n638), .A2(new_n647), .A3(new_n643), .A4(new_n639), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT103), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n653), .A3(new_n650), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n642), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  OR2_X1    g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n651), .A2(new_n641), .A3(new_n658), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n637), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n595), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n460), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n370), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G8gat), .B1(new_n665), .B2(new_n369), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  MUX2_X1   g471(.A(new_n670), .B(new_n672), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n665), .B2(new_n527), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n417), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n665), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n665), .A2(new_n501), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n636), .A3(new_n616), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT104), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n595), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(G29gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n684), .A3(new_n460), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT45), .ZN(new_n686));
  INV_X1    g485(.A(new_n616), .ZN(new_n687));
  AND4_X1   g486(.A1(new_n517), .A2(new_n498), .A3(new_n501), .A4(new_n513), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n517), .B1(new_n516), .B2(new_n498), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n529), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n469), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT106), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n695), .B(KEYINPUT44), .C1(new_n530), .C2(new_n687), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n690), .A2(KEYINPUT107), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n519), .A2(new_n700), .A3(new_n529), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n469), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n687), .A2(KEYINPUT44), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n698), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n700), .B1(new_n519), .B2(new_n529), .ZN(new_n706));
  AOI211_X1 g505(.A(KEYINPUT107), .B(new_n528), .C1(new_n515), .C2(new_n518), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n691), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(KEYINPUT108), .A3(new_n703), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n697), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n661), .B(KEYINPUT105), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n581), .A2(new_n584), .B1(new_n589), .B2(new_n570), .ZN(new_n712));
  INV_X1    g511(.A(new_n636), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n710), .A2(KEYINPUT109), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT109), .B1(new_n710), .B2(new_n714), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n715), .A2(new_n716), .A3(new_n461), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n686), .B1(new_n717), .B2(new_n684), .ZN(G1328gat));
  NOR3_X1   g517(.A1(new_n682), .A2(new_n369), .A3(new_n538), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT46), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n715), .A2(new_n716), .A3(new_n369), .ZN(new_n721));
  INV_X1    g520(.A(new_n538), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n683), .A2(new_n724), .A3(new_n467), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n715), .A2(new_n716), .A3(new_n527), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(new_n724), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n710), .A2(new_n714), .ZN(new_n732));
  OAI21_X1  g531(.A(G43gat), .B1(new_n732), .B2(new_n527), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n726), .B1(new_n733), .B2(new_n725), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n730), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n527), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n710), .A2(KEYINPUT109), .A3(new_n714), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n727), .B1(new_n741), .B2(G43gat), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT110), .B1(new_n742), .B2(new_n734), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n743), .ZN(G1330gat));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n501), .A2(G50gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n682), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n710), .A2(new_n287), .A3(new_n714), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n745), .B(new_n747), .C1(new_n748), .C2(G50gat), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n749), .A2(KEYINPUT111), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(KEYINPUT111), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n738), .A2(new_n287), .A3(new_n740), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n747), .B1(new_n752), .B2(G50gat), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n750), .A2(new_n751), .B1(new_n753), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g553(.A1(new_n708), .A2(new_n712), .A3(new_n637), .A4(new_n711), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n461), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n756), .B(G57gat), .Z(G1332gat));
  XOR2_X1   g556(.A(new_n755), .B(KEYINPUT112), .Z(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n370), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT49), .B(G64gat), .Z(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(G1333gat));
  NAND3_X1  g561(.A1(new_n758), .A2(G71gat), .A3(new_n739), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n619), .B1(new_n755), .B2(new_n417), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g565(.A1(new_n758), .A2(new_n287), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G78gat), .ZN(G1335gat));
  INV_X1    g567(.A(new_n712), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n713), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n708), .A2(new_n616), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n661), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n599), .A3(new_n460), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n710), .A2(new_n661), .A3(new_n770), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT113), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(new_n460), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n778), .B2(new_n599), .ZN(G1336gat));
  OAI21_X1  g578(.A(G92gat), .B1(new_n776), .B2(new_n369), .ZN(new_n780));
  INV_X1    g579(.A(new_n711), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n781), .A2(G92gat), .A3(new_n369), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT115), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n784), .A2(KEYINPUT115), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n780), .A2(new_n783), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n773), .A2(KEYINPUT114), .A3(new_n782), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n776), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n792), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n370), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n791), .B1(new_n795), .B2(G92gat), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n787), .B1(new_n796), .B2(new_n784), .ZN(G1337gat));
  INV_X1    g596(.A(G99gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n774), .A2(new_n798), .A3(new_n467), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n777), .A2(new_n739), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(new_n798), .ZN(G1338gat));
  NOR3_X1   g600(.A1(new_n781), .A2(G106gat), .A3(new_n501), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n773), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(KEYINPUT53), .ZN(new_n804));
  OAI21_X1  g603(.A(G106gat), .B1(new_n776), .B2(new_n501), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n793), .A2(new_n287), .A3(new_n794), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n803), .B1(new_n807), .B2(G106gat), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(G1339gat));
  AND2_X1   g609(.A1(new_n559), .A2(new_n561), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n811), .A2(new_n560), .B1(new_n577), .B2(new_n576), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n581), .A2(new_n584), .B1(new_n569), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n661), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n815));
  NAND3_X1  g614(.A1(new_n652), .A2(new_n654), .A3(new_n815), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n649), .A2(new_n650), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n649), .B2(new_n650), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n658), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n816), .A2(new_n820), .A3(KEYINPUT55), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n660), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n821), .A2(new_n827), .A3(new_n822), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n824), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n814), .B1(new_n829), .B2(new_n712), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n687), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n830), .A2(new_n687), .B1(new_n831), .B2(new_n813), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n832), .A2(new_n713), .B1(new_n769), .B2(new_n663), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n460), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n287), .A2(new_n417), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n834), .A2(new_n370), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n769), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n370), .A2(new_n461), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n833), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n380), .B1(new_n594), .B2(new_n592), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(G1340gat));
  AOI21_X1  g641(.A(G120gat), .B1(new_n837), .B2(new_n661), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n781), .A2(new_n378), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n840), .B2(new_n844), .ZN(G1341gat));
  NAND3_X1  g644(.A1(new_n837), .A2(new_n373), .A3(new_n713), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n840), .A2(new_n713), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n846), .B1(new_n373), .B2(new_n847), .ZN(G1342gat));
  NAND3_X1  g647(.A1(new_n837), .A2(new_n371), .A3(new_n616), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(KEYINPUT56), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT118), .Z(new_n851));
  AOI21_X1  g650(.A(new_n371), .B1(new_n840), .B2(new_n616), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n849), .B2(KEYINPUT56), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1343gat));
  INV_X1    g653(.A(new_n834), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n739), .A2(new_n370), .A3(new_n501), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n594), .A2(new_n592), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n858), .A2(new_n217), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(KEYINPUT58), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n839), .A2(new_n527), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n663), .A2(new_n769), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n830), .A2(new_n687), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n831), .A2(new_n813), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n866), .B2(new_n636), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(KEYINPUT57), .A3(new_n501), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n821), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n825), .A2(new_n660), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT120), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n826), .A2(new_n874), .A3(new_n870), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n873), .B(new_n875), .C1(new_n593), .C2(new_n591), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n616), .B1(new_n876), .B2(new_n814), .ZN(new_n877));
  INV_X1    g676(.A(new_n865), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n636), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n287), .B1(new_n880), .B2(new_n863), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n862), .B(new_n868), .C1(new_n881), .C2(KEYINPUT57), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(KEYINPUT121), .A3(new_n859), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n214), .B2(new_n213), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT121), .B1(new_n882), .B2(new_n859), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n861), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n882), .A2(new_n769), .B1(new_n204), .B2(new_n206), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT58), .B1(new_n887), .B2(new_n860), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1344gat));
  NAND3_X1  g688(.A1(new_n858), .A2(new_n215), .A3(new_n661), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n501), .A2(KEYINPUT57), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n664), .A2(new_n592), .A3(new_n594), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n879), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n833), .B2(new_n287), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n899), .A2(new_n662), .A3(new_n862), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n900), .A2(KEYINPUT122), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n215), .B1(new_n900), .B2(KEYINPUT122), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n891), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n215), .C1(new_n882), .C2(new_n661), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n890), .B1(new_n903), .B2(new_n904), .ZN(G1345gat));
  NOR3_X1   g704(.A1(new_n857), .A2(G155gat), .A3(new_n636), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n882), .A2(new_n713), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(G155gat), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT123), .ZN(G1346gat));
  AOI21_X1  g708(.A(G162gat), .B1(new_n858), .B2(new_n616), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n687), .A2(new_n210), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n882), .B2(new_n911), .ZN(G1347gat));
  NAND2_X1  g711(.A1(new_n370), .A2(new_n461), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n836), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n833), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n769), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n859), .A2(G169gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n915), .B2(new_n781), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n662), .A2(G176gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n915), .B2(new_n921), .ZN(G1349gat));
  NOR3_X1   g721(.A1(new_n915), .A2(KEYINPUT27), .A3(new_n636), .ZN(new_n923));
  XOR2_X1   g722(.A(KEYINPUT60), .B(G183gat), .Z(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(G1350gat));
  OAI22_X1  g724(.A1(new_n915), .A2(new_n687), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n926));
  NAND2_X1  g725(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(G1351gat));
  NOR2_X1   g727(.A1(new_n867), .A2(new_n501), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n739), .A2(new_n913), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n769), .ZN(new_n933));
  INV_X1    g732(.A(new_n930), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n899), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n859), .A2(G197gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1352gat));
  NOR3_X1   g736(.A1(new_n931), .A2(G204gat), .A3(new_n662), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT124), .Z(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n940));
  INV_X1    g739(.A(new_n935), .ZN(new_n941));
  OAI21_X1  g740(.A(G204gat), .B1(new_n941), .B2(new_n781), .ZN(new_n942));
  XOR2_X1   g741(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n943));
  OAI211_X1 g742(.A(new_n940), .B(new_n942), .C1(new_n939), .C2(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n932), .A2(new_n241), .A3(new_n713), .ZN(new_n945));
  INV_X1    g744(.A(G211gat), .ZN(new_n946));
  NOR4_X1   g745(.A1(new_n895), .A2(new_n897), .A3(new_n636), .A4(new_n934), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n879), .A2(new_n894), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n892), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT57), .B1(new_n867), .B2(new_n501), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n951), .A2(new_n952), .A3(new_n713), .A4(new_n930), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT126), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n898), .A2(new_n948), .A3(new_n713), .A4(new_n930), .ZN(new_n956));
  AND4_X1   g755(.A1(KEYINPUT63), .A2(new_n954), .A3(G211gat), .A4(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n945), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT127), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n960), .B(new_n945), .C1(new_n955), .C2(new_n957), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n941), .B2(new_n687), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n932), .A2(new_n224), .A3(new_n616), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


