//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n452), .A2(G567), .B1(G2106), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n459), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(new_n468), .ZN(G160));
  OAI21_X1  g044(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G112), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G2105), .ZN(new_n472));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n459), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT67), .Z(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n478));
  AOI211_X1 g053(.A(new_n472), .B(new_n477), .C1(G136), .C2(new_n478), .ZN(G162));
  OAI21_X1  g054(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G114), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n486), .A2(KEYINPUT68), .A3(G126), .A4(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n482), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n486), .A2(new_n491), .A3(G138), .A4(new_n459), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  AND2_X1   g070(.A1(KEYINPUT69), .A2(KEYINPUT5), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT69), .A2(KEYINPUT5), .ZN(new_n497));
  OAI211_X1 g072(.A(KEYINPUT70), .B(G543), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT69), .A2(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(KEYINPUT70), .B1(new_n499), .B2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n498), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(new_n499), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  INV_X1    g090(.A(new_n513), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n507), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n510), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  XNOR2_X1  g096(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n522), .B(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(G51), .B2(new_n514), .ZN(new_n525));
  OAI21_X1  g100(.A(G543), .B1(new_n496), .B2(new_n497), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n505), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n513), .B1(new_n527), .B2(new_n498), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n525), .A2(new_n529), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AND2_X1   g107(.A1(new_n507), .A2(G64), .ZN(new_n533));
  AND2_X1   g108(.A1(G77), .A2(G543), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n528), .A2(G90), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n514), .A2(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(KEYINPUT72), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n536), .B2(new_n537), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n535), .B1(new_n539), .B2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND3_X1  g118(.A1(new_n507), .A2(G81), .A3(new_n516), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n514), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  AND2_X1   g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n507), .B2(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n550), .B2(new_n509), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n527), .B2(new_n498), .ZN(new_n553));
  OAI211_X1 g128(.A(KEYINPUT73), .B(G651), .C1(new_n553), .C2(new_n549), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n547), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT75), .Z(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n507), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI211_X1 g141(.A(KEYINPUT76), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n566), .B1(new_n527), .B2(new_n498), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n569), .B2(new_n563), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(G651), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n517), .A2(KEYINPUT74), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n528), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n574), .A3(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n514), .A2(G53), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n571), .A2(new_n575), .A3(new_n577), .ZN(G299));
  OAI21_X1  g153(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n514), .A2(G49), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n572), .A2(new_n574), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n572), .A2(new_n574), .A3(G86), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n527), .B2(new_n498), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n514), .A2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g169(.A1(new_n585), .A2(KEYINPUT77), .A3(new_n591), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n509), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  INV_X1    g174(.A(new_n514), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT78), .B(G47), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n517), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n514), .A2(G54), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT79), .B(G66), .Z(new_n607));
  AOI22_X1  g182(.A1(new_n507), .A2(new_n607), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n606), .B1(new_n608), .B2(new_n509), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n572), .A2(new_n574), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI211_X1 g187(.A(KEYINPUT74), .B(new_n513), .C1(new_n527), .C2(new_n498), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n573), .B1(new_n507), .B2(new_n516), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n615), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n609), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT80), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n605), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n605), .B1(new_n618), .B2(G868), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  INV_X1    g196(.A(G299), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G297));
  OAI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n618), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n486), .A2(new_n466), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n478), .A2(G135), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n459), .A2(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n475), .A2(new_n638), .A3(G123), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n638), .B1(new_n475), .B2(G123), .ZN(new_n640));
  OAI221_X1 g215(.A(new_n635), .B1(new_n636), .B2(new_n637), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  AOI22_X1  g216(.A1(new_n634), .A2(G2100), .B1(G2096), .B2(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n642), .B(new_n643), .C1(G2100), .C2(new_n634), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(G156));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT85), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(G14), .B1(new_n653), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n653), .ZN(G401));
  XOR2_X1   g237(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n666), .B2(new_n663), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n669), .B(new_n671), .Z(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1971), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n695), .A2(G23), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G288), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT33), .B(G1976), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n702), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n698), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(G305), .A2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G6), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G16), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT32), .B(G1981), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n709), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n706), .B(new_n711), .C1(new_n707), .C2(G16), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n705), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n714));
  AOI22_X1  g289(.A1(G119), .A2(new_n475), .B1(new_n478), .B2(G131), .ZN(new_n715));
  NOR2_X1   g290(.A1(G95), .A2(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT87), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n715), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G25), .B(new_n722), .S(G29), .Z(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT35), .B(G1991), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT89), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n695), .A2(G24), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n728), .B(new_n729), .C1(new_n603), .C2(new_n695), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n726), .B1(G1986), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G1986), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n713), .B2(KEYINPUT34), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n714), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n734), .A2(new_n735), .A3(KEYINPUT36), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT91), .B(KEYINPUT36), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n714), .B2(new_n733), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G160), .A2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n741), .B2(KEYINPUT24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(KEYINPUT24), .B2(new_n741), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n740), .A2(G2084), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G29), .A2(G33), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT94), .Z(new_n746));
  AND2_X1   g321(.A1(new_n486), .A2(G127), .ZN(new_n747));
  AND2_X1   g322(.A1(G115), .A2(G2104), .ZN(new_n748));
  OAI21_X1  g323(.A(G2105), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n750));
  NAND2_X1  g325(.A1(G103), .A2(G2104), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n478), .A2(G139), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n746), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n744), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT95), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n475), .A2(G129), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n466), .A2(G105), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G141), .B2(new_n478), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT96), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT26), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(new_n756), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(KEYINPUT97), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G29), .B2(G32), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n771), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n759), .B(new_n761), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(KEYINPUT98), .ZN(new_n778));
  NOR2_X1   g353(.A1(G168), .A2(new_n695), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n695), .B2(G21), .ZN(new_n780));
  INV_X1    g355(.A(G1966), .ZN(new_n781));
  INV_X1    g356(.A(new_n776), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n780), .A2(new_n781), .B1(new_n774), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G2078), .ZN(new_n784));
  NOR2_X1   g359(.A1(G164), .A2(new_n756), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G27), .B2(new_n756), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n783), .B1(new_n781), .B2(new_n780), .C1(new_n784), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n756), .A2(G35), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G162), .B2(new_n756), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT29), .B(G2090), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(G2084), .B1(new_n740), .B2(new_n743), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n786), .B2(new_n784), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT31), .B(G11), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT99), .B(G28), .Z(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(KEYINPUT30), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT30), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(new_n756), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n794), .B1(new_n796), .B2(new_n798), .C1(new_n641), .C2(new_n756), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT100), .Z(new_n800));
  NAND3_X1  g375(.A1(new_n791), .A2(new_n793), .A3(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n778), .A2(new_n787), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n695), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n622), .B2(new_n695), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n777), .A2(KEYINPUT98), .B1(G1956), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n802), .B(new_n806), .C1(G1956), .C2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n695), .A2(G5), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G171), .B2(new_n695), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT101), .ZN(new_n810));
  INV_X1    g385(.A(G1961), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n695), .A2(G4), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n618), .B2(new_n695), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G1348), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(G1348), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n695), .A2(G19), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n556), .B2(new_n695), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G1341), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n756), .A2(G26), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT92), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT28), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n478), .A2(G140), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n475), .A2(G128), .ZN(new_n825));
  OR2_X1    g400(.A1(G104), .A2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n823), .B1(new_n829), .B2(new_n756), .ZN(new_n830));
  INV_X1    g405(.A(G2067), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n816), .A2(new_n817), .A3(new_n820), .A4(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT93), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n813), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n739), .A2(new_n837), .ZN(G311));
  AND2_X1   g413(.A1(new_n813), .A2(new_n836), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n839), .A2(new_n835), .A3(new_n738), .A4(new_n736), .ZN(G150));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n841));
  AND2_X1   g416(.A1(G80), .A2(G543), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n507), .B2(G67), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n843), .B2(new_n509), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n507), .A2(G93), .A3(new_n516), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n514), .A2(G55), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G67), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n527), .B2(new_n498), .ZN(new_n849));
  OAI211_X1 g424(.A(KEYINPUT102), .B(G651), .C1(new_n849), .C2(new_n842), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n844), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT103), .B(G860), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n618), .A2(G559), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n555), .A2(new_n851), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n555), .A2(new_n851), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n857), .B(KEYINPUT38), .ZN(new_n864));
  INV_X1    g439(.A(new_n862), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n856), .B1(new_n871), .B2(new_n852), .ZN(new_n872));
  AOI211_X1 g447(.A(KEYINPUT104), .B(new_n853), .C1(new_n868), .C2(new_n870), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n855), .B1(new_n872), .B2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n722), .B(new_n632), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n769), .B(new_n755), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT105), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT105), .B1(new_n490), .B2(new_n492), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n488), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n829), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n475), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n459), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(G142), .B2(new_n478), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n881), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n877), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n641), .B(G160), .ZN(new_n889));
  XNOR2_X1  g464(.A(G162), .B(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n890), .B2(new_n888), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g468(.A(new_n862), .B(KEYINPUT106), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n627), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT107), .B1(new_n617), .B2(G299), .ZN(new_n896));
  INV_X1    g471(.A(new_n609), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT10), .B1(new_n615), .B2(G92), .ZN(new_n898));
  AND4_X1   g473(.A1(KEYINPUT10), .A2(new_n572), .A3(G92), .A4(new_n574), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n622), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n617), .A2(G299), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n896), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT41), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n896), .A2(new_n902), .A3(new_n906), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n895), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G305), .A2(G290), .ZN(new_n911));
  XNOR2_X1  g486(.A(G288), .B(G303), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n603), .B1(new_n594), .B2(new_n595), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n904), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n895), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n910), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n910), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(G868), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G868), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n851), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(G295));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n925), .ZN(G331));
  OAI21_X1  g502(.A(G651), .B1(new_n553), .B2(new_n549), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n546), .B1(new_n548), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n845), .A2(new_n846), .ZN(new_n930));
  OAI21_X1  g505(.A(G651), .B1(new_n849), .B2(new_n842), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n841), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n929), .A2(new_n932), .A3(new_n554), .A4(new_n850), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n555), .A2(new_n851), .ZN(new_n934));
  NAND2_X1  g509(.A1(G168), .A2(KEYINPUT108), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(G301), .B1(KEYINPUT108), .B2(G168), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n940));
  NAND2_X1  g515(.A1(G286), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(G301), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n935), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n860), .B2(new_n861), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n939), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT109), .B1(new_n908), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n904), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n938), .B1(new_n936), .B2(new_n937), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n944), .A2(new_n942), .A3(new_n945), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n905), .A4(new_n907), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n948), .A2(new_n916), .A3(new_n949), .A4(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n948), .A2(new_n949), .A3(new_n954), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n914), .B2(new_n915), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT43), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n956), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n952), .A2(new_n905), .A3(new_n907), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n962), .A2(KEYINPUT110), .B1(new_n904), .B2(new_n947), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n909), .A2(new_n964), .A3(new_n952), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n916), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n961), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT44), .B1(new_n960), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n967), .B1(new_n957), .B2(new_n959), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n961), .A2(new_n966), .A3(KEYINPUT43), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(G397));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n465), .A2(new_n467), .ZN(new_n976));
  INV_X1    g551(.A(G125), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n473), .B2(new_n474), .ZN(new_n978));
  INV_X1    g553(.A(new_n463), .ZN(new_n979));
  OAI21_X1  g554(.A(G2105), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n980), .A3(G40), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND3_X1  g559(.A1(G160), .A2(KEYINPUT111), .A3(G40), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n880), .A2(new_n983), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n975), .B1(new_n986), .B2(G8), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n975), .A3(G8), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  NOR2_X1   g566(.A1(G288), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n990), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n988), .B2(new_n989), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT114), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n993), .A2(new_n997), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n988), .A2(new_n989), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n528), .A2(G86), .ZN(new_n1002));
  OAI21_X1  g577(.A(G1981), .B1(new_n591), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1981), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n584), .A2(new_n589), .A3(new_n1004), .A4(new_n590), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT49), .B1(new_n1007), .B2(KEYINPUT116), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT115), .B1(KEYINPUT116), .B2(KEYINPUT49), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1001), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(KEYINPUT117), .B(new_n1001), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n880), .A2(new_n1017), .A3(new_n984), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n494), .A2(new_n984), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT50), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n983), .A2(new_n985), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1022), .A2(G2090), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n880), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1384), .B1(new_n488), .B2(new_n493), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1024), .B(new_n1021), .C1(KEYINPUT45), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1971), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1016), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G303), .A2(G8), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1000), .A2(new_n1015), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1005), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G288), .A2(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n1015), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n990), .B(KEYINPUT118), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1034), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n880), .A2(new_n984), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT50), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1025), .A2(KEYINPUT119), .A3(new_n1017), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1041), .A2(new_n1021), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1028), .B1(new_n1045), .B2(G2090), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1032), .B1(new_n1046), .B2(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1033), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1021), .B1(new_n1049), .B2(new_n1019), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n880), .B2(new_n984), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n781), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G2084), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1016), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1055), .A2(G168), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1000), .A2(new_n1048), .A3(new_n1015), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1000), .A2(new_n1015), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1056), .B1(new_n1032), .B2(new_n1029), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1061), .A2(new_n1058), .A3(new_n1033), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1039), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1066));
  OAI211_X1 g641(.A(G8), .B(new_n1065), .C1(new_n1066), .C2(G286), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1055), .A2(G286), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G168), .A2(new_n1016), .ZN(new_n1070));
  AND2_X1   g645(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1071), .A2(new_n1065), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1055), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT62), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  OR3_X1    g649(.A1(new_n1055), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n1068), .A4(new_n1067), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  OR4_X1    g653(.A1(new_n1078), .A2(new_n1050), .A3(G2078), .A4(new_n1051), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1022), .A2(new_n811), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1026), .B2(G2078), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1082), .A2(G171), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1074), .A2(new_n1077), .A3(new_n1083), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT56), .B(G2072), .Z(new_n1085));
  OR2_X1    g660(.A1(new_n1026), .A2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1025), .A2(KEYINPUT119), .A3(new_n1017), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n1025), .B2(new_n1017), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n983), .A2(new_n985), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1040), .B2(KEYINPUT50), .ZN(new_n1091));
  AOI211_X1 g666(.A(KEYINPUT120), .B(G1956), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n1093));
  INV_X1    g668(.A(G1956), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1045), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1086), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(G299), .B(KEYINPUT57), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1021), .A2(KEYINPUT121), .A3(new_n984), .A4(new_n880), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n986), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1348), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1102), .A2(new_n831), .B1(new_n1103), .B2(new_n1022), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n900), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1097), .B(KEYINPUT122), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1098), .A2(new_n1105), .B1(new_n1096), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(new_n831), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1022), .A2(new_n1103), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n1109), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n900), .A2(KEYINPUT124), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n617), .B(KEYINPUT124), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n1104), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT58), .B(G1341), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1102), .A2(new_n1119), .B1(G1996), .B2(new_n1026), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n556), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(KEYINPUT123), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1120), .B(new_n556), .C1(KEYINPUT123), .C2(new_n1122), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT61), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1118), .B(new_n1126), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1096), .A2(KEYINPUT61), .A3(new_n1097), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1107), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G301), .B(KEYINPUT54), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1051), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n981), .A2(new_n1078), .A3(G2078), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n1024), .A3(new_n1136), .ZN(new_n1137));
  AND4_X1   g712(.A1(new_n1080), .A2(new_n1134), .A3(new_n1081), .A4(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1082), .A2(new_n1133), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1132), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1084), .B1(new_n1131), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1060), .A2(new_n1048), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1064), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1135), .A2(new_n1090), .ZN(new_n1144));
  INV_X1    g719(.A(G1996), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n769), .B(new_n1145), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n722), .A2(new_n724), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n828), .B(new_n831), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n722), .A2(new_n724), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n603), .B(G1986), .Z(new_n1151));
  OAI21_X1  g726(.A(new_n1144), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1143), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(G290), .A2(G1986), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT48), .B1(new_n1144), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1144), .A2(new_n1154), .A3(KEYINPUT48), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1155), .B(new_n1156), .C1(new_n1144), .C2(new_n1150), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT46), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1148), .A2(new_n765), .A3(new_n768), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1144), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1144), .A2(KEYINPUT46), .A3(new_n1145), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1161), .A2(KEYINPUT126), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(KEYINPUT126), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT47), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1166), .A2(new_n1147), .B1(G2067), .B2(new_n828), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1157), .B(new_n1165), .C1(new_n1144), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1153), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g744(.A1(new_n971), .A2(new_n972), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n674), .A2(G319), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1172), .A2(G401), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n693), .A2(new_n1173), .ZN(new_n1174));
  AND2_X1   g748(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1176));
  OAI21_X1  g750(.A(new_n892), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g751(.A1(new_n1171), .A2(new_n1177), .ZN(G308));
  OAI221_X1 g752(.A(new_n892), .B1(new_n1175), .B2(new_n1176), .C1(new_n971), .C2(new_n972), .ZN(G225));
endmodule


