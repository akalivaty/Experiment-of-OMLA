//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT0), .A4(G128), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n190), .A2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n188), .A2(G143), .ZN(new_n199));
  OAI211_X1 g013(.A(G128), .B(new_n197), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n189), .B(new_n191), .C1(KEYINPUT1), .C2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n196), .B1(new_n204), .B2(G125), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n206));
  INV_X1    g020(.A(G224), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G953), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n205), .B1(new_n206), .B2(new_n208), .ZN(new_n210));
  XNOR2_X1  g024(.A(G110), .B(G122), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n211), .B(KEYINPUT82), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n213));
  XNOR2_X1  g027(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G104), .ZN(new_n219));
  INV_X1    g033(.A(G101), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(G107), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n216), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n215), .A2(G107), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(G101), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G116), .ZN(new_n229));
  INV_X1    g043(.A(G116), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  OR2_X1    g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT5), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(G113), .B1(new_n229), .B2(KEYINPUT5), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n214), .B1(new_n227), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n235), .B2(KEYINPUT85), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(KEYINPUT85), .B2(new_n235), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n226), .B1(new_n241), .B2(new_n234), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n209), .B(new_n210), .C1(new_n239), .C2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n216), .A2(new_n219), .A3(new_n221), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n232), .B(new_n233), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n248), .A3(G101), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT81), .A4(new_n249), .ZN(new_n253));
  OR2_X1    g067(.A1(new_n238), .A2(new_n226), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(new_n212), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n187), .B1(new_n243), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n258), .A3(new_n212), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT83), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT83), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n255), .A2(new_n261), .A3(new_n258), .A4(new_n212), .ZN(new_n262));
  INV_X1    g076(.A(new_n256), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n258), .B1(new_n255), .B2(new_n212), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n260), .A2(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n205), .B(new_n208), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n257), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT87), .ZN(new_n268));
  OAI21_X1  g082(.A(G210), .B1(G237), .B2(G902), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(KEYINPUT86), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n269), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT87), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n270), .A2(KEYINPUT86), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n267), .A2(KEYINPUT87), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G214), .B1(G237), .B2(G902), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT80), .ZN(new_n280));
  INV_X1    g094(.A(G469), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(new_n187), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT64), .ZN(new_n283));
  INV_X1    g097(.A(G137), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(KEYINPUT64), .A2(G137), .ZN(new_n286));
  AND2_X1   g100(.A1(KEYINPUT11), .A2(G134), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT11), .B1(new_n284), .B2(G134), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G134), .ZN(new_n291));
  AOI21_X1  g105(.A(G131), .B1(new_n291), .B2(G137), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT65), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT65), .A4(new_n292), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n288), .B(new_n290), .C1(G134), .C2(new_n284), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n295), .A2(new_n296), .B1(G131), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT10), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n204), .A2(new_n227), .A3(KEYINPUT78), .A4(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n200), .A2(new_n222), .A3(new_n225), .A4(new_n202), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n193), .A2(new_n194), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n249), .A2(new_n305), .A3(new_n192), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT77), .B1(new_n306), .B2(new_n246), .ZN(new_n307));
  INV_X1    g121(.A(new_n195), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n246), .A2(KEYINPUT77), .A3(new_n308), .A4(new_n249), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n298), .B(new_n304), .C1(new_n307), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT12), .ZN(new_n312));
  AND4_X1   g126(.A1(new_n202), .A2(new_n200), .A3(new_n222), .A4(new_n225), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n202), .A2(new_n200), .B1(new_n222), .B2(new_n225), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n312), .B1(new_n315), .B2(new_n298), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n297), .A2(G131), .ZN(new_n317));
  AND2_X1   g131(.A1(KEYINPUT64), .A2(G137), .ZN(new_n318));
  NOR2_X1   g132(.A1(KEYINPUT64), .A2(G137), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n289), .B1(new_n320), .B2(new_n287), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT65), .B1(new_n321), .B2(new_n292), .ZN(new_n322));
  INV_X1    g136(.A(new_n296), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n203), .A2(new_n226), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n301), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n324), .A2(KEYINPUT79), .A3(KEYINPUT12), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n316), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n295), .A2(new_n296), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n329), .A2(new_n317), .B1(new_n325), .B2(new_n301), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT79), .B1(new_n330), .B2(KEYINPUT12), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n311), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G140), .ZN(new_n333));
  INV_X1    g147(.A(G227), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G953), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT76), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n249), .A2(new_n305), .A3(new_n192), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n341), .A2(new_n309), .B1(new_n300), .B2(new_n303), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n336), .B1(new_n342), .B2(new_n298), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n304), .B1(new_n307), .B2(new_n310), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n324), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n332), .A2(new_n337), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n282), .B1(new_n346), .B2(G469), .ZN(new_n347));
  INV_X1    g161(.A(new_n336), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n311), .B(new_n348), .C1(new_n328), .C2(new_n331), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n348), .B1(new_n345), .B2(new_n311), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n281), .B(new_n187), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT9), .B(G234), .ZN(new_n354));
  OAI21_X1  g168(.A(G221), .B1(new_n354), .B2(G902), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n280), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n355), .ZN(new_n357));
  AOI211_X1 g171(.A(KEYINPUT80), .B(new_n357), .C1(new_n347), .C2(new_n352), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G113), .B(G122), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(new_n215), .ZN(new_n361));
  XNOR2_X1  g175(.A(G125), .B(G140), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT16), .ZN(new_n363));
  INV_X1    g177(.A(G125), .ZN(new_n364));
  OR3_X1    g178(.A1(new_n364), .A2(KEYINPUT16), .A3(G140), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(G146), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT74), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(KEYINPUT74), .A3(new_n365), .A4(G146), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n363), .A2(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n188), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(G237), .A2(G953), .ZN(new_n374));
  AOI21_X1  g188(.A(G143), .B1(new_n374), .B2(G214), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(G143), .A3(G214), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT17), .A3(G131), .ZN(new_n379));
  INV_X1    g193(.A(new_n377), .ZN(new_n380));
  OAI21_X1  g194(.A(G131), .B1(new_n380), .B2(new_n375), .ZN(new_n381));
  INV_X1    g195(.A(G131), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n382), .A3(new_n377), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT89), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT89), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(new_n383), .A3(new_n387), .A4(new_n384), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n373), .A2(new_n379), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n380), .A2(new_n375), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT18), .A2(G131), .ZN(new_n391));
  XOR2_X1   g205(.A(G125), .B(G140), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G146), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n362), .A2(new_n188), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n390), .A2(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n378), .A2(KEYINPUT18), .A3(G131), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n361), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n389), .A2(new_n399), .A3(new_n361), .A4(new_n397), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n386), .A2(new_n388), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n368), .A2(new_n379), .A3(new_n371), .A4(new_n369), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n361), .B(new_n397), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT90), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n398), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G475), .B1(new_n405), .B2(G902), .ZN(new_n406));
  NOR2_X1   g220(.A1(G475), .A2(G902), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n400), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n362), .B(KEYINPUT19), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n188), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n381), .A2(new_n383), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n366), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n361), .B1(new_n413), .B2(new_n397), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n415), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n408), .B1(new_n409), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(KEYINPUT91), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n400), .A2(new_n404), .B1(new_n416), .B2(new_n417), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT20), .B1(new_n422), .B2(new_n408), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT91), .B1(new_n419), .B2(new_n420), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n406), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G478), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(KEYINPUT15), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n190), .A2(G128), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n201), .A2(G143), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(new_n291), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n230), .A2(KEYINPUT14), .A3(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(G116), .B(G122), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(G107), .B(new_n433), .C1(new_n435), .C2(KEYINPUT14), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n432), .B(new_n436), .C1(G107), .C2(new_n435), .ZN(new_n437));
  INV_X1    g251(.A(new_n429), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n438), .A2(KEYINPUT13), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n430), .B1(new_n438), .B2(KEYINPUT13), .ZN(new_n440));
  OAI21_X1  g254(.A(G134), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n431), .A2(new_n291), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n434), .B(new_n218), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n437), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G217), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n354), .A2(new_n446), .A3(G953), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n445), .B(new_n447), .Z(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n187), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT92), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n428), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n450), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(KEYINPUT92), .A3(new_n187), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(new_n454), .B2(new_n428), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT93), .B(G952), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(G953), .ZN(new_n457));
  NAND2_X1  g271(.A1(G234), .A2(G237), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n458), .A2(G902), .A3(G953), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(G898), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  NOR4_X1   g278(.A1(new_n279), .A2(new_n359), .A3(new_n426), .A4(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G472), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n187), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT66), .B1(new_n320), .B2(G134), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n284), .A2(G134), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT66), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n471), .B(new_n291), .C1(new_n318), .C2(new_n319), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n473), .A2(G131), .B1(new_n295), .B2(new_n296), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n204), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n324), .A2(new_n308), .ZN(new_n476));
  INV_X1    g290(.A(new_n247), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n374), .A2(G210), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT27), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT26), .B(G101), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n298), .A2(new_n195), .ZN(new_n487));
  AOI21_X1  g301(.A(G134), .B1(new_n285), .B2(new_n286), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n470), .B1(new_n488), .B2(new_n471), .ZN(new_n489));
  INV_X1    g303(.A(new_n472), .ZN(new_n490));
  OAI21_X1  g304(.A(G131), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n329), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT67), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n203), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n487), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT68), .B1(new_n496), .B2(KEYINPUT30), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n204), .B1(new_n474), .B2(KEYINPUT67), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n492), .A2(new_n493), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n476), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT68), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n475), .A2(new_n476), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n477), .B1(new_n505), .B2(KEYINPUT30), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n486), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT31), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n468), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n505), .A2(KEYINPUT30), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n247), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n503), .B2(new_n497), .ZN(new_n512));
  OAI211_X1 g326(.A(KEYINPUT69), .B(KEYINPUT31), .C1(new_n512), .C2(new_n486), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n505), .A2(new_n515), .A3(new_n477), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n478), .A2(KEYINPUT28), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n500), .A2(new_n247), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n507), .A2(new_n508), .B1(new_n484), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n467), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT70), .B1(new_n522), .B2(KEYINPUT32), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n475), .A2(new_n476), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n247), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n483), .A2(KEYINPUT29), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n187), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n484), .B1(new_n512), .B2(new_n479), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n518), .A2(new_n483), .A3(new_n519), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n529), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n524), .B1(new_n534), .B2(new_n466), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n532), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n496), .A2(KEYINPUT68), .A3(KEYINPUT30), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n501), .B1(new_n500), .B2(new_n502), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n506), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n478), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n536), .B1(new_n540), .B2(new_n484), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT71), .B(G472), .C1(new_n541), .C2(new_n529), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT70), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT32), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n520), .A2(new_n484), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n539), .A2(new_n485), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(new_n547), .B2(KEYINPUT31), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n509), .B2(new_n513), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n544), .B(new_n545), .C1(new_n549), .C2(new_n467), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n522), .A2(KEYINPUT32), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n523), .A2(new_n543), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n446), .B1(G234), .B2(new_n187), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT25), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT24), .B(G110), .Z(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT72), .ZN(new_n557));
  XNOR2_X1  g371(.A(G119), .B(G128), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT23), .B1(new_n201), .B2(G119), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT73), .B1(new_n228), .B2(G128), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n560), .B(new_n561), .Z(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G110), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n366), .B(new_n394), .C1(new_n559), .C2(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n557), .A2(new_n558), .B1(new_n562), .B2(G110), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT75), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n565), .A2(new_n566), .A3(new_n372), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(new_n565), .B2(new_n372), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n564), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT22), .B(G137), .ZN(new_n570));
  INV_X1    g384(.A(G953), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n571), .A2(G221), .A3(G234), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n570), .B(new_n572), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n564), .B(new_n573), .C1(new_n567), .C2(new_n568), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n555), .B1(new_n577), .B2(G902), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n575), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n576), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n554), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n577), .A2(G902), .A3(new_n553), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n465), .A2(new_n552), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  INV_X1    g398(.A(new_n522), .ZN(new_n585));
  AOI21_X1  g399(.A(G902), .B1(new_n514), .B2(new_n521), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n585), .B1(new_n466), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n582), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n587), .A2(new_n588), .A3(new_n359), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n272), .A2(KEYINPUT94), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n265), .A2(new_n266), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT95), .B(new_n270), .C1(new_n591), .C2(new_n257), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT95), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n267), .B2(new_n269), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT94), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n267), .A2(new_n595), .A3(new_n269), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n590), .A2(new_n592), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(new_n278), .ZN(new_n598));
  NAND2_X1  g412(.A1(G478), .A2(G902), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n449), .B2(G478), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n445), .B(new_n447), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n445), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n601), .B(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n600), .B1(G478), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n426), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n598), .A2(new_n463), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n589), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  XOR2_X1   g426(.A(new_n463), .B(KEYINPUT98), .Z(new_n613));
  INV_X1    g427(.A(new_n455), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n406), .A2(KEYINPUT97), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n406), .A2(KEYINPUT97), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n419), .A2(new_n420), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n423), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n614), .A2(new_n615), .A3(new_n616), .A4(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n598), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n589), .A2(new_n613), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  INV_X1    g437(.A(new_n587), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n574), .A2(KEYINPUT36), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n569), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n569), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n629), .A2(G902), .A3(new_n553), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n580), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n465), .A2(new_n624), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT37), .B(G110), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G12));
  NAND2_X1  g448(.A1(new_n597), .A2(new_n278), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n631), .B1(new_n358), .B2(new_n356), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(G900), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n460), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n459), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n619), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n552), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  NAND2_X1  g457(.A1(new_n526), .A2(new_n478), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT99), .B1(new_n644), .B2(new_n484), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n644), .A2(KEYINPUT99), .A3(new_n484), .ZN(new_n646));
  OR3_X1    g460(.A1(new_n507), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n466), .B1(new_n647), .B2(new_n187), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n522), .B2(KEYINPUT32), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n523), .A2(new_n649), .A3(new_n550), .ZN(new_n650));
  INV_X1    g464(.A(new_n278), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n580), .A2(new_n630), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n426), .A3(new_n614), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n277), .A2(KEYINPUT38), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT38), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n271), .A2(new_n274), .A3(new_n655), .A4(new_n276), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT100), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n640), .B(KEYINPUT39), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n660), .B1(new_n356), .B2(new_n358), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT101), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n664), .B(new_n660), .C1(new_n356), .C2(new_n358), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n663), .B1(new_n662), .B2(new_n665), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n650), .A2(new_n669), .A3(new_n657), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n659), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G143), .ZN(G45));
  INV_X1    g486(.A(new_n640), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n607), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n552), .A2(new_n637), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  OR2_X1    g490(.A1(new_n350), .A2(new_n351), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n187), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G469), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n355), .A3(new_n352), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT102), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n679), .A2(new_n682), .A3(new_n355), .A4(new_n352), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n681), .A2(new_n582), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n609), .A2(new_n552), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NAND4_X1  g501(.A1(new_n620), .A2(new_n552), .A3(new_n613), .A4(new_n684), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  NAND2_X1  g503(.A1(new_n679), .A2(new_n352), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n597), .A2(new_n278), .A3(new_n355), .A4(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n426), .ZN(new_n694));
  AND4_X1   g508(.A1(new_n694), .A2(new_n631), .A3(new_n463), .A4(new_n455), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n552), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  AOI22_X1  g511(.A1(new_n507), .A2(new_n508), .B1(new_n484), .B2(new_n527), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n547), .A2(KEYINPUT31), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n467), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n586), .B2(new_n466), .ZN(new_n702));
  OAI211_X1 g516(.A(KEYINPUT103), .B(G472), .C1(new_n549), .C2(G902), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n426), .A2(new_n614), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n635), .A2(new_n705), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n681), .A2(new_n613), .A3(new_n683), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n704), .A2(new_n582), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT104), .B(G122), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G24));
  NAND4_X1  g524(.A1(new_n704), .A2(new_n631), .A3(new_n674), .A4(new_n693), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  INV_X1    g526(.A(new_n353), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n355), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n271), .A2(new_n274), .A3(new_n278), .A4(new_n276), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n552), .A2(new_n582), .A3(new_n674), .A4(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n543), .A2(new_n551), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n585), .A2(new_n545), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n588), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n674), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n720), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  NAND4_X1  g543(.A1(new_n552), .A2(new_n582), .A3(new_n641), .A4(new_n718), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G134), .ZN(G36));
  OAI211_X1 g545(.A(new_n606), .B(new_n406), .C1(new_n424), .C2(new_n425), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n587), .A2(new_n631), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n332), .A2(new_n337), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n343), .A2(new_n345), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n281), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n741), .B2(new_n740), .ZN(new_n743));
  INV_X1    g557(.A(new_n282), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT46), .B1(new_n743), .B2(new_n744), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n352), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n355), .B(new_n660), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n717), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n587), .A2(new_n734), .A3(KEYINPUT44), .A4(new_n631), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n737), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  NAND2_X1  g570(.A1(new_n674), .A2(new_n588), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n552), .A2(new_n717), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n355), .B1(new_n748), .B2(new_n749), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(KEYINPUT47), .B(new_n355), .C1(new_n748), .C2(new_n749), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  NOR2_X1   g579(.A1(new_n717), .A2(new_n680), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT115), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n767), .A2(new_n588), .A3(new_n650), .A4(new_n459), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n608), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n457), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n704), .A2(new_n582), .ZN(new_n771));
  INV_X1    g585(.A(new_n459), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n734), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n693), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n734), .A2(new_n772), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n767), .A2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n777), .A2(KEYINPUT48), .A3(new_n724), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT48), .B1(new_n777), .B2(new_n724), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n770), .A2(new_n775), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n654), .A2(new_n656), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n278), .A3(new_n680), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n773), .A3(new_n582), .A4(new_n704), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(KEYINPUT113), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(KEYINPUT113), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n771), .A2(new_n773), .A3(new_n786), .A4(new_n782), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n752), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n691), .A2(KEYINPUT112), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n691), .A2(KEYINPUT112), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n790), .A2(new_n791), .A3(new_n355), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n774), .B(new_n789), .C1(new_n763), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n704), .A2(new_n631), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n767), .A3(new_n776), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n426), .A2(new_n606), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n795), .B1(new_n768), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n798), .A3(KEYINPUT51), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n780), .B1(new_n788), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n785), .A2(new_n787), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(new_n785), .B2(new_n787), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(KEYINPUT116), .B(new_n798), .C1(new_n802), .C2(new_n803), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n807), .A3(new_n793), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n800), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n455), .A2(new_n640), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n636), .A2(new_n717), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n552), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n730), .B(new_n814), .C1(new_n794), .C2(new_n725), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n815), .A2(KEYINPUT110), .B1(new_n721), .B2(new_n727), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n552), .B(new_n637), .C1(new_n641), .C2(new_n674), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(new_n711), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n716), .A2(new_n631), .A3(new_n673), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n650), .A2(new_n706), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT52), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n589), .A2(new_n613), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n426), .B2(new_n455), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n607), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n426), .A2(new_n824), .A3(new_n455), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(new_n279), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n632), .B(new_n696), .C1(new_n823), .C2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n688), .A2(new_n685), .A3(new_n708), .A4(new_n583), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n794), .A2(new_n725), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n730), .A3(new_n814), .A4(new_n834), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n816), .A2(new_n822), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n817), .A2(new_n711), .A3(new_n821), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT111), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT53), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n816), .A2(new_n832), .A3(new_n835), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n841), .A2(new_n842), .A3(new_n838), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n816), .A2(new_n832), .A3(new_n835), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n839), .A3(KEYINPUT53), .A4(new_n822), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n842), .B1(new_n841), .B2(new_n838), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n810), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(G952), .B2(G953), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n588), .A2(new_n732), .A3(new_n651), .A4(new_n357), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT108), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n690), .B(KEYINPUT49), .ZN(new_n854));
  OR4_X1    g668(.A1(new_n650), .A2(new_n853), .A3(new_n781), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(G75));
  NAND2_X1  g670(.A1(new_n846), .A2(new_n847), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(G210), .A3(G902), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n265), .A2(new_n266), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n591), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT55), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n862), .B1(new_n858), .B2(new_n859), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n571), .A2(G952), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G51));
  XNOR2_X1  g680(.A(new_n282), .B(KEYINPUT57), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n848), .B1(new_n846), .B2(new_n847), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n677), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n857), .A2(G902), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(new_n743), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n865), .B1(new_n871), .B2(new_n873), .ZN(G54));
  NAND2_X1  g688(.A1(KEYINPUT58), .A2(G475), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n422), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n865), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n872), .A2(new_n422), .A3(new_n875), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(G60));
  XOR2_X1   g694(.A(new_n599), .B(KEYINPUT59), .Z(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n844), .B2(new_n849), .ZN(new_n882));
  INV_X1    g696(.A(new_n605), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n605), .A2(new_n881), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n868), .B2(new_n869), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n877), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n884), .A2(new_n887), .ZN(G63));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n889));
  XOR2_X1   g703(.A(KEYINPUT117), .B(KEYINPUT60), .Z(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT119), .ZN(new_n891));
  NAND2_X1  g705(.A1(G217), .A2(G902), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT118), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n891), .B(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n846), .B2(new_n847), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n629), .B(KEYINPUT120), .Z(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n577), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n877), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n889), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n896), .A2(new_n900), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(KEYINPUT61), .A3(new_n877), .A4(new_n898), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(G66));
  OAI21_X1  g719(.A(G953), .B1(new_n461), .B2(new_n207), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n832), .B2(G953), .ZN(new_n907));
  INV_X1    g721(.A(new_n265), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(G898), .B2(new_n571), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n907), .B(new_n909), .ZN(G69));
  NAND2_X1  g724(.A1(new_n504), .A2(new_n510), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n410), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(G900), .B2(G953), .ZN(new_n913));
  INV_X1    g727(.A(new_n750), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n724), .A2(new_n706), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n818), .A2(new_n730), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n764), .A2(new_n755), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n728), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n913), .B1(new_n920), .B2(G953), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(G953), .B1(new_n334), .B2(new_n638), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n921), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n828), .A2(new_n661), .A3(new_n717), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n552), .A3(new_n582), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n764), .A2(new_n928), .A3(new_n755), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n818), .A2(new_n671), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(KEYINPUT62), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n818), .A2(new_n671), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT121), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n650), .A2(new_n669), .A3(new_n657), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n669), .B1(new_n650), .B2(new_n657), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n666), .A2(new_n667), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n817), .A2(new_n711), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT62), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n764), .A2(new_n928), .A3(new_n755), .ZN(new_n941));
  AND4_X1   g755(.A1(KEYINPUT121), .A2(new_n940), .A3(new_n933), .A4(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n571), .B1(new_n934), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n912), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n926), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(KEYINPUT122), .A3(new_n912), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n925), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n940), .A2(new_n933), .A3(new_n941), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n931), .A2(KEYINPUT121), .A3(new_n933), .ZN(new_n952));
  AOI21_X1  g766(.A(G953), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n912), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND4_X1   g769(.A1(new_n921), .A2(new_n955), .A3(new_n925), .A4(new_n947), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n948), .A2(new_n956), .ZN(G72));
  NOR2_X1   g771(.A1(new_n840), .A2(new_n843), .ZN(new_n958));
  XNOR2_X1  g772(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n466), .A2(new_n187), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n530), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n961), .B1(new_n962), .B2(new_n507), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT127), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n540), .B(KEYINPUT126), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n951), .A2(new_n952), .A3(new_n832), .ZN(new_n967));
  AOI211_X1 g781(.A(new_n484), .B(new_n966), .C1(new_n967), .C2(new_n961), .ZN(new_n968));
  INV_X1    g782(.A(new_n832), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n961), .B1(new_n920), .B2(new_n969), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n970), .A2(new_n484), .A3(new_n966), .ZN(new_n971));
  NOR4_X1   g785(.A1(new_n965), .A2(new_n968), .A3(new_n865), .A4(new_n971), .ZN(G57));
endmodule


