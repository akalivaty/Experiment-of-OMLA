//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G101), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT28), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G113), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G116), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(G119), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n202), .A2(G119), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n201), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  AND4_X1   g025(.A1(new_n211), .A2(new_n206), .A3(new_n208), .A4(new_n201), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n207), .B1(new_n198), .B2(new_n200), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n213), .B2(new_n206), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OR2_X1    g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G143), .B(G146), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G134), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G137), .ZN(new_n228));
  INV_X1    g042(.A(G137), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT64), .B1(new_n229), .B2(G134), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI211_X1 g046(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n229), .C2(G134), .ZN(new_n233));
  OAI21_X1  g047(.A(G131), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n229), .A2(G134), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n227), .B2(G137), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n235), .B1(new_n237), .B2(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n230), .A2(new_n231), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n226), .B1(new_n234), .B2(new_n241), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n232), .A2(G131), .A3(new_n233), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT1), .B1(new_n218), .B2(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n218), .A2(G146), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n216), .A2(G143), .ZN(new_n246));
  OAI211_X1 g060(.A(G128), .B(new_n244), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n217), .B(new_n219), .C1(KEYINPUT1), .C2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n227), .A2(G137), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n250), .B2(new_n235), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n247), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n243), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n215), .B1(new_n242), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n226), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n239), .B1(new_n238), .B2(new_n240), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n243), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n206), .A2(new_n208), .A3(new_n201), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n213), .A2(new_n211), .A3(new_n206), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n209), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n241), .A2(new_n249), .A3(new_n247), .A4(new_n251), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n196), .B1(new_n254), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n242), .A2(new_n253), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT28), .B1(new_n265), .B2(new_n261), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n195), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT68), .B(new_n195), .C1(new_n264), .C2(new_n266), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n242), .A2(new_n253), .A3(KEYINPUT30), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n257), .B2(new_n262), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n215), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n263), .A3(new_n194), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n263), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT30), .B1(new_n242), .B2(new_n253), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n257), .A2(new_n262), .A3(new_n273), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(new_n282), .B2(new_n215), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT31), .A3(new_n194), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n188), .B1(new_n271), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT31), .B1(new_n283), .B2(new_n194), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n261), .B1(new_n280), .B2(new_n281), .ZN(new_n288));
  NOR4_X1   g102(.A1(new_n288), .A2(new_n279), .A3(new_n277), .A4(new_n195), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n269), .B(new_n270), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT69), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n187), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n187), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n290), .A2(KEYINPUT69), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n285), .A2(new_n188), .A3(new_n269), .A4(new_n270), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n264), .ZN(new_n300));
  INV_X1    g114(.A(new_n266), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(KEYINPUT29), .A3(new_n194), .A4(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n264), .A2(new_n266), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT29), .B1(new_n306), .B2(new_n194), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n195), .B1(new_n288), .B2(new_n279), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n304), .A2(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n302), .A2(KEYINPUT71), .A3(new_n303), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n299), .A2(KEYINPUT32), .B1(G472), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT70), .B1(new_n299), .B2(KEYINPUT32), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n295), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G128), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n248), .A2(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT24), .B(G110), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT23), .B1(new_n248), .B2(G119), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n248), .A2(G119), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n248), .A2(KEYINPUT23), .A3(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n320), .B1(new_n325), .B2(G110), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n328), .A2(new_n330), .A3(KEYINPUT72), .A4(KEYINPUT16), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n328), .A2(new_n330), .A3(KEYINPUT16), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(new_n328), .B2(KEYINPUT16), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n216), .B(new_n331), .C1(new_n332), .C2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n328), .A2(new_n330), .A3(KEYINPUT16), .ZN(new_n337));
  OR3_X1    g151(.A1(new_n329), .A2(KEYINPUT16), .A3(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n333), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n216), .B1(new_n339), .B2(new_n331), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n326), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G110), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n323), .A2(KEYINPUT73), .A3(new_n342), .A4(new_n324), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n315), .B2(G128), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n345), .A2(new_n324), .A3(new_n342), .A4(new_n316), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n318), .A2(new_n319), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n343), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n331), .B1(new_n332), .B2(new_n334), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G146), .ZN(new_n352));
  XNOR2_X1  g166(.A(G125), .B(G140), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n216), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n341), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G137), .ZN(new_n357));
  INV_X1    g171(.A(G953), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(G221), .A3(G234), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n357), .B(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n341), .A2(new_n355), .A3(new_n360), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT75), .ZN(new_n365));
  INV_X1    g179(.A(G217), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(G234), .B2(new_n303), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n362), .A2(new_n303), .A3(new_n363), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT74), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(KEYINPUT74), .A3(KEYINPUT25), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n367), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  AOI22_X1  g194(.A1(KEYINPUT76), .A2(new_n379), .B1(new_n380), .B2(G107), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n382));
  INV_X1    g196(.A(G107), .ZN(new_n383));
  AND4_X1   g197(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT3), .A4(G104), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n382), .A2(KEYINPUT3), .B1(new_n383), .B2(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G101), .ZN(new_n387));
  INV_X1    g201(.A(G101), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(new_n381), .C1(new_n384), .C2(new_n385), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n390));
  OAI22_X1  g204(.A1(KEYINPUT76), .A2(new_n379), .B1(new_n380), .B2(G107), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT3), .A4(G104), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n388), .B1(new_n393), .B2(new_n381), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT77), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI22_X1  g210(.A1(new_n382), .A2(KEYINPUT3), .B1(new_n383), .B2(G104), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n391), .B2(new_n392), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT77), .ZN(new_n399));
  NOR4_X1   g213(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT4), .A4(new_n388), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n215), .B(new_n390), .C1(new_n396), .C2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n197), .B1(new_n403), .B2(new_n207), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n206), .A2(new_n208), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n212), .B2(new_n214), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT78), .B1(new_n383), .B2(G104), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n383), .A2(G104), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n383), .A2(KEYINPUT78), .A3(G104), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n389), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n402), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n413), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n259), .A2(new_n260), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT81), .A4(new_n406), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n401), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n401), .A2(new_n414), .A3(new_n419), .A4(new_n417), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n223), .B(new_n222), .C1(new_n245), .C2(new_n246), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n329), .B1(new_n424), .B2(new_n221), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n247), .A2(new_n249), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n425), .A2(new_n426), .B1(new_n427), .B2(new_n329), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n226), .A2(G125), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT82), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n358), .A2(G224), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT83), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n431), .B(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n418), .A2(new_n435), .A3(new_n420), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n423), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n432), .A2(KEYINPUT7), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n428), .B2(new_n430), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n427), .A2(new_n329), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n226), .A2(new_n426), .A3(G125), .ZN(new_n441));
  AND4_X1   g255(.A1(new_n430), .A2(new_n440), .A3(new_n441), .A4(new_n438), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n422), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n407), .A2(new_n415), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n419), .B(KEYINPUT84), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT8), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n403), .A2(new_n207), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G113), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n206), .A2(KEYINPUT5), .A3(new_n208), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n452), .A2(new_n451), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n453), .A2(new_n454), .B1(new_n260), .B2(new_n259), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n415), .B1(new_n455), .B2(new_n456), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n448), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n444), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n437), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n437), .A2(new_n460), .A3(new_n462), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n378), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n358), .A2(G952), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(G234), .B2(G237), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n303), .B(new_n358), .C1(G234), .C2(G237), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G469), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n255), .B(new_n390), .C1(new_n396), .C2(new_n400), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT10), .B1(new_n413), .B2(new_n427), .ZN(new_n476));
  INV_X1    g290(.A(new_n427), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT10), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n389), .A4(new_n412), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n243), .A2(new_n256), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n475), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT79), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n386), .A2(new_n395), .A3(G101), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n399), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n394), .A2(KEYINPUT77), .A3(new_n395), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n395), .B1(new_n398), .B2(new_n388), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n226), .B1(new_n488), .B2(new_n387), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n487), .A2(new_n489), .B1(new_n476), .B2(new_n479), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT79), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n481), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G110), .B(G140), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n358), .A2(G227), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n481), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n415), .A2(new_n477), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n413), .A2(new_n427), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT12), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT12), .B(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n493), .A2(new_n497), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n490), .A2(new_n481), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n497), .B1(new_n493), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n474), .B(new_n303), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n474), .A2(new_n303), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n491), .B1(new_n490), .B2(new_n481), .ZN(new_n512));
  AND4_X1   g326(.A1(new_n491), .A2(new_n475), .A3(new_n481), .A4(new_n480), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n507), .B(new_n497), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n483), .A2(new_n492), .B1(new_n503), .B2(new_n504), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n514), .B(G469), .C1(new_n515), .C2(new_n497), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n509), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT9), .B(G234), .ZN(new_n518));
  OAI21_X1  g332(.A(G221), .B1(new_n518), .B2(G902), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n518), .A2(new_n366), .A3(G953), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT14), .A4(G122), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT91), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n203), .A2(new_n205), .A3(G122), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT14), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n202), .A2(G122), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n203), .A2(new_n205), .A3(new_n525), .A4(G122), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT91), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n383), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n524), .A2(new_n383), .A3(new_n526), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT90), .B1(new_n218), .B2(G128), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n248), .A3(G143), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT88), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n248), .B2(G143), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n218), .A2(KEYINPUT88), .A3(G128), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(new_n541), .A3(new_n227), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n227), .B1(new_n537), .B2(new_n541), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n533), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT92), .B1(new_n531), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n537), .A2(new_n541), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G134), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n532), .B1(new_n548), .B2(new_n542), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n523), .A2(new_n527), .B1(KEYINPUT91), .B2(new_n529), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(new_n383), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n383), .B1(new_n524), .B2(new_n526), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n542), .B1(new_n532), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n539), .A2(KEYINPUT13), .A3(new_n540), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT13), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n541), .A2(KEYINPUT89), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT89), .B1(new_n541), .B2(new_n557), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n537), .B(new_n556), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n555), .B1(new_n560), .B2(G134), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n520), .B1(new_n553), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n520), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n564), .B(new_n561), .C1(new_n546), .C2(new_n552), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n303), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G478), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(KEYINPUT15), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI221_X1 g383(.A(new_n303), .B1(KEYINPUT15), .B2(new_n567), .C1(new_n563), .C2(new_n565), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n574));
  OAI21_X1  g388(.A(G131), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n576));
  INV_X1    g390(.A(G237), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(new_n358), .A3(G214), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n218), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n239), .A3(new_n572), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n239), .B1(new_n579), .B2(new_n572), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT17), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n581), .A2(new_n352), .A3(new_n335), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(KEYINPUT18), .A2(G131), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n573), .B2(new_n574), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n328), .A2(new_n330), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G146), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n354), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n579), .A2(new_n572), .A3(new_n585), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G113), .B(G122), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(new_n380), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n584), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n595), .B1(new_n584), .B2(new_n593), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n303), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G475), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT19), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n588), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n353), .A2(KEYINPUT19), .ZN(new_n603));
  AOI21_X1  g417(.A(G146), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n340), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n575), .A2(new_n580), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n592), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT87), .B1(new_n607), .B2(new_n595), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT87), .ZN(new_n609));
  INV_X1    g423(.A(new_n595), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n573), .A2(new_n574), .A3(G131), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n582), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n612), .A2(new_n340), .A3(new_n604), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n609), .B(new_n610), .C1(new_n613), .C2(new_n592), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n608), .A2(new_n596), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT20), .ZN(new_n616));
  NOR2_X1   g430(.A1(G475), .A2(G902), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(new_n615), .B2(new_n617), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n600), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n571), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n517), .A2(new_n519), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n473), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n314), .A2(new_n376), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  OAI21_X1  g439(.A(new_n303), .B1(new_n286), .B2(new_n291), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n299), .B1(new_n626), .B2(G472), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n496), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n493), .A2(new_n497), .A3(new_n505), .ZN(new_n630));
  AOI211_X1 g444(.A(G469), .B(G902), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n516), .A2(new_n511), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n519), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n376), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n437), .A2(new_n462), .A3(new_n460), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n462), .B1(new_n437), .B2(new_n460), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n377), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT93), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(KEYINPUT93), .B(new_n377), .C1(new_n637), .C2(new_n638), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n567), .A2(new_n303), .ZN(new_n644));
  INV_X1    g458(.A(new_n566), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(new_n567), .ZN(new_n646));
  OR3_X1    g460(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT33), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT33), .B1(new_n563), .B2(new_n565), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(G478), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n620), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n650), .A2(new_n651), .A3(new_n471), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n636), .A2(new_n643), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G104), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  AND2_X1   g470(.A1(new_n569), .A2(new_n570), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n614), .A2(new_n596), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n602), .A2(new_n603), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n352), .B1(G146), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n593), .B1(new_n660), .B2(new_n612), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n609), .B1(new_n661), .B2(new_n610), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n617), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT20), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(KEYINPUT95), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT95), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n615), .A2(new_n667), .A3(new_n616), .A4(new_n617), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n668), .A2(new_n600), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n657), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n636), .A2(new_n472), .A3(new_n643), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  INV_X1    g488(.A(KEYINPUT96), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n370), .A2(KEYINPUT74), .A3(KEYINPUT25), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT25), .B1(new_n370), .B2(KEYINPUT74), .ZN(new_n677));
  INV_X1    g491(.A(new_n367), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n361), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n356), .B(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n681), .A2(new_n368), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n675), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n375), .A2(KEYINPUT96), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n627), .A2(KEYINPUT97), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(G472), .ZN(new_n688));
  AOI21_X1  g502(.A(G902), .B1(new_n297), .B2(new_n298), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n292), .B(new_n686), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT97), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n687), .A2(new_n692), .A3(new_n623), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT37), .B(G110), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G12));
  INV_X1    g509(.A(G900), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n468), .B1(new_n469), .B2(new_n696), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n657), .A2(new_n670), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n314), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n686), .A2(new_n519), .A3(new_n517), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n641), .B2(new_n642), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  INV_X1    g517(.A(new_n519), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n493), .A2(new_n505), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n496), .B1(new_n483), .B2(new_n492), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n705), .A2(new_n496), .B1(new_n706), .B2(new_n507), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n510), .B1(new_n707), .B2(G469), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n704), .B1(new_n708), .B2(new_n509), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n697), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT98), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT40), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n637), .A2(new_n638), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT38), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n678), .B1(new_n371), .B2(new_n372), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n675), .B(new_n682), .C1(new_n717), .C2(new_n374), .ZN(new_n718));
  AOI21_X1  g532(.A(KEYINPUT96), .B1(new_n375), .B2(new_n684), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n571), .A2(new_n620), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n377), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n295), .A2(new_n313), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n283), .A2(new_n195), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n254), .A2(new_n263), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(G902), .B1(new_n728), .B2(new_n195), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n688), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n299), .B2(KEYINPUT32), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n716), .B(new_n723), .C1(new_n724), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n714), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT99), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT100), .B(G143), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G45));
  AND3_X1   g550(.A1(new_n295), .A2(new_n312), .A3(new_n313), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n633), .A2(new_n720), .ZN(new_n738));
  INV_X1    g552(.A(new_n697), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n646), .A2(new_n649), .A3(new_n620), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n643), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT101), .B1(new_n737), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n700), .A2(new_n740), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT101), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n314), .A2(new_n744), .A3(new_n745), .A4(new_n643), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G146), .ZN(G48));
  AOI22_X1  g562(.A1(new_n628), .A2(new_n496), .B1(new_n706), .B2(new_n505), .ZN(new_n749));
  OAI21_X1  g563(.A(G469), .B1(new_n749), .B2(G902), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n519), .A3(new_n509), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n471), .B(new_n751), .C1(new_n641), .C2(new_n642), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n650), .A2(new_n651), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n314), .A3(new_n376), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(KEYINPUT41), .B(G113), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT102), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n754), .B(new_n756), .ZN(G15));
  NAND4_X1  g571(.A1(new_n752), .A2(new_n314), .A3(new_n376), .A4(new_n671), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G116), .ZN(G18));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n314), .A3(new_n621), .A4(new_n686), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G119), .ZN(G21));
  INV_X1    g575(.A(KEYINPUT104), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT103), .B(G472), .Z(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n626), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n285), .A2(new_n267), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n187), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT104), .B1(new_n689), .B2(new_n763), .ZN(new_n768));
  AND4_X1   g582(.A1(new_n376), .A2(new_n765), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n751), .A2(new_n471), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT105), .B1(new_n643), .B2(new_n722), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT105), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n772), .B(new_n721), .C1(new_n641), .C2(new_n642), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n769), .B(new_n770), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  NAND4_X1  g589(.A1(new_n765), .A2(new_n768), .A3(new_n686), .A4(new_n767), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g591(.A(new_n740), .B(new_n751), .C1(new_n641), .C2(new_n642), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  NAND2_X1  g594(.A1(new_n311), .A2(G472), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n292), .B2(new_n294), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n299), .A2(KEYINPUT32), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n376), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n637), .A2(new_n638), .A3(new_n378), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n741), .A2(new_n709), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT42), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n786), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT42), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n314), .A2(new_n788), .A3(new_n789), .A4(new_n376), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G131), .ZN(G33));
  NAND3_X1  g606(.A1(new_n464), .A2(new_n377), .A3(new_n465), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n633), .A2(new_n634), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n314), .A2(new_n794), .A3(new_n698), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  OR2_X1    g610(.A1(new_n707), .A2(KEYINPUT45), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n707), .A2(KEYINPUT45), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(G469), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT106), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT106), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n511), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(KEYINPUT46), .A3(new_n511), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n509), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n519), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT43), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT107), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n812));
  NAND3_X1  g626(.A1(new_n651), .A2(new_n646), .A3(new_n649), .ZN(new_n813));
  MUX2_X1   g627(.A(new_n811), .B(new_n812), .S(new_n813), .Z(new_n814));
  INV_X1    g628(.A(new_n627), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n686), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT44), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n793), .B1(new_n816), .B2(new_n817), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n809), .A2(new_n710), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G137), .ZN(G39));
  NOR3_X1   g635(.A1(new_n740), .A2(new_n793), .A3(new_n376), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n737), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n807), .A2(KEYINPUT108), .A3(new_n519), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT108), .B1(new_n807), .B2(new_n519), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n824), .B(new_n825), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT108), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n808), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n831), .A2(new_n833), .A3(new_n826), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n823), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(new_n327), .ZN(G42));
  NOR2_X1   g651(.A1(G952), .A2(G953), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT118), .Z(new_n839));
  NOR2_X1   g653(.A1(new_n751), .A2(new_n793), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n468), .A3(new_n814), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n784), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT48), .Z(new_n846));
  NAND3_X1  g660(.A1(new_n769), .A2(new_n468), .A3(new_n814), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n751), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n643), .A3(new_n849), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n467), .B(KEYINPUT117), .Z(new_n851));
  NAND3_X1  g665(.A1(new_n842), .A2(new_n468), .A3(new_n843), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n724), .A2(new_n731), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n852), .A2(new_n634), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n851), .B1(new_n854), .B2(new_n753), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n846), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n750), .A2(new_n704), .A3(new_n509), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n829), .A2(new_n835), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n847), .A2(new_n793), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n620), .B1(new_n646), .B2(new_n649), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n776), .B2(new_n844), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n716), .A2(new_n378), .A3(new_n849), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT113), .Z(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n848), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n867));
  XOR2_X1   g681(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n868));
  AOI211_X1 g682(.A(new_n863), .B(new_n867), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n856), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n860), .A2(KEYINPUT51), .A3(new_n869), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n699), .A2(new_n701), .B1(new_n777), .B2(new_n778), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n633), .A2(new_n679), .A3(new_n682), .A4(new_n697), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n853), .B(new_n879), .C1(new_n771), .C2(new_n773), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n747), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n878), .A2(new_n747), .A3(new_n880), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT110), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n627), .A2(new_n635), .A3(new_n466), .A4(new_n652), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n624), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n624), .B2(new_n887), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n651), .A2(new_n571), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT111), .ZN(new_n892));
  INV_X1    g706(.A(new_n473), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n635), .A3(new_n893), .A4(new_n627), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n693), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n774), .A2(new_n754), .A3(new_n758), .A4(new_n760), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n787), .A2(new_n790), .A3(new_n795), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n569), .A2(new_n570), .A3(new_n739), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n670), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n785), .A2(new_n901), .A3(KEYINPUT112), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT112), .B1(new_n785), .B2(new_n901), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n700), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n314), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n776), .B2(new_n786), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n896), .A2(new_n898), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n877), .B1(new_n885), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n895), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n624), .A2(new_n887), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT110), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n912), .A3(new_n888), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n777), .A2(new_n788), .B1(new_n904), .B2(new_n314), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(new_n787), .A3(new_n790), .A4(new_n795), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n913), .A2(new_n915), .A3(new_n897), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n882), .A3(new_n884), .ZN(new_n917));
  INV_X1    g731(.A(new_n878), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT53), .B1(new_n918), .B2(KEYINPUT52), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n909), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT54), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n877), .B1(new_n918), .B2(KEYINPUT52), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n916), .A2(new_n882), .A3(new_n884), .A4(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n909), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n921), .B(new_n925), .C1(new_n873), .C2(new_n874), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n839), .B1(new_n876), .B2(new_n926), .ZN(new_n927));
  NOR4_X1   g741(.A1(new_n813), .A2(new_n634), .A3(new_n378), .A4(new_n704), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n750), .A2(new_n509), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n929), .A2(KEYINPUT49), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(KEYINPUT49), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n928), .A2(new_n716), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n927), .B1(new_n853), .B2(new_n932), .ZN(G75));
  NOR2_X1   g747(.A1(new_n358), .A2(G952), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n303), .B1(new_n909), .B2(new_n923), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT56), .B1(new_n936), .B2(G210), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n423), .A2(new_n436), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n434), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT55), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n935), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n937), .B2(new_n940), .ZN(G51));
  NAND2_X1  g756(.A1(new_n909), .A2(new_n923), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT54), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n945), .A3(new_n925), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n510), .B(KEYINPUT57), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT120), .ZN(new_n950));
  INV_X1    g764(.A(new_n749), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n946), .A2(new_n952), .A3(new_n947), .A4(new_n948), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n936), .A2(new_n800), .A3(new_n801), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n934), .B1(new_n954), .B2(new_n955), .ZN(G54));
  AND2_X1   g770(.A1(KEYINPUT58), .A2(G475), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n936), .A2(new_n615), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n615), .B1(new_n936), .B2(new_n957), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n934), .ZN(G60));
  XNOR2_X1  g774(.A(new_n644), .B(KEYINPUT59), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n921), .B2(new_n925), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n647), .A2(new_n648), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n647), .B2(new_n648), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n946), .A2(new_n947), .A3(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n964), .A2(KEYINPUT121), .A3(new_n935), .A4(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT121), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n935), .B1(new_n962), .B2(new_n963), .ZN(new_n969));
  INV_X1    g783(.A(new_n966), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n909), .B2(new_n923), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(new_n681), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n365), .B(KEYINPUT122), .Z(new_n977));
  OAI21_X1  g791(.A(new_n935), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT61), .ZN(new_n979));
  OAI22_X1  g793(.A1(new_n976), .A2(new_n978), .B1(KEYINPUT123), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(KEYINPUT123), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT124), .Z(new_n982));
  XOR2_X1   g796(.A(new_n980), .B(new_n982), .Z(G66));
  INV_X1    g797(.A(G224), .ZN(new_n984));
  OAI21_X1  g798(.A(G953), .B1(new_n470), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n913), .A2(new_n897), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n938), .B1(G898), .B2(new_n358), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  NOR2_X1   g803(.A1(new_n696), .A2(new_n358), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n899), .B(KEYINPUT126), .ZN(new_n991));
  INV_X1    g805(.A(new_n771), .ZN(new_n992));
  INV_X1    g806(.A(new_n773), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n784), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n809), .A2(new_n710), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n878), .A2(new_n747), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n820), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n836), .A2(new_n991), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n990), .B1(new_n999), .B2(new_n358), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G227), .A2(G900), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n282), .B(KEYINPUT125), .Z(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(new_n659), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1001), .A2(G953), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1004), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n892), .A2(new_n753), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1007), .A2(new_n793), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1008), .A2(new_n314), .A3(new_n376), .A4(new_n713), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n820), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT99), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n733), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n997), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1010), .B1(new_n1013), .B2(KEYINPUT62), .ZN(new_n1014));
  OR3_X1    g828(.A1(new_n734), .A2(KEYINPUT62), .A3(new_n996), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n358), .B(new_n1006), .C1(new_n1016), .C2(new_n836), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1002), .A2(G953), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1017), .B(new_n1018), .C1(new_n1000), .C2(new_n1006), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n1005), .A2(new_n1019), .ZN(G72));
  AND2_X1   g834(.A1(new_n999), .A2(new_n986), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n283), .B(new_n195), .C1(new_n1021), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n836), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1014), .A2(new_n1026), .A3(new_n1015), .A4(new_n986), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n1023), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n725), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1024), .B1(new_n276), .B2(new_n308), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n934), .B1(new_n920), .B2(new_n1030), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n1025), .A2(new_n1029), .A3(new_n1031), .ZN(G57));
endmodule


