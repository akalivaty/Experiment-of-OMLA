//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n457), .B1(G567), .B2(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT68), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n465), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(new_n469), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n479), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(G137), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n477), .A2(new_n478), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n480), .A2(new_n476), .A3(new_n482), .A4(new_n469), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT70), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n463), .A2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n483), .A2(new_n485), .B1(G101), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n475), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT71), .ZN(G160));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G112), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n480), .A2(new_n469), .A3(new_n476), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT72), .Z(new_n496));
  NAND4_X1  g071(.A1(new_n480), .A2(new_n476), .A3(G2105), .A4(new_n469), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI211_X1 g073(.A(new_n492), .B(new_n496), .C1(G124), .C2(new_n498), .ZN(G162));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n470), .B1(new_n468), .B2(new_n469), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n501), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(G102), .A2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(G2105), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n509), .B(G2104), .C1(G114), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n493), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G126), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n497), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n500), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n467), .A2(new_n471), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT4), .B1(new_n518), .B2(new_n506), .ZN(new_n519));
  NOR3_X1   g094(.A1(new_n501), .A2(new_n505), .A3(G2105), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n520), .A2(new_n469), .A3(new_n480), .A4(new_n476), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n521), .B(new_n511), .C1(new_n514), .C2(new_n497), .ZN(new_n522));
  NOR3_X1   g097(.A1(new_n519), .A2(new_n522), .A3(KEYINPUT73), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(G164));
  OR2_X1    g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n527), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G50), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n527), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G88), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n530), .A2(new_n539), .ZN(G166));
  NAND3_X1  g115(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT74), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n534), .A2(G51), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  INV_X1    g120(.A(G89), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n543), .B(new_n545), .C1(new_n537), .C2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n542), .A2(new_n547), .ZN(G168));
  AOI22_X1  g123(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n529), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n534), .A2(G52), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n537), .B2(new_n552), .ZN(new_n553));
  OR3_X1    g128(.A1(new_n550), .A2(new_n553), .A3(KEYINPUT75), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT75), .B1(new_n550), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(G171));
  AOI22_X1  g131(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n529), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n534), .A2(G43), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n537), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n534), .A2(G53), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT9), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n525), .A2(new_n526), .B1(new_n532), .B2(new_n533), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G91), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n527), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n570), .B(new_n572), .C1(new_n529), .C2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n534), .A2(G49), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n537), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT76), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n583), .B(G651), .C1(new_n527), .C2(G74), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n534), .A2(G48), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n537), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n527), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n529), .ZN(new_n592));
  AND2_X1   g167(.A1(KEYINPUT5), .A2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(KEYINPUT5), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G61), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n597), .A2(KEYINPUT77), .A3(G651), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n589), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G305));
  AOI22_X1  g175(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n529), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n534), .A2(G47), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n537), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G301), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n571), .A2(G92), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT10), .Z(new_n611));
  NAND2_X1  g186(.A1(new_n527), .A2(G66), .ZN(new_n612));
  INV_X1    g187(.A(G79), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n531), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(G54), .B2(new_n534), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n611), .A2(KEYINPUT78), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(KEYINPUT78), .B1(new_n611), .B2(new_n615), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n609), .B1(new_n619), .B2(new_n608), .ZN(G284));
  XOR2_X1   g195(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n608), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n608), .B2(G168), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(new_n608), .B2(G168), .ZN(G280));
  XOR2_X1   g199(.A(KEYINPUT80), .B(G559), .Z(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(G860), .B2(new_n625), .ZN(G148));
  NAND2_X1  g201(.A1(new_n619), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G111), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G2105), .ZN(new_n633));
  AND2_X1   g208(.A1(new_n498), .A2(G123), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT81), .Z(new_n635));
  AOI211_X1 g210(.A(new_n633), .B(new_n635), .C1(G135), .C2(new_n494), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n518), .A2(new_n486), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2100), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n663), .A2(KEYINPUT82), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(KEYINPUT82), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(KEYINPUT17), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n664), .B(new_n665), .C1(new_n660), .C2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n661), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(new_n659), .A3(new_n658), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n660), .A3(new_n658), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(new_n684), .B(new_n683), .S(new_n676), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT84), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT83), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  MUX2_X1   g271(.A(G6), .B(G305), .S(G16), .Z(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT87), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT85), .B(G16), .Z(new_n702));
  MUX2_X1   g277(.A(G303), .B(G22), .S(new_n702), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1971), .ZN(new_n704));
  INV_X1    g279(.A(G23), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G16), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G288), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n704), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n700), .A2(new_n701), .A3(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n714));
  MUX2_X1   g289(.A(G290), .B(G24), .S(new_n702), .Z(new_n715));
  XOR2_X1   g290(.A(KEYINPUT86), .B(G1986), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G25), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n494), .A2(G131), .ZN(new_n720));
  INV_X1    g295(.A(G119), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n510), .A2(G107), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n723));
  OAI22_X1  g298(.A1(new_n497), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n719), .B1(new_n725), .B2(new_n718), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n726), .A2(new_n728), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n717), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n713), .A2(new_n714), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n733));
  OR3_X1    g308(.A1(new_n732), .A2(KEYINPUT88), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT88), .B(KEYINPUT36), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n718), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n718), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT29), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G2090), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G2090), .ZN(new_n741));
  NAND2_X1  g316(.A1(G160), .A2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n743), .B2(KEYINPUT24), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(KEYINPUT24), .B2(new_n743), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G2084), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(G2084), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n740), .A2(new_n741), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G4), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G16), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n618), .B2(G16), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n562), .ZN(new_n755));
  MUX2_X1   g330(.A(new_n755), .B(G19), .S(new_n702), .Z(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT89), .B(G1341), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT90), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n757), .A2(new_n759), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  INV_X1    g337(.A(G28), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n760), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n754), .B(new_n767), .C1(G29), .C2(new_n636), .ZN(new_n768));
  NAND2_X1  g343(.A1(G168), .A2(G16), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(KEYINPUT92), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(KEYINPUT92), .B2(new_n769), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1966), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n718), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  INV_X1    g350(.A(G128), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n510), .A2(G116), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  OAI22_X1  g353(.A1(new_n497), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G140), .B2(new_n494), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(new_n718), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2067), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n752), .B2(new_n753), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n718), .A2(G32), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n494), .A2(G141), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT26), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n788), .A2(new_n789), .B1(G105), .B2(new_n486), .ZN(new_n790));
  INV_X1    g365(.A(G129), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n497), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n785), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n784), .B1(new_n793), .B2(new_n718), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT27), .B(G1996), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT91), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G5), .B(G301), .S(G16), .Z(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G1961), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n718), .A2(G33), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n510), .A2(G103), .A3(G2104), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT25), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n518), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(new_n510), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n802), .B(new_n804), .C1(G139), .C2(new_n494), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n800), .B1(new_n805), .B2(new_n718), .ZN(new_n806));
  AOI211_X1 g381(.A(new_n797), .B(new_n799), .C1(G2072), .C2(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n768), .A2(new_n773), .A3(new_n783), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G164), .A2(new_n718), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G27), .B2(new_n718), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n702), .A2(G20), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT23), .Z(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G299), .B2(G16), .ZN(new_n815));
  INV_X1    g390(.A(G1956), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n798), .B2(G1961), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n810), .A2(new_n811), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n818), .B(new_n819), .C1(G2072), .C2(new_n806), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n749), .A2(new_n808), .A3(new_n812), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n734), .A2(new_n736), .A3(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  NAND2_X1  g398(.A1(new_n619), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n529), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n534), .A2(G55), .ZN(new_n828));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n537), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n562), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n825), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n834));
  AOI21_X1  g409(.A(G860), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT93), .ZN(new_n837));
  OAI21_X1  g412(.A(G860), .B1(new_n827), .B2(new_n830), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  NOR2_X1   g415(.A1(new_n519), .A2(new_n522), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(new_n780), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n793), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n841), .B(new_n780), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n785), .B2(new_n792), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n843), .B(new_n845), .C1(KEYINPUT94), .C2(new_n805), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n805), .A2(KEYINPUT94), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n498), .A2(G130), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n510), .A2(G118), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G142), .B2(new_n494), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n639), .B(new_n853), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n725), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n848), .B(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n636), .B(G160), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G162), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT95), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n856), .A2(new_n858), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(G37), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(KEYINPUT40), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT40), .B1(new_n860), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(G395));
  NAND2_X1  g441(.A1(new_n611), .A2(new_n615), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(G299), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT41), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n832), .B(KEYINPUT96), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n627), .B(new_n871), .ZN(new_n872));
  MUX2_X1   g447(.A(new_n870), .B(new_n868), .S(new_n872), .Z(new_n873));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  XOR2_X1   g451(.A(G166), .B(new_n606), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n599), .B(new_n585), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  OAI21_X1  g456(.A(G868), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(G868), .B2(new_n831), .ZN(G295));
  OAI21_X1  g458(.A(new_n882), .B1(G868), .B2(new_n831), .ZN(G331));
  NAND2_X1  g459(.A1(G171), .A2(KEYINPUT97), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(new_n832), .Z(new_n886));
  OAI21_X1  g461(.A(G286), .B1(G171), .B2(KEYINPUT97), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n889), .A3(new_n868), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n869), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n879), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n897));
  INV_X1    g472(.A(new_n892), .ZN(new_n898));
  INV_X1    g473(.A(new_n879), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n890), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n893), .A2(new_n900), .A3(new_n894), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT99), .B1(new_n902), .B2(KEYINPUT43), .ZN(new_n903));
  OAI211_X1 g478(.A(KEYINPUT98), .B(new_n879), .C1(new_n891), .C2(new_n892), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n879), .A2(KEYINPUT98), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n898), .A2(new_n890), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n894), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n903), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(KEYINPUT101), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(KEYINPUT101), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n904), .A2(new_n906), .A3(new_n897), .A4(new_n894), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT100), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n915), .B2(new_n917), .ZN(G397));
  AOI21_X1  g493(.A(G1384), .B1(new_n508), .B2(new_n516), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n919), .A2(KEYINPUT102), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(KEYINPUT102), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n475), .A2(new_n487), .A3(G40), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n930));
  OR3_X1    g505(.A1(new_n929), .A2(new_n930), .A3(G1996), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n929), .B2(G1996), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n780), .B(G2067), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n933), .A2(new_n793), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n931), .B(new_n932), .C1(new_n929), .C2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n935), .B(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n929), .ZN(new_n938));
  NOR2_X1   g513(.A1(G290), .A2(G1986), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(KEYINPUT48), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n793), .B(G1996), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n728), .B1(new_n720), .B2(new_n724), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n725), .A2(new_n727), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n941), .A2(new_n933), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n940), .B1(new_n929), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT48), .B1(new_n938), .B2(new_n939), .ZN(new_n947));
  AND4_X1   g522(.A1(new_n727), .A2(new_n941), .A3(new_n725), .A4(new_n933), .ZN(new_n948));
  INV_X1    g523(.A(G2067), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(new_n780), .ZN(new_n950));
  OAI22_X1  g525(.A1(new_n946), .A2(new_n947), .B1(new_n929), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n937), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G8), .ZN(new_n953));
  NOR2_X1   g528(.A1(G168), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n519), .B2(new_n522), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n955), .C1(new_n519), .C2(new_n522), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n924), .B1(new_n960), .B2(new_n921), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n508), .A2(new_n516), .A3(new_n500), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT73), .B1(new_n519), .B2(new_n522), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n965));
  AOI21_X1  g540(.A(G1966), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n957), .A2(new_n967), .A3(new_n959), .ZN(new_n968));
  INV_X1    g543(.A(new_n924), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n964), .A2(new_n967), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT115), .B(G2084), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n954), .B1(new_n966), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n976));
  OAI21_X1  g551(.A(G8), .B1(new_n966), .B2(new_n974), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT122), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n954), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n960), .A2(new_n921), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(new_n969), .A3(new_n965), .ZN(new_n981));
  INV_X1    g556(.A(G1966), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n955), .B1(new_n517), .B2(new_n523), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n985), .A2(new_n969), .A3(new_n968), .A4(new_n972), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n953), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT122), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n976), .B1(new_n979), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT123), .ZN(new_n990));
  INV_X1    g565(.A(new_n954), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n976), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n977), .A2(KEYINPUT123), .A3(new_n976), .A4(new_n991), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n975), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n970), .B2(new_n971), .ZN(new_n999));
  INV_X1    g574(.A(G1961), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n985), .A2(KEYINPUT118), .A3(new_n969), .A4(new_n968), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(G2078), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n961), .A2(new_n965), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n924), .B1(KEYINPUT45), .B2(new_n919), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1006), .B(new_n811), .C1(KEYINPUT45), .C2(new_n964), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT124), .B1(new_n1007), .B2(new_n1003), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1007), .A2(KEYINPUT124), .A3(new_n1003), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1002), .B(new_n1005), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT125), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1010), .A2(new_n1011), .A3(G171), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n1010), .B2(G171), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT45), .B(new_n955), .C1(new_n519), .C2(new_n522), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1015), .A2(G40), .A3(new_n475), .A4(new_n487), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n984), .B2(new_n921), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT104), .B1(new_n1017), .B2(G1971), .ZN(new_n1018));
  INV_X1    g593(.A(G2090), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n985), .A2(new_n1019), .A3(new_n969), .A4(new_n968), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1006), .B1(KEYINPUT45), .B2(new_n964), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT104), .ZN(new_n1022));
  INV_X1    g597(.A(G1971), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1018), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G166), .A2(new_n953), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT106), .B(KEYINPUT55), .Z(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  OAI22_X1  g604(.A1(G166), .A2(new_n953), .B1(KEYINPUT106), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1025), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT107), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1025), .A2(KEYINPUT107), .A3(G8), .A4(new_n1031), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n924), .B1(new_n964), .B2(new_n967), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1039), .A2(G2090), .B1(G1971), .B2(new_n1017), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1031), .B1(new_n1040), .B2(G8), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n969), .A2(new_n957), .A3(new_n959), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n1043));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n571), .A2(G86), .B1(new_n534), .B2(G48), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n597), .A2(G651), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n599), .B2(new_n1044), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1043), .B1(new_n1048), .B2(KEYINPUT49), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G1981), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT77), .B1(new_n597), .B2(G651), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n590), .B(new_n529), .C1(new_n595), .C2(new_n596), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1044), .B(new_n1045), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1055), .A2(KEYINPUT111), .A3(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(G8), .B(new_n1042), .C1(new_n1049), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT109), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT49), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1048), .A2(KEYINPUT109), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1062), .A3(new_n1059), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1058), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n582), .A2(new_n584), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  NOR4_X1   g643(.A1(new_n1067), .A2(KEYINPUT108), .A3(new_n1068), .A4(new_n580), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT108), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n585), .B2(G1976), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(G8), .A3(new_n1042), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT52), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1072), .A2(new_n1042), .A3(G8), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT114), .B1(new_n1066), .B2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1042), .A2(G8), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1057), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT111), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1065), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1079), .B(new_n1082), .C1(new_n1083), .C2(new_n1063), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1041), .B1(new_n1078), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1036), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1014), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(new_n975), .C1(new_n989), .C2(new_n995), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n997), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT112), .B1(new_n1066), .B2(new_n1077), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1084), .A2(new_n1094), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1066), .A2(G1976), .A3(G288), .ZN(new_n1098));
  XOR2_X1   g673(.A(new_n1054), .B(KEYINPUT113), .Z(new_n1099));
  OAI21_X1  g674(.A(new_n1079), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n977), .A2(G286), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1036), .A2(new_n1087), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT63), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1025), .A2(G8), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n977), .A2(new_n1104), .A3(G286), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1036), .A2(new_n1107), .A3(new_n1096), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1101), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1092), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1042), .A2(G2067), .ZN(new_n1112));
  XOR2_X1   g687(.A(new_n1112), .B(KEYINPUT117), .Z(new_n1113));
  NAND3_X1  g688(.A1(new_n999), .A2(new_n753), .A3(new_n1001), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(G299), .B(KEYINPUT57), .Z(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1017), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1039), .B2(new_n816), .ZN(new_n1120));
  AOI211_X1 g695(.A(KEYINPUT116), .B(G1956), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1116), .B(new_n1118), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1115), .A2(new_n1122), .A3(new_n619), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1116), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT119), .B(G1996), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1017), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(G1341), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1042), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n755), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT59), .Z(new_n1134));
  NAND3_X1  g709(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n619), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n619), .A2(KEYINPUT60), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n619), .A2(KEYINPUT60), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1113), .A2(new_n1114), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1134), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT61), .B1(new_n1126), .B2(new_n1122), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1126), .A2(KEYINPUT61), .A3(new_n1122), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT121), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1126), .A2(new_n1144), .A3(KEYINPUT61), .A4(new_n1122), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1127), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n1006), .A3(new_n1004), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1002), .B(new_n1148), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G171), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1150), .B(KEYINPUT54), .C1(G171), .C2(new_n1010), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n996), .A2(new_n1036), .A3(new_n1087), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1010), .A2(G171), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT125), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1010), .A2(new_n1011), .A3(G171), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1155), .B(new_n1156), .C1(G171), .C2(new_n1149), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1157), .A2(KEYINPUT126), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT126), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1111), .B1(new_n1153), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n606), .B(G1986), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n929), .B1(new_n945), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n952), .B1(new_n1162), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g740(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n695), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g742(.A(new_n1168), .B1(new_n860), .B2(new_n862), .ZN(new_n1169));
  AND2_X1   g743(.A1(new_n1169), .A2(new_n909), .ZN(G308));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n909), .ZN(G225));
endmodule


