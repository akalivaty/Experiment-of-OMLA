

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U321 ( .A(n368), .B(n367), .ZN(n369) );
  NOR2_X1 U322 ( .A1(n502), .A2(n501), .ZN(n508) );
  XOR2_X1 U323 ( .A(n463), .B(KEYINPUT28), .Z(n528) );
  XOR2_X1 U324 ( .A(G29GAT), .B(G43GAT), .Z(n289) );
  AND2_X1 U325 ( .A1(n562), .A2(n396), .ZN(n397) );
  XNOR2_X1 U326 ( .A(KEYINPUT109), .B(KEYINPUT47), .ZN(n399) );
  INV_X1 U327 ( .A(KEYINPUT118), .ZN(n422) );
  XNOR2_X1 U328 ( .A(n400), .B(n399), .ZN(n406) );
  XNOR2_X1 U329 ( .A(n370), .B(n369), .ZN(n372) );
  XNOR2_X1 U330 ( .A(n422), .B(KEYINPUT54), .ZN(n423) );
  XNOR2_X1 U331 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U332 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U333 ( .A(n380), .B(n379), .ZN(n403) );
  XNOR2_X1 U334 ( .A(n443), .B(n442), .ZN(n444) );
  NOR2_X1 U335 ( .A1(n561), .A2(n530), .ZN(n449) );
  XOR2_X1 U336 ( .A(n420), .B(n419), .Z(n516) );
  INV_X1 U337 ( .A(G190GAT), .ZN(n448) );
  XOR2_X1 U338 ( .A(KEYINPUT11), .B(KEYINPUT73), .Z(n291) );
  XNOR2_X1 U339 ( .A(G50GAT), .B(G190GAT), .ZN(n290) );
  XNOR2_X1 U340 ( .A(n291), .B(n290), .ZN(n298) );
  XOR2_X1 U341 ( .A(G92GAT), .B(KEYINPUT10), .Z(n293) );
  XNOR2_X1 U342 ( .A(KEYINPUT64), .B(KEYINPUT9), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U344 ( .A(n294), .B(KEYINPUT65), .Z(n296) );
  XOR2_X1 U345 ( .A(G134GAT), .B(KEYINPUT74), .Z(n333) );
  XNOR2_X1 U346 ( .A(G218GAT), .B(n333), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n307) );
  XOR2_X1 U349 ( .A(G106GAT), .B(G162GAT), .Z(n300) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U352 ( .A(G99GAT), .B(G85GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n301), .B(KEYINPUT72), .ZN(n384) );
  XOR2_X1 U354 ( .A(n302), .B(n384), .Z(n305) );
  XNOR2_X1 U355 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n289), .B(n303), .ZN(n366) );
  XNOR2_X1 U357 ( .A(G36GAT), .B(n366), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U359 ( .A(n307), .B(n306), .Z(n552) );
  INV_X1 U360 ( .A(n552), .ZN(n537) );
  XOR2_X1 U361 ( .A(KEYINPUT77), .B(G176GAT), .Z(n309) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(KEYINPUT78), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n325) );
  XOR2_X1 U364 ( .A(G120GAT), .B(G99GAT), .Z(n311) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(G134GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U367 ( .A(n312), .B(KEYINPUT79), .Z(n314) );
  XOR2_X1 U368 ( .A(KEYINPUT0), .B(G127GAT), .Z(n332) );
  XNOR2_X1 U369 ( .A(G15GAT), .B(n332), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U371 ( .A(KEYINPUT20), .B(G71GAT), .Z(n316) );
  NAND2_X1 U372 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U374 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U375 ( .A(KEYINPUT18), .B(G190GAT), .Z(n320) );
  XNOR2_X1 U376 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U378 ( .A(KEYINPUT19), .B(n321), .ZN(n418) );
  XOR2_X1 U379 ( .A(G113GAT), .B(n418), .Z(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n465) );
  INV_X1 U382 ( .A(n465), .ZN(n526) );
  XOR2_X1 U383 ( .A(KEYINPUT5), .B(G85GAT), .Z(n327) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(G29GAT), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U386 ( .A(KEYINPUT86), .B(KEYINPUT4), .Z(n329) );
  XNOR2_X1 U387 ( .A(KEYINPUT85), .B(KEYINPUT1), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U389 ( .A(n331), .B(n330), .Z(n338) );
  XOR2_X1 U390 ( .A(G113GAT), .B(G1GAT), .Z(n368) );
  XOR2_X1 U391 ( .A(n333), .B(n332), .Z(n335) );
  NAND2_X1 U392 ( .A1(G225GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n368), .B(n336), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U396 ( .A(n339), .B(KEYINPUT84), .Z(n342) );
  XNOR2_X1 U397 ( .A(G120GAT), .B(G148GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n340), .B(G57GAT), .ZN(n385) );
  XNOR2_X1 U399 ( .A(n385), .B(KEYINPUT6), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n347) );
  XOR2_X1 U401 ( .A(KEYINPUT3), .B(G162GAT), .Z(n344) );
  XNOR2_X1 U402 ( .A(KEYINPUT81), .B(G155GAT), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U404 ( .A(KEYINPUT2), .B(n345), .ZN(n436) );
  INV_X1 U405 ( .A(n436), .ZN(n346) );
  XOR2_X1 U406 ( .A(n347), .B(n346), .Z(n461) );
  XNOR2_X1 U407 ( .A(KEYINPUT87), .B(n461), .ZN(n513) );
  XOR2_X1 U408 ( .A(G64GAT), .B(G57GAT), .Z(n349) );
  XNOR2_X1 U409 ( .A(G1GAT), .B(G211GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n365) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(KEYINPUT70), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n350), .B(KEYINPUT13), .ZN(n383) );
  XOR2_X1 U413 ( .A(n383), .B(KEYINPUT75), .Z(n355) );
  XOR2_X1 U414 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n352) );
  XNOR2_X1 U415 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U417 ( .A(G8GAT), .B(n353), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n363) );
  NAND2_X1 U419 ( .A1(G233GAT), .A2(G231GAT), .ZN(n361) );
  XOR2_X1 U420 ( .A(G78GAT), .B(G155GAT), .Z(n357) );
  XNOR2_X1 U421 ( .A(G22GAT), .B(G15GAT), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n359) );
  XOR2_X1 U423 ( .A(G183GAT), .B(G127GAT), .Z(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U425 ( .A(n361), .B(n360), .Z(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U427 ( .A(n365), .B(n364), .Z(n562) );
  XNOR2_X1 U428 ( .A(n366), .B(KEYINPUT67), .ZN(n370) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U430 ( .A(G15GAT), .B(G197GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n380) );
  XNOR2_X1 U432 ( .A(G50GAT), .B(G22GAT), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n373), .B(G141GAT), .ZN(n437) );
  XNOR2_X1 U434 ( .A(G169GAT), .B(G36GAT), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n374), .B(G8GAT), .ZN(n415) );
  XOR2_X1 U436 ( .A(n437), .B(n415), .Z(n378) );
  XOR2_X1 U437 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n376) );
  XNOR2_X1 U438 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U440 ( .A(G64GAT), .B(G92GAT), .Z(n382) );
  XNOR2_X1 U441 ( .A(G176GAT), .B(G204GAT), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n411) );
  XOR2_X1 U443 ( .A(n411), .B(n383), .Z(n387) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n394) );
  XOR2_X1 U446 ( .A(G106GAT), .B(G78GAT), .Z(n431) );
  XOR2_X1 U447 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n389) );
  XNOR2_X1 U448 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U450 ( .A(n431), .B(n390), .Z(n392) );
  NAND2_X1 U451 ( .A1(G230GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n570) );
  XOR2_X1 U454 ( .A(KEYINPUT41), .B(n570), .Z(n548) );
  NAND2_X1 U455 ( .A1(n403), .A2(n548), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n395), .B(KEYINPUT46), .ZN(n396) );
  XNOR2_X1 U457 ( .A(KEYINPUT108), .B(n397), .ZN(n398) );
  NAND2_X1 U458 ( .A1(n398), .A2(n537), .ZN(n400) );
  XOR2_X1 U459 ( .A(n552), .B(KEYINPUT36), .Z(n580) );
  NOR2_X1 U460 ( .A1(n562), .A2(n580), .ZN(n401) );
  XOR2_X1 U461 ( .A(KEYINPUT45), .B(n401), .Z(n402) );
  NOR2_X1 U462 ( .A1(n570), .A2(n402), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n403), .B(KEYINPUT69), .ZN(n530) );
  NAND2_X1 U464 ( .A1(n404), .A2(n530), .ZN(n405) );
  NAND2_X1 U465 ( .A1(n406), .A2(n405), .ZN(n408) );
  XOR2_X1 U466 ( .A(KEYINPUT110), .B(KEYINPUT48), .Z(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n525) );
  XOR2_X1 U468 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n410) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n412) );
  XOR2_X1 U471 ( .A(n412), .B(n411), .Z(n417) );
  XOR2_X1 U472 ( .A(G211GAT), .B(KEYINPUT21), .Z(n414) );
  XNOR2_X1 U473 ( .A(G197GAT), .B(G218GAT), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n434) );
  XNOR2_X1 U475 ( .A(n415), .B(n434), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n420) );
  INV_X1 U477 ( .A(n418), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n516), .B(KEYINPUT117), .ZN(n421) );
  NOR2_X1 U479 ( .A1(n525), .A2(n421), .ZN(n424) );
  NOR2_X1 U480 ( .A1(n513), .A2(n425), .ZN(n566) );
  XOR2_X1 U481 ( .A(G204GAT), .B(KEYINPUT22), .Z(n427) );
  XNOR2_X1 U482 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n441) );
  XOR2_X1 U484 ( .A(G148GAT), .B(KEYINPUT83), .Z(n429) );
  XNOR2_X1 U485 ( .A(KEYINPUT80), .B(KEYINPUT82), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U487 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U490 ( .A(n435), .B(n434), .Z(n439) );
  XOR2_X1 U491 ( .A(n437), .B(n436), .Z(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U493 ( .A(n441), .B(n440), .Z(n463) );
  NAND2_X1 U494 ( .A1(n566), .A2(n463), .ZN(n443) );
  XOR2_X1 U495 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n442) );
  NAND2_X1 U496 ( .A1(n526), .A2(n444), .ZN(n561) );
  NOR2_X1 U497 ( .A1(n537), .A2(n561), .ZN(n446) );
  XNOR2_X1 U498 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  INV_X1 U501 ( .A(G169GAT), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n449), .B(KEYINPUT120), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(G1348GAT) );
  XOR2_X1 U504 ( .A(KEYINPUT93), .B(KEYINPUT34), .Z(n472) );
  NOR2_X1 U505 ( .A1(n530), .A2(n570), .ZN(n487) );
  INV_X1 U506 ( .A(n487), .ZN(n470) );
  NOR2_X1 U507 ( .A1(n552), .A2(n562), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n452), .B(KEYINPUT16), .ZN(n469) );
  NAND2_X1 U509 ( .A1(n516), .A2(n526), .ZN(n453) );
  NAND2_X1 U510 ( .A1(n453), .A2(n463), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n454), .B(KEYINPUT91), .ZN(n455) );
  XNOR2_X1 U512 ( .A(KEYINPUT25), .B(n455), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n463), .A2(n526), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT26), .ZN(n565) );
  XNOR2_X1 U515 ( .A(n516), .B(KEYINPUT27), .ZN(n464) );
  NAND2_X1 U516 ( .A1(n565), .A2(n464), .ZN(n457) );
  XNOR2_X1 U517 ( .A(KEYINPUT90), .B(n457), .ZN(n458) );
  NAND2_X1 U518 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U519 ( .A(KEYINPUT92), .B(n460), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n462), .A2(n461), .ZN(n468) );
  NAND2_X1 U521 ( .A1(n513), .A2(n464), .ZN(n524) );
  NOR2_X1 U522 ( .A1(n528), .A2(n524), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n484) );
  NAND2_X1 U525 ( .A1(n469), .A2(n484), .ZN(n501) );
  NOR2_X1 U526 ( .A1(n470), .A2(n501), .ZN(n480) );
  NAND2_X1 U527 ( .A1(n480), .A2(n513), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  NAND2_X1 U530 ( .A1(n480), .A2(n516), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(KEYINPUT94), .ZN(n475) );
  XNOR2_X1 U532 ( .A(G8GAT), .B(n475), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT35), .B(KEYINPUT96), .Z(n477) );
  NAND2_X1 U534 ( .A1(n480), .A2(n526), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n479) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT95), .Z(n478) );
  XNOR2_X1 U537 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n482) );
  NAND2_X1 U539 ( .A1(n480), .A2(n528), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U541 ( .A(G22GAT), .B(n483), .ZN(G1327GAT) );
  INV_X1 U542 ( .A(n562), .ZN(n574) );
  NOR2_X1 U543 ( .A1(n574), .A2(n580), .ZN(n485) );
  NAND2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(n486), .ZN(n512) );
  NAND2_X1 U546 ( .A1(n487), .A2(n512), .ZN(n488) );
  XOR2_X1 U547 ( .A(KEYINPUT38), .B(n488), .Z(n499) );
  NAND2_X1 U548 ( .A1(n499), .A2(n513), .ZN(n493) );
  XOR2_X1 U549 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n490) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(KEYINPUT99), .B(n491), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n495) );
  NAND2_X1 U555 ( .A1(n516), .A2(n499), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n499), .A2(n526), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U561 ( .A1(n499), .A2(n528), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U563 ( .A(n548), .ZN(n555) );
  NOR2_X1 U564 ( .A1(n403), .A2(n555), .ZN(n511) );
  INV_X1 U565 ( .A(n511), .ZN(n502) );
  NAND2_X1 U566 ( .A1(n513), .A2(n508), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n516), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n508), .A2(n526), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U575 ( .A1(n508), .A2(n528), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  XOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT105), .Z(n515) );
  AND2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n520) );
  NAND2_X1 U579 ( .A1(n520), .A2(n513), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n520), .A2(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n526), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT106), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n522) );
  NAND2_X1 U587 ( .A1(n520), .A2(n528), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n543) );
  NAND2_X1 U591 ( .A1(n526), .A2(n543), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(KEYINPUT111), .B(n529), .ZN(n538) );
  NOR2_X1 U594 ( .A1(n530), .A2(n538), .ZN(n531) );
  XOR2_X1 U595 ( .A(G113GAT), .B(n531), .Z(G1340GAT) );
  NOR2_X1 U596 ( .A1(n555), .A2(n538), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n562), .A2(n538), .ZN(n535) );
  XNOR2_X1 U600 ( .A(KEYINPUT112), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U602 ( .A(G127GAT), .B(n536), .Z(G1342GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n542) );
  XOR2_X1 U604 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n540) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  AND2_X1 U608 ( .A1(n543), .A2(n565), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n403), .A2(n553), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(KEYINPUT115), .B(n547), .Z(n550) );
  NAND2_X1 U615 ( .A1(n553), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n553), .A2(n574), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n561), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(KEYINPUT56), .B(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n579) );
  INV_X1 U631 ( .A(n579), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n575), .A2(n403), .ZN(n569) );
  XOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .Z(n567) );
  XNOR2_X1 U634 ( .A(KEYINPUT59), .B(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U637 ( .A1(n575), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(n582), .B(n581), .Z(G1355GAT) );
endmodule

