

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(G651), .A2(n625), .ZN(n646) );
  NOR2_X4 U550 ( .A1(G2105), .A2(G2104), .ZN(n555) );
  INV_X1 U551 ( .A(KEYINPUT17), .ZN(n554) );
  AND2_X1 U552 ( .A1(n557), .A2(n556), .ZN(G164) );
  AND2_X2 U553 ( .A1(n552), .A2(G2104), .ZN(n893) );
  NOR2_X2 U554 ( .A1(G543), .A2(G651), .ZN(n642) );
  INV_X1 U555 ( .A(G651), .ZN(n523) );
  XNOR2_X1 U556 ( .A(n705), .B(KEYINPUT28), .ZN(n712) );
  INV_X1 U557 ( .A(KEYINPUT96), .ZN(n715) );
  NOR2_X2 U558 ( .A1(n625), .A2(n523), .ZN(n643) );
  NOR2_X1 U559 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U560 ( .A1(G543), .A2(n523), .ZN(n516) );
  XOR2_X1 U561 ( .A(n715), .B(KEYINPUT29), .Z(n513) );
  AND2_X1 U562 ( .A1(n551), .A2(n550), .ZN(n514) );
  INV_X1 U563 ( .A(KEYINPUT94), .ZN(n692) );
  BUF_X1 U564 ( .A(n701), .Z(n717) );
  INV_X1 U565 ( .A(KEYINPUT97), .ZN(n722) );
  INV_X1 U566 ( .A(KEYINPUT99), .ZN(n739) );
  XNOR2_X1 U567 ( .A(KEYINPUT100), .B(KEYINPUT32), .ZN(n742) );
  INV_X1 U568 ( .A(n779), .ZN(n757) );
  INV_X1 U569 ( .A(n968), .ZN(n764) );
  INV_X1 U570 ( .A(KEYINPUT1), .ZN(n515) );
  AND2_X2 U571 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NOR2_X1 U572 ( .A1(n539), .A2(n538), .ZN(G171) );
  XNOR2_X2 U573 ( .A(n516), .B(n515), .ZN(n650) );
  NAND2_X1 U574 ( .A1(n650), .A2(G63), .ZN(n517) );
  XNOR2_X1 U575 ( .A(n517), .B(KEYINPUT72), .ZN(n519) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n625) );
  NAND2_X1 U577 ( .A1(G51), .A2(n646), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U579 ( .A(KEYINPUT6), .B(n520), .ZN(n529) );
  NAND2_X1 U580 ( .A1(G89), .A2(n642), .ZN(n521) );
  XNOR2_X1 U581 ( .A(n521), .B(KEYINPUT70), .ZN(n522) );
  XNOR2_X1 U582 ( .A(n522), .B(KEYINPUT4), .ZN(n525) );
  NAND2_X1 U583 ( .A1(G76), .A2(n643), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U585 ( .A(KEYINPUT71), .B(n526), .ZN(n527) );
  XNOR2_X1 U586 ( .A(KEYINPUT5), .B(n527), .ZN(n528) );
  NOR2_X1 U587 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U588 ( .A(KEYINPUT7), .B(n530), .Z(G168) );
  XNOR2_X1 U589 ( .A(G168), .B(KEYINPUT8), .ZN(n531) );
  XNOR2_X1 U590 ( .A(n531), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U591 ( .A1(G90), .A2(n642), .ZN(n533) );
  NAND2_X1 U592 ( .A1(G77), .A2(n643), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U594 ( .A(n534), .B(KEYINPUT9), .ZN(n536) );
  NAND2_X1 U595 ( .A1(G52), .A2(n646), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n539) );
  NAND2_X1 U597 ( .A1(G64), .A2(n650), .ZN(n537) );
  XNOR2_X1 U598 ( .A(KEYINPUT65), .B(n537), .ZN(n538) );
  XOR2_X1 U599 ( .A(G2438), .B(G2454), .Z(n541) );
  XNOR2_X1 U600 ( .A(G2435), .B(G2430), .ZN(n540) );
  XNOR2_X1 U601 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U602 ( .A(n542), .B(G2427), .Z(n544) );
  XNOR2_X1 U603 ( .A(G1341), .B(G1348), .ZN(n543) );
  XNOR2_X1 U604 ( .A(n544), .B(n543), .ZN(n548) );
  XOR2_X1 U605 ( .A(G2443), .B(G2446), .Z(n546) );
  XNOR2_X1 U606 ( .A(KEYINPUT106), .B(G2451), .ZN(n545) );
  XNOR2_X1 U607 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U608 ( .A(n548), .B(n547), .Z(n549) );
  AND2_X1 U609 ( .A1(G14), .A2(n549), .ZN(G401) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U611 ( .A1(G114), .A2(n897), .ZN(n551) );
  NOR2_X1 U612 ( .A1(n552), .A2(G2104), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G126), .A2(n558), .ZN(n550) );
  INV_X1 U614 ( .A(G2105), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G102), .A2(n893), .ZN(n553) );
  AND2_X1 U616 ( .A1(n514), .A2(n553), .ZN(n557) );
  XNOR2_X2 U617 ( .A(n555), .B(n554), .ZN(n892) );
  NAND2_X1 U618 ( .A1(n892), .A2(G138), .ZN(n556) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  INV_X1 U621 ( .A(G120), .ZN(G236) );
  INV_X1 U622 ( .A(G69), .ZN(G235) );
  BUF_X1 U623 ( .A(n558), .Z(n896) );
  NAND2_X1 U624 ( .A1(n896), .A2(G125), .ZN(n561) );
  NAND2_X1 U625 ( .A1(G101), .A2(n893), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT23), .B(n559), .Z(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n685) );
  NAND2_X1 U628 ( .A1(n892), .A2(G137), .ZN(n563) );
  NAND2_X1 U629 ( .A1(G113), .A2(n897), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n683) );
  NOR2_X1 U631 ( .A1(n685), .A2(n683), .ZN(G160) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n837) );
  NAND2_X1 U635 ( .A1(n837), .A2(G567), .ZN(n565) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U637 ( .A1(G81), .A2(n642), .ZN(n566) );
  XNOR2_X1 U638 ( .A(n566), .B(KEYINPUT12), .ZN(n567) );
  XNOR2_X1 U639 ( .A(n567), .B(KEYINPUT66), .ZN(n569) );
  NAND2_X1 U640 ( .A1(G68), .A2(n643), .ZN(n568) );
  NAND2_X1 U641 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U642 ( .A(n570), .B(KEYINPUT13), .ZN(n572) );
  NAND2_X1 U643 ( .A1(G43), .A2(n646), .ZN(n571) );
  NAND2_X1 U644 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n650), .A2(G56), .ZN(n573) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(n573), .Z(n574) );
  NOR2_X2 U647 ( .A1(n575), .A2(n574), .ZN(n971) );
  NAND2_X1 U648 ( .A1(n971), .A2(G860), .ZN(G153) );
  XNOR2_X1 U649 ( .A(G171), .B(KEYINPUT67), .ZN(G301) );
  NAND2_X1 U650 ( .A1(n646), .A2(G54), .ZN(n582) );
  NAND2_X1 U651 ( .A1(G92), .A2(n642), .ZN(n577) );
  NAND2_X1 U652 ( .A1(G79), .A2(n643), .ZN(n576) );
  NAND2_X1 U653 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U654 ( .A1(n650), .A2(G66), .ZN(n578) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(n578), .Z(n579) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U657 ( .A(KEYINPUT15), .B(n583), .Z(n974) );
  INV_X1 U658 ( .A(n974), .ZN(n617) );
  NOR2_X1 U659 ( .A1(n617), .A2(G868), .ZN(n584) );
  XNOR2_X1 U660 ( .A(n584), .B(KEYINPUT69), .ZN(n586) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U662 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G53), .A2(n646), .ZN(n588) );
  NAND2_X1 U664 ( .A1(G65), .A2(n650), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G91), .A2(n642), .ZN(n590) );
  NAND2_X1 U667 ( .A1(G78), .A2(n643), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n977) );
  INV_X1 U670 ( .A(n977), .ZN(G299) );
  NOR2_X1 U671 ( .A1(G868), .A2(G299), .ZN(n594) );
  INV_X1 U672 ( .A(G868), .ZN(n662) );
  NOR2_X1 U673 ( .A1(G286), .A2(n662), .ZN(n593) );
  NOR2_X1 U674 ( .A1(n594), .A2(n593), .ZN(G297) );
  INV_X1 U675 ( .A(G860), .ZN(n619) );
  NAND2_X1 U676 ( .A1(n619), .A2(G559), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n595), .A2(n617), .ZN(n596) );
  XNOR2_X1 U678 ( .A(n596), .B(KEYINPUT16), .ZN(n597) );
  XNOR2_X1 U679 ( .A(KEYINPUT74), .B(n597), .ZN(G148) );
  NAND2_X1 U680 ( .A1(n617), .A2(G868), .ZN(n598) );
  NOR2_X1 U681 ( .A1(G559), .A2(n598), .ZN(n600) );
  AND2_X1 U682 ( .A1(n662), .A2(n971), .ZN(n599) );
  NOR2_X1 U683 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G123), .A2(n896), .ZN(n601) );
  XNOR2_X1 U685 ( .A(n601), .B(KEYINPUT18), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n893), .A2(G99), .ZN(n602) );
  NAND2_X1 U687 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U688 ( .A1(G135), .A2(n892), .ZN(n605) );
  NAND2_X1 U689 ( .A1(G111), .A2(n897), .ZN(n604) );
  NAND2_X1 U690 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n1007) );
  XNOR2_X1 U692 ( .A(G2096), .B(n1007), .ZN(n609) );
  INV_X1 U693 ( .A(G2100), .ZN(n608) );
  NAND2_X1 U694 ( .A1(n609), .A2(n608), .ZN(G156) );
  NAND2_X1 U695 ( .A1(G55), .A2(n646), .ZN(n611) );
  NAND2_X1 U696 ( .A1(G67), .A2(n650), .ZN(n610) );
  NAND2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n616) );
  NAND2_X1 U698 ( .A1(G93), .A2(n642), .ZN(n613) );
  NAND2_X1 U699 ( .A1(G80), .A2(n643), .ZN(n612) );
  NAND2_X1 U700 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U701 ( .A(KEYINPUT75), .B(n614), .Z(n615) );
  OR2_X1 U702 ( .A1(n616), .A2(n615), .ZN(n661) );
  XNOR2_X1 U703 ( .A(n661), .B(KEYINPUT76), .ZN(n621) );
  NAND2_X1 U704 ( .A1(G559), .A2(n617), .ZN(n618) );
  XNOR2_X1 U705 ( .A(n618), .B(n971), .ZN(n658) );
  NAND2_X1 U706 ( .A1(n658), .A2(n619), .ZN(n620) );
  XNOR2_X1 U707 ( .A(n621), .B(n620), .ZN(G145) );
  NAND2_X1 U708 ( .A1(G49), .A2(n646), .ZN(n623) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n622) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U711 ( .A1(n650), .A2(n624), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n625), .A2(G87), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G48), .A2(n646), .ZN(n629) );
  NAND2_X1 U715 ( .A1(G86), .A2(n642), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n643), .A2(G73), .ZN(n630) );
  XOR2_X1 U718 ( .A(KEYINPUT2), .B(n630), .Z(n631) );
  NOR2_X1 U719 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U720 ( .A1(n650), .A2(G61), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G88), .A2(n642), .ZN(n636) );
  NAND2_X1 U723 ( .A1(G75), .A2(n643), .ZN(n635) );
  NAND2_X1 U724 ( .A1(n636), .A2(n635), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G62), .A2(n650), .ZN(n637) );
  XOR2_X1 U726 ( .A(KEYINPUT77), .B(n637), .Z(n639) );
  NAND2_X1 U727 ( .A1(n646), .A2(G50), .ZN(n638) );
  NAND2_X1 U728 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U729 ( .A1(n641), .A2(n640), .ZN(G166) );
  NAND2_X1 U730 ( .A1(G85), .A2(n642), .ZN(n645) );
  NAND2_X1 U731 ( .A1(G72), .A2(n643), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U733 ( .A1(G47), .A2(n646), .ZN(n647) );
  XOR2_X1 U734 ( .A(KEYINPUT64), .B(n647), .Z(n648) );
  NOR2_X1 U735 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n650), .A2(G60), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(G290) );
  XNOR2_X1 U738 ( .A(KEYINPUT19), .B(G288), .ZN(n657) );
  XNOR2_X1 U739 ( .A(G166), .B(n661), .ZN(n653) );
  XNOR2_X1 U740 ( .A(G305), .B(n653), .ZN(n654) );
  XNOR2_X1 U741 ( .A(n977), .B(n654), .ZN(n655) );
  XNOR2_X1 U742 ( .A(n655), .B(G290), .ZN(n656) );
  XNOR2_X1 U743 ( .A(n657), .B(n656), .ZN(n864) );
  XNOR2_X1 U744 ( .A(n864), .B(n658), .ZN(n659) );
  NAND2_X1 U745 ( .A1(n659), .A2(G868), .ZN(n660) );
  XNOR2_X1 U746 ( .A(n660), .B(KEYINPUT78), .ZN(n664) );
  NAND2_X1 U747 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XNOR2_X1 U750 ( .A(n665), .B(KEYINPUT20), .ZN(n666) );
  XNOR2_X1 U751 ( .A(n666), .B(KEYINPUT79), .ZN(n667) );
  NAND2_X1 U752 ( .A1(n667), .A2(G2090), .ZN(n668) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U756 ( .A1(G235), .A2(G236), .ZN(n670) );
  XNOR2_X1 U757 ( .A(KEYINPUT80), .B(n670), .ZN(n671) );
  NAND2_X1 U758 ( .A1(n671), .A2(G57), .ZN(n672) );
  XNOR2_X1 U759 ( .A(KEYINPUT81), .B(n672), .ZN(n673) );
  NAND2_X1 U760 ( .A1(n673), .A2(G108), .ZN(n842) );
  NAND2_X1 U761 ( .A1(G567), .A2(n842), .ZN(n678) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U764 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U765 ( .A1(G96), .A2(n676), .ZN(n843) );
  NAND2_X1 U766 ( .A1(G2106), .A2(n843), .ZN(n677) );
  NAND2_X1 U767 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U768 ( .A(KEYINPUT82), .B(n679), .Z(G319) );
  INV_X1 U769 ( .A(G319), .ZN(n913) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n680) );
  XOR2_X1 U771 ( .A(KEYINPUT83), .B(n680), .Z(n681) );
  NOR2_X1 U772 ( .A1(n913), .A2(n681), .ZN(n839) );
  NAND2_X1 U773 ( .A1(n839), .A2(G36), .ZN(G176) );
  XOR2_X1 U774 ( .A(KEYINPUT84), .B(G166), .Z(G303) );
  INV_X1 U775 ( .A(G40), .ZN(n682) );
  OR2_X2 U776 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U777 ( .A1(n685), .A2(n684), .ZN(n783) );
  NOR2_X2 U778 ( .A1(G164), .A2(G1384), .ZN(n785) );
  AND2_X2 U779 ( .A1(n783), .A2(n785), .ZN(n701) );
  NAND2_X1 U780 ( .A1(n701), .A2(G1996), .ZN(n687) );
  XNOR2_X1 U781 ( .A(n687), .B(KEYINPUT26), .ZN(n689) );
  INV_X1 U782 ( .A(n701), .ZN(n733) );
  NAND2_X1 U783 ( .A1(G1341), .A2(n733), .ZN(n688) );
  NAND2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U785 ( .A(n690), .B(KEYINPUT93), .ZN(n691) );
  NAND2_X1 U786 ( .A1(n691), .A2(n971), .ZN(n699) );
  NOR2_X2 U787 ( .A1(n699), .A2(n974), .ZN(n693) );
  XNOR2_X1 U788 ( .A(n693), .B(n692), .ZN(n698) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n733), .ZN(n695) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n717), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U792 ( .A(KEYINPUT95), .B(n696), .Z(n697) );
  NAND2_X1 U793 ( .A1(n698), .A2(n697), .ZN(n709) );
  BUF_X1 U794 ( .A(n699), .Z(n700) );
  NAND2_X1 U795 ( .A1(n700), .A2(n974), .ZN(n707) );
  NAND2_X1 U796 ( .A1(n701), .A2(G2072), .ZN(n702) );
  XNOR2_X1 U797 ( .A(n702), .B(KEYINPUT27), .ZN(n704) );
  XOR2_X1 U798 ( .A(KEYINPUT92), .B(G1956), .Z(n948) );
  NOR2_X1 U799 ( .A1(n717), .A2(n948), .ZN(n703) );
  NOR2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n710) );
  NOR2_X1 U801 ( .A1(n977), .A2(n710), .ZN(n705) );
  INV_X1 U802 ( .A(n712), .ZN(n706) );
  AND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n977), .A2(n710), .ZN(n711) );
  OR2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n716) );
  XNOR2_X1 U808 ( .A(n716), .B(n513), .ZN(n721) );
  INV_X1 U809 ( .A(G1961), .ZN(n961) );
  NAND2_X1 U810 ( .A1(n733), .A2(n961), .ZN(n719) );
  XNOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .ZN(n928) );
  NAND2_X1 U812 ( .A1(n717), .A2(n928), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n724) );
  NAND2_X1 U814 ( .A1(G171), .A2(n724), .ZN(n720) );
  NAND2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U816 ( .A(n723), .B(n722), .ZN(n732) );
  NOR2_X1 U817 ( .A1(G171), .A2(n724), .ZN(n729) );
  NAND2_X1 U818 ( .A1(G8), .A2(n733), .ZN(n779) );
  NOR2_X1 U819 ( .A1(G1966), .A2(n779), .ZN(n747) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n733), .ZN(n749) );
  NOR2_X1 U821 ( .A1(n747), .A2(n749), .ZN(n725) );
  NAND2_X1 U822 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U824 ( .A1(G168), .A2(n727), .ZN(n728) );
  NOR2_X1 U825 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U826 ( .A(KEYINPUT31), .B(n730), .Z(n731) );
  NAND2_X1 U827 ( .A1(n732), .A2(n731), .ZN(n744) );
  NAND2_X1 U828 ( .A1(n744), .A2(G286), .ZN(n738) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n779), .ZN(n735) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U831 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U832 ( .A1(G303), .A2(n736), .ZN(n737) );
  NAND2_X1 U833 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U834 ( .A(n740), .B(n739), .ZN(n741) );
  NAND2_X1 U835 ( .A1(n741), .A2(G8), .ZN(n743) );
  XNOR2_X1 U836 ( .A(n743), .B(n742), .ZN(n753) );
  BUF_X1 U837 ( .A(n744), .Z(n745) );
  INV_X1 U838 ( .A(n745), .ZN(n746) );
  NOR2_X1 U839 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U840 ( .A(n748), .B(KEYINPUT98), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n749), .A2(G8), .ZN(n750) );
  NAND2_X1 U842 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n768) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n761) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U846 ( .A1(n761), .A2(n754), .ZN(n981) );
  NAND2_X1 U847 ( .A1(n768), .A2(n981), .ZN(n755) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n980) );
  NAND2_X1 U849 ( .A1(n755), .A2(n980), .ZN(n756) );
  XNOR2_X1 U850 ( .A(n756), .B(KEYINPUT101), .ZN(n758) );
  NAND2_X1 U851 ( .A1(n758), .A2(n757), .ZN(n760) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U853 ( .A1(n760), .A2(n759), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n761), .A2(KEYINPUT33), .ZN(n762) );
  NOR2_X1 U855 ( .A1(n762), .A2(n779), .ZN(n765) );
  XOR2_X1 U856 ( .A(G1981), .B(KEYINPUT102), .Z(n763) );
  XNOR2_X1 U857 ( .A(G305), .B(n763), .ZN(n968) );
  NOR2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U859 ( .A1(n767), .A2(n766), .ZN(n775) );
  BUF_X1 U860 ( .A(n768), .Z(n771) );
  NOR2_X1 U861 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U862 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n779), .A2(n772), .ZN(n773) );
  XOR2_X1 U865 ( .A(KEYINPUT103), .B(n773), .Z(n774) );
  NAND2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U867 ( .A(n776), .B(KEYINPUT104), .ZN(n781) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U869 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  NOR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X2 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U872 ( .A(n782), .B(KEYINPUT105), .ZN(n821) );
  INV_X1 U873 ( .A(n783), .ZN(n784) );
  NOR2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n832) );
  NAND2_X1 U875 ( .A1(G117), .A2(n897), .ZN(n786) );
  XOR2_X1 U876 ( .A(KEYINPUT88), .B(n786), .Z(n789) );
  NAND2_X1 U877 ( .A1(n893), .A2(G105), .ZN(n787) );
  XOR2_X1 U878 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n896), .A2(G129), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n792), .B(KEYINPUT89), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G141), .A2(n892), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n876) );
  NAND2_X1 U885 ( .A1(G1996), .A2(n876), .ZN(n803) );
  NAND2_X1 U886 ( .A1(G131), .A2(n892), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G95), .A2(n893), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G119), .A2(n896), .ZN(n797) );
  XNOR2_X1 U890 ( .A(KEYINPUT87), .B(n797), .ZN(n798) );
  NOR2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n897), .A2(G107), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n886) );
  NAND2_X1 U894 ( .A1(G1991), .A2(n886), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U896 ( .A(KEYINPUT90), .B(n804), .Z(n1017) );
  INV_X1 U897 ( .A(n1017), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n832), .A2(n805), .ZN(n822) );
  NAND2_X1 U899 ( .A1(G140), .A2(n892), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G104), .A2(n893), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U902 ( .A(KEYINPUT34), .B(n808), .ZN(n813) );
  NAND2_X1 U903 ( .A1(G128), .A2(n896), .ZN(n810) );
  NAND2_X1 U904 ( .A1(G116), .A2(n897), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U906 ( .A(KEYINPUT35), .B(n811), .Z(n812) );
  NOR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U908 ( .A(KEYINPUT36), .B(n814), .ZN(n907) );
  XNOR2_X1 U909 ( .A(KEYINPUT37), .B(G2067), .ZN(n830) );
  NOR2_X1 U910 ( .A1(n907), .A2(n830), .ZN(n999) );
  NAND2_X1 U911 ( .A1(n832), .A2(n999), .ZN(n828) );
  NAND2_X1 U912 ( .A1(n822), .A2(n828), .ZN(n815) );
  XNOR2_X1 U913 ( .A(n815), .B(KEYINPUT91), .ZN(n819) );
  XOR2_X1 U914 ( .A(G1986), .B(KEYINPUT85), .Z(n816) );
  XNOR2_X1 U915 ( .A(G290), .B(n816), .ZN(n976) );
  NAND2_X1 U916 ( .A1(n976), .A2(n832), .ZN(n817) );
  XNOR2_X1 U917 ( .A(KEYINPUT86), .B(n817), .ZN(n818) );
  AND2_X1 U918 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n821), .A2(n820), .ZN(n835) );
  NOR2_X1 U920 ( .A1(G1996), .A2(n876), .ZN(n1015) );
  INV_X1 U921 ( .A(n822), .ZN(n825) );
  NOR2_X1 U922 ( .A1(G1991), .A2(n886), .ZN(n1008) );
  NOR2_X1 U923 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U924 ( .A1(n1008), .A2(n823), .ZN(n824) );
  NOR2_X1 U925 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U926 ( .A1(n1015), .A2(n826), .ZN(n827) );
  XNOR2_X1 U927 ( .A(n827), .B(KEYINPUT39), .ZN(n829) );
  NAND2_X1 U928 ( .A1(n829), .A2(n828), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n907), .A2(n830), .ZN(n998) );
  NAND2_X1 U930 ( .A1(n831), .A2(n998), .ZN(n833) );
  NAND2_X1 U931 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U932 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U936 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U938 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U939 ( .A(KEYINPUT107), .B(n841), .Z(G188) );
  XNOR2_X1 U940 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G57), .ZN(G237) );
  NOR2_X1 U944 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XOR2_X1 U946 ( .A(KEYINPUT110), .B(G1971), .Z(n845) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1976), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U949 ( .A(n846), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U952 ( .A(G1966), .B(G1956), .Z(n850) );
  XNOR2_X1 U953 ( .A(G1981), .B(G1961), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U955 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U956 ( .A(KEYINPUT109), .B(G2474), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(G229) );
  XOR2_X1 U958 ( .A(G2096), .B(KEYINPUT43), .Z(n856) );
  XNOR2_X1 U959 ( .A(G2072), .B(KEYINPUT108), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U961 ( .A(n857), .B(G2678), .Z(n859) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2090), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U964 ( .A(KEYINPUT42), .B(G2100), .Z(n861) );
  XNOR2_X1 U965 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n863), .B(n862), .ZN(G227) );
  XOR2_X1 U968 ( .A(n864), .B(n971), .Z(n866) );
  XNOR2_X1 U969 ( .A(G286), .B(G171), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(n974), .B(n867), .Z(n868) );
  NOR2_X1 U972 ( .A1(G37), .A2(n868), .ZN(G397) );
  NAND2_X1 U973 ( .A1(G124), .A2(n896), .ZN(n869) );
  XNOR2_X1 U974 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n893), .A2(G100), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G136), .A2(n892), .ZN(n873) );
  NAND2_X1 U978 ( .A1(G112), .A2(n897), .ZN(n872) );
  NAND2_X1 U979 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U980 ( .A1(n875), .A2(n874), .ZN(G162) );
  XNOR2_X1 U981 ( .A(G160), .B(n876), .ZN(n889) );
  NAND2_X1 U982 ( .A1(G118), .A2(n897), .ZN(n885) );
  NAND2_X1 U983 ( .A1(n896), .A2(G130), .ZN(n877) );
  XNOR2_X1 U984 ( .A(KEYINPUT111), .B(n877), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G142), .A2(n892), .ZN(n879) );
  NAND2_X1 U986 ( .A1(G106), .A2(n893), .ZN(n878) );
  NAND2_X1 U987 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U988 ( .A(KEYINPUT112), .B(n880), .Z(n881) );
  XNOR2_X1 U989 ( .A(KEYINPUT45), .B(n881), .ZN(n882) );
  NOR2_X1 U990 ( .A1(n883), .A2(n882), .ZN(n884) );
  NAND2_X1 U991 ( .A1(n885), .A2(n884), .ZN(n887) );
  XNOR2_X1 U992 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U993 ( .A(n889), .B(n888), .ZN(n909) );
  XOR2_X1 U994 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n891) );
  XNOR2_X1 U995 ( .A(G164), .B(KEYINPUT113), .ZN(n890) );
  XNOR2_X1 U996 ( .A(n891), .B(n890), .ZN(n903) );
  NAND2_X1 U997 ( .A1(G139), .A2(n892), .ZN(n895) );
  NAND2_X1 U998 ( .A1(G103), .A2(n893), .ZN(n894) );
  NAND2_X1 U999 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(G127), .A2(n896), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(G115), .A2(n897), .ZN(n898) );
  NAND2_X1 U1002 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1003 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(n1001) );
  XOR2_X1 U1005 ( .A(n903), .B(n1001), .Z(n905) );
  XNOR2_X1 U1006 ( .A(G162), .B(n1007), .ZN(n904) );
  XNOR2_X1 U1007 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n910), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n911) );
  XNOR2_X1 U1013 ( .A(n912), .B(n911), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(n913), .A2(G401), .ZN(n914) );
  XOR2_X1 U1015 ( .A(KEYINPUT114), .B(n914), .Z(n915) );
  NOR2_X1 U1016 ( .A1(G397), .A2(n915), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n918), .A2(G395), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n919), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1020 ( .A(G308), .ZN(G225) );
  XNOR2_X1 U1021 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n1022) );
  XNOR2_X1 U1022 ( .A(G1991), .B(G25), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(G33), .B(G2072), .ZN(n920) );
  NOR2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n927) );
  XOR2_X1 U1025 ( .A(G1996), .B(G32), .Z(n922) );
  NAND2_X1 U1026 ( .A1(n922), .A2(G28), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(KEYINPUT120), .B(G2067), .ZN(n923) );
  XNOR2_X1 U1028 ( .A(G26), .B(n923), .ZN(n924) );
  NOR2_X1 U1029 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1031 ( .A(G27), .B(n928), .Z(n929) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1033 ( .A(KEYINPUT53), .B(n931), .Z(n934) );
  XOR2_X1 U1034 ( .A(KEYINPUT54), .B(G34), .Z(n932) );
  XNOR2_X1 U1035 ( .A(G2084), .B(n932), .ZN(n933) );
  NAND2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(G35), .B(G2090), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1039 ( .A(n1022), .B(n937), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(G29), .A2(n938), .ZN(n939) );
  XOR2_X1 U1041 ( .A(KEYINPUT121), .B(n939), .Z(n995) );
  XNOR2_X1 U1042 ( .A(G1986), .B(G24), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(G1976), .B(G23), .ZN(n941) );
  XNOR2_X1 U1044 ( .A(G1971), .B(G22), .ZN(n940) );
  NOR2_X1 U1045 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1046 ( .A(KEYINPUT125), .B(n942), .ZN(n943) );
  NOR2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1048 ( .A(KEYINPUT58), .B(n945), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(KEYINPUT123), .B(G1341), .ZN(n946) );
  XNOR2_X1 U1050 ( .A(n946), .B(G19), .ZN(n952) );
  XOR2_X1 U1051 ( .A(G1348), .B(KEYINPUT59), .Z(n947) );
  XNOR2_X1 U1052 ( .A(G4), .B(n947), .ZN(n950) );
  XOR2_X1 U1053 ( .A(n948), .B(G20), .Z(n949) );
  NOR2_X1 U1054 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1055 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1056 ( .A(KEYINPUT124), .B(G1981), .ZN(n953) );
  XNOR2_X1 U1057 ( .A(G6), .B(n953), .ZN(n954) );
  NOR2_X1 U1058 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1059 ( .A(KEYINPUT60), .B(n956), .Z(n958) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G21), .ZN(n957) );
  NOR2_X1 U1061 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1062 ( .A1(n960), .A2(n959), .ZN(n964) );
  XOR2_X1 U1063 ( .A(KEYINPUT122), .B(n961), .Z(n962) );
  XNOR2_X1 U1064 ( .A(G5), .B(n962), .ZN(n963) );
  NOR2_X1 U1065 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1066 ( .A(KEYINPUT61), .B(n965), .Z(n966) );
  NOR2_X1 U1067 ( .A1(G16), .A2(n966), .ZN(n967) );
  XOR2_X1 U1068 ( .A(KEYINPUT126), .B(n967), .Z(n993) );
  XNOR2_X1 U1069 ( .A(KEYINPUT56), .B(G16), .ZN(n991) );
  XNOR2_X1 U1070 ( .A(G168), .B(G1966), .ZN(n969) );
  NAND2_X1 U1071 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1072 ( .A(n970), .B(KEYINPUT57), .ZN(n989) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n971), .ZN(n973) );
  NAND2_X1 U1074 ( .A1(G303), .A2(G1971), .ZN(n972) );
  NAND2_X1 U1075 ( .A1(n973), .A2(n972), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(n974), .B(G1348), .ZN(n975) );
  NOR2_X1 U1077 ( .A1(n976), .A2(n975), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n977), .B(G1956), .ZN(n979) );
  XNOR2_X1 U1079 ( .A(G171), .B(G1961), .ZN(n978) );
  NAND2_X1 U1080 ( .A1(n979), .A2(n978), .ZN(n983) );
  NAND2_X1 U1081 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1082 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1083 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1085 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(G11), .A2(n996), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(n997), .B(KEYINPUT127), .ZN(n1026) );
  INV_X1 U1091 ( .A(n998), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1013) );
  XOR2_X1 U1093 ( .A(G2072), .B(n1001), .Z(n1003) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(G160), .B(G2084), .ZN(n1005) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1100 ( .A(KEYINPUT118), .B(n1009), .Z(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1105 ( .A(KEYINPUT51), .B(n1016), .Z(n1018) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(G29), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

