//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT14), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n204), .A2(KEYINPUT90), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(KEYINPUT90), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n205), .A2(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n208), .B(new_n209), .C1(new_n204), .C2(KEYINPUT90), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(KEYINPUT91), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n208), .B2(new_n209), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT91), .B1(new_n207), .B2(new_n210), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n203), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT92), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n203), .B1(new_n207), .B2(new_n210), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n216), .B(new_n217), .C1(new_n208), .C2(new_n209), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT93), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n214), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT17), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(new_n214), .C1(new_n220), .C2(new_n221), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT7), .ZN(new_n228));
  INV_X1    g027(.A(G99gat), .ZN(new_n229));
  INV_X1    g028(.A(G106gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT8), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n228), .B(new_n231), .C1(G85gat), .C2(G92gat), .ZN(new_n232));
  XOR2_X1   g031(.A(G99gat), .B(G106gat), .Z(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n234), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n240));
  OR2_X1    g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n240), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G190gat), .B(G218gat), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G134gat), .B(G162gat), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n242), .A3(new_n248), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G15gat), .B(G22gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT16), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(G1gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(G1gat), .B2(new_n254), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(G8gat), .Z(new_n258));
  NAND2_X1  g057(.A1(G71gat), .A2(G78gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT96), .ZN(new_n260));
  INV_X1    g059(.A(G71gat), .ZN(new_n261));
  INV_X1    g060(.A(G78gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G57gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G64gat), .ZN(new_n265));
  INV_X1    g064(.A(G64gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G57gat), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n259), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n260), .B(new_n263), .C1(new_n268), .C2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n267), .B(KEYINPUT98), .Z(new_n272));
  XOR2_X1   g071(.A(new_n265), .B(KEYINPUT97), .Z(new_n273));
  OAI22_X1  g072(.A1(new_n272), .A2(new_n273), .B1(KEYINPUT9), .B2(new_n269), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n263), .A2(new_n259), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n275), .B(KEYINPUT99), .Z(new_n276));
  OAI21_X1  g075(.A(new_n271), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n258), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G183gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n278), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n285), .ZN(new_n287));
  XOR2_X1   g086(.A(KEYINPUT101), .B(G211gat), .Z(new_n288));
  NAND2_X1  g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G127gat), .B(G155gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT100), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n290), .B(new_n292), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n286), .A2(new_n287), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n286), .B2(new_n287), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G230gat), .A2(G233gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n277), .B(new_n234), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n277), .A2(new_n234), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n298), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G120gat), .B(G148gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(G176gat), .B(G204gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT104), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT104), .ZN(new_n312));
  NOR4_X1   g111(.A1(new_n303), .A2(new_n312), .A3(new_n305), .A4(new_n309), .ZN(new_n313));
  OAI22_X1  g112(.A1(new_n311), .A2(new_n313), .B1(new_n306), .B2(new_n310), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n253), .A2(new_n296), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(G50gat), .ZN(new_n318));
  XOR2_X1   g117(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G22gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT83), .ZN(new_n323));
  XOR2_X1   g122(.A(G197gat), .B(G204gat), .Z(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n326));
  INV_X1    g125(.A(G218gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(KEYINPUT71), .A2(G218gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(G211gat), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT22), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n330), .A2(KEYINPUT72), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT72), .B1(new_n330), .B2(new_n331), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n325), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n338));
  AND2_X1   g137(.A1(KEYINPUT71), .A2(G218gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(KEYINPUT71), .A2(G218gat), .ZN(new_n340));
  INV_X1    g139(.A(G211gat), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n338), .B1(new_n342), .B2(KEYINPUT22), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n330), .A2(KEYINPUT72), .A3(new_n331), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(new_n325), .A3(new_n335), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G155gat), .ZN(new_n348));
  INV_X1    g147(.A(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(G141gat), .B(G148gat), .Z(new_n353));
  INV_X1    g152(.A(KEYINPUT2), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n351), .B1(new_n350), .B2(KEYINPUT2), .ZN(new_n356));
  INV_X1    g155(.A(G148gat), .ZN(new_n357));
  OR2_X1    g156(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G141gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(G148gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n356), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT78), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n365), .B(new_n356), .C1(new_n360), .C2(new_n362), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n355), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n347), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n335), .B1(new_n345), .B2(new_n325), .ZN(new_n373));
  AOI211_X1 g172(.A(new_n324), .B(new_n336), .C1(new_n343), .C2(new_n344), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT82), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n347), .A2(new_n377), .A3(new_n371), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n368), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n355), .ZN(new_n380));
  INV_X1    g179(.A(new_n366), .ZN(new_n381));
  AND2_X1   g180(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n383));
  OAI21_X1  g182(.A(G148gat), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n362), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n365), .B1(new_n386), .B2(new_n356), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n380), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n372), .B1(new_n379), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n323), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT3), .B1(new_n375), .B2(KEYINPUT82), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n367), .B1(new_n393), .B2(new_n378), .ZN(new_n394));
  OAI211_X1 g193(.A(KEYINPUT83), .B(new_n390), .C1(new_n394), .C2(new_n372), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n337), .B2(new_n346), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n397), .B2(KEYINPUT84), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n373), .A2(new_n374), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(KEYINPUT29), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n367), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n402), .A2(new_n390), .A3(new_n372), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n322), .B1(new_n396), .B2(new_n404), .ZN(new_n405));
  AOI211_X1 g204(.A(G22gat), .B(new_n403), .C1(new_n392), .C2(new_n395), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n321), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n370), .B1(new_n337), .B2(new_n346), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n368), .B1(new_n408), .B2(new_n377), .ZN(new_n409));
  AOI211_X1 g208(.A(KEYINPUT82), .B(new_n370), .C1(new_n337), .C2(new_n346), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n388), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n372), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT83), .B1(new_n413), .B2(new_n390), .ZN(new_n414));
  AOI211_X1 g213(.A(new_n323), .B(new_n391), .C1(new_n411), .C2(new_n412), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n404), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G22gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n396), .A2(new_n322), .A3(new_n404), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(new_n320), .ZN(new_n419));
  XOR2_X1   g218(.A(G15gat), .B(G43gat), .Z(new_n420));
  XOR2_X1   g219(.A(G71gat), .B(G99gat), .Z(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G183gat), .A2(G190gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT24), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n426));
  INV_X1    g225(.A(G190gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n280), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT25), .B1(new_n429), .B2(KEYINPUT64), .ZN(new_n430));
  AND2_X1   g229(.A1(G169gat), .A2(G176gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(KEYINPUT23), .B2(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n432), .A2(KEYINPUT23), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(new_n435), .ZN(new_n437));
  AND2_X1   g236(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n427), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT28), .ZN(new_n441));
  NAND2_X1  g240(.A1(G169gat), .A2(G176gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT26), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n432), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT65), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT28), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n446), .B(new_n427), .C1(new_n438), .C2(new_n439), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n441), .A2(new_n445), .A3(new_n423), .A4(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NOR3_X1   g248(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n444), .A2(KEYINPUT65), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n436), .A2(new_n437), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454));
  INV_X1    g253(.A(G113gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(G120gat), .ZN(new_n456));
  INV_X1    g255(.A(G120gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(G113gat), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n454), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT1), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(G113gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(G120gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT67), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT66), .B(G127gat), .Z(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G134gat), .ZN(new_n466));
  OR2_X1    g265(.A1(G127gat), .A2(G134gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G127gat), .B(G134gat), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n469), .B(new_n460), .C1(new_n456), .C2(new_n458), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n430), .A2(new_n435), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n430), .A2(new_n435), .ZN(new_n475));
  OAI22_X1  g274(.A1(new_n474), .A2(new_n475), .B1(new_n451), .B2(new_n448), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n471), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(G227gat), .A2(G233gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n481));
  INV_X1    g280(.A(KEYINPUT32), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n422), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n473), .B2(new_n477), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n422), .A2(KEYINPUT69), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n422), .A2(KEYINPUT69), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n486), .A2(new_n482), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT34), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n485), .A3(new_n477), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n480), .A2(KEYINPUT32), .A3(new_n489), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n496));
  INV_X1    g295(.A(new_n422), .ZN(new_n497));
  INV_X1    g296(.A(new_n483), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n486), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n492), .A2(new_n494), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n494), .B1(new_n492), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n407), .A2(new_n419), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G8gat), .B(G36gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(G64gat), .B(G92gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G226gat), .ZN(new_n508));
  INV_X1    g307(.A(G233gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT29), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n476), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n510), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n430), .B(new_n435), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n449), .A2(new_n452), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n347), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n476), .A2(new_n510), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n370), .B1(new_n514), .B2(new_n515), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n518), .B(new_n400), .C1(new_n519), .C2(new_n510), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n507), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT74), .B1(new_n521), .B2(KEYINPUT30), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(new_n520), .ZN(new_n525));
  INV_X1    g324(.A(new_n507), .ZN(new_n526));
  OAI22_X1  g325(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT75), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n525), .B2(new_n526), .ZN(new_n530));
  AOI211_X1 g329(.A(KEYINPUT75), .B(new_n507), .C1(new_n517), .C2(new_n520), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT76), .B(new_n528), .C1(new_n530), .C2(new_n531), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n527), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n388), .B(new_n471), .ZN(new_n537));
  NAND2_X1  g336(.A1(G225gat), .A2(G233gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(new_n369), .A3(new_n471), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT79), .B(KEYINPUT4), .C1(new_n388), .C2(new_n471), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT4), .B1(new_n388), .B2(new_n471), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n367), .A2(new_n546), .A3(new_n468), .A4(new_n470), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT79), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(KEYINPUT5), .B(new_n540), .C1(new_n544), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n547), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n539), .A2(KEYINPUT5), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n542), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G57gat), .B(G85gat), .Z(new_n555));
  XNOR2_X1  g354(.A(G1gat), .B(G29gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n561));
  INV_X1    g360(.A(new_n559), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n550), .A2(new_n562), .A3(new_n553), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n554), .A2(KEYINPUT6), .A3(new_n559), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n536), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT35), .B1(new_n504), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT89), .ZN(new_n569));
  INV_X1    g368(.A(new_n504), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT35), .B1(new_n567), .B2(KEYINPUT88), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n534), .A2(new_n535), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n525), .A2(new_n526), .ZN(new_n573));
  INV_X1    g372(.A(new_n524), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n522), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n572), .A2(new_n566), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT88), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n570), .A2(new_n571), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n580), .B(KEYINPUT35), .C1(new_n504), .C2(new_n567), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n569), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n513), .B1(new_n453), .B2(KEYINPUT29), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n400), .B1(new_n583), .B2(new_n518), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n510), .B1(new_n476), .B2(new_n371), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n585), .A2(new_n516), .A3(new_n347), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n526), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT75), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n521), .A2(new_n529), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT76), .B1(new_n590), .B2(new_n528), .ZN(new_n591));
  INV_X1    g390(.A(new_n535), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n575), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n538), .B1(new_n551), .B2(new_n542), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n595), .B(KEYINPUT39), .C1(new_n539), .C2(new_n537), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT85), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT40), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n559), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n598), .B1(new_n596), .B2(new_n600), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n593), .A2(new_n603), .A3(new_n560), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT86), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n407), .A2(new_n419), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n526), .B1(new_n525), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n608), .B1(new_n607), .B2(new_n525), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n609), .A2(KEYINPUT87), .A3(KEYINPUT38), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT87), .B1(new_n609), .B2(KEYINPUT38), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n566), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n583), .A2(new_n518), .A3(new_n400), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n347), .B1(new_n585), .B2(new_n516), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n616), .A3(KEYINPUT37), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n608), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n612), .A2(new_n613), .A3(new_n590), .A4(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT86), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n593), .A2(new_n603), .A3(new_n620), .A4(new_n560), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n619), .A4(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT70), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(new_n501), .B2(new_n502), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT36), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n623), .B(KEYINPUT36), .C1(new_n501), .C2(new_n502), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n407), .A2(new_n419), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n567), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n582), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G113gat), .B(G141gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G197gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT11), .B(G169gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n226), .A2(new_n258), .ZN(new_n638));
  INV_X1    g437(.A(new_n258), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n222), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G229gat), .A2(G233gat), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n638), .A2(KEYINPUT18), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n640), .B1(new_n226), .B2(new_n258), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n646), .A2(KEYINPUT94), .A3(KEYINPUT18), .A4(new_n642), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n642), .ZN(new_n649));
  AOI211_X1 g448(.A(new_n649), .B(new_n640), .C1(new_n226), .C2(new_n258), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n222), .B(new_n258), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n642), .B(KEYINPUT13), .ZN(new_n652));
  OAI22_X1  g451(.A1(new_n650), .A2(KEYINPUT18), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n637), .B1(new_n648), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n646), .A2(new_n642), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT18), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n637), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n658), .A2(new_n645), .A3(new_n647), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n632), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT95), .ZN(new_n663));
  INV_X1    g462(.A(new_n661), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n582), .B2(new_n631), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n316), .B1(new_n663), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n613), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n593), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT16), .B(G8gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(G8gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n673), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n668), .A2(KEYINPUT42), .A3(new_n593), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1325gat));
  AOI21_X1  g479(.A(G15gat), .B1(new_n668), .B2(new_n503), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n628), .A2(G15gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT106), .Z(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n668), .B2(new_n683), .ZN(G1326gat));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n629), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  NAND2_X1  g486(.A1(new_n663), .A2(new_n667), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n296), .A2(new_n314), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n252), .A3(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(G29gat), .A3(new_n566), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT45), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  AOI211_X1 g493(.A(new_n694), .B(new_n253), .C1(new_n582), .C2(new_n631), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n622), .A2(KEYINPUT107), .A3(new_n630), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT107), .B1(new_n622), .B2(new_n630), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n582), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n252), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n695), .B1(new_n699), .B2(new_n694), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n661), .A3(new_n689), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(new_n566), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n693), .B1(new_n702), .B2(G29gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n692), .B1(new_n703), .B2(new_n691), .ZN(G1328gat));
  NOR3_X1   g503(.A1(new_n690), .A2(G36gat), .A3(new_n536), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G36gat), .B1(new_n701), .B2(new_n536), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(G1329gat));
  INV_X1    g509(.A(new_n628), .ZN(new_n711));
  OAI21_X1  g510(.A(G43gat), .B1(new_n701), .B2(new_n711), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n296), .B(new_n314), .C1(new_n663), .C2(new_n667), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n503), .A3(new_n252), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n714), .B2(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1330gat));
  OAI21_X1  g516(.A(G50gat), .B1(new_n701), .B2(new_n606), .ZN(new_n718));
  INV_X1    g517(.A(G50gat), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n713), .A2(new_n719), .A3(new_n629), .A4(new_n252), .ZN(new_n720));
  OR2_X1    g519(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1331gat));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n631), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n622), .A2(new_n630), .A3(KEYINPUT107), .ZN(new_n727));
  INV_X1    g526(.A(new_n581), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n576), .A2(new_n503), .A3(new_n419), .A4(new_n407), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n580), .B1(new_n729), .B2(KEYINPUT35), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n726), .A2(new_n727), .B1(new_n731), .B2(new_n579), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n661), .ZN(new_n733));
  INV_X1    g532(.A(new_n296), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(new_n252), .A3(new_n315), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n566), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n264), .ZN(G1332gat));
  INV_X1    g537(.A(new_n736), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n536), .B(KEYINPUT109), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n266), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT110), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n266), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1333gat));
  NAND3_X1  g545(.A1(new_n733), .A2(new_n503), .A3(new_n735), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n733), .A2(KEYINPUT111), .A3(new_n503), .A4(new_n735), .ZN(new_n750));
  AOI21_X1  g549(.A(G71gat), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n261), .B1(new_n739), .B2(new_n628), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g553(.A1(new_n736), .A2(new_n606), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n262), .ZN(G1335gat));
  OAI21_X1  g555(.A(new_n694), .B1(new_n732), .B2(new_n253), .ZN(new_n757));
  INV_X1    g556(.A(new_n695), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n661), .A2(new_n296), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n757), .A2(new_n314), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(G85gat), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n760), .A2(new_n761), .A3(new_n566), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n698), .A2(new_n252), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT51), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n698), .A2(new_n759), .A3(new_n765), .A4(new_n252), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n613), .A3(new_n314), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n762), .B1(new_n769), .B2(new_n761), .ZN(G1336gat));
  NAND4_X1  g569(.A1(new_n700), .A2(new_n593), .A3(new_n314), .A4(new_n759), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n771), .A2(new_n772), .A3(G92gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n764), .A2(new_n766), .B1(KEYINPUT113), .B2(new_n763), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n763), .A2(KEYINPUT113), .A3(new_n765), .ZN(new_n775));
  INV_X1    g574(.A(new_n740), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(G92gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n314), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n774), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n772), .B1(new_n771), .B2(G92gat), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n773), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n700), .A2(new_n314), .A3(new_n740), .A4(new_n759), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(new_n783), .B2(G92gat), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n764), .A2(new_n314), .A3(new_n766), .A4(new_n777), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT114), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G92gat), .B1(new_n760), .B2(new_n776), .ZN(new_n787));
  AND4_X1   g586(.A1(KEYINPUT114), .A2(new_n787), .A3(new_n782), .A4(new_n785), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n781), .A2(new_n782), .B1(new_n786), .B2(new_n788), .ZN(G1337gat));
  NAND4_X1  g588(.A1(new_n768), .A2(new_n229), .A3(new_n503), .A4(new_n314), .ZN(new_n790));
  OAI21_X1  g589(.A(G99gat), .B1(new_n760), .B2(new_n711), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1338gat));
  NOR2_X1   g591(.A1(new_n760), .A2(new_n606), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n230), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n629), .A2(new_n230), .A3(new_n314), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n774), .A2(new_n775), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n767), .B2(new_n795), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n799), .B2(new_n794), .ZN(G1339gat));
  INV_X1    g599(.A(new_n313), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n300), .A2(new_n302), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n297), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n304), .A3(new_n310), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n312), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n300), .A2(new_n302), .A3(new_n298), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n310), .B1(new_n303), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(KEYINPUT55), .A3(new_n810), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n806), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n654), .B2(new_n660), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n646), .A2(new_n642), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n651), .A2(new_n652), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n636), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n660), .A2(new_n314), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n253), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n660), .A2(new_n819), .ZN(new_n823));
  INV_X1    g622(.A(new_n815), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n252), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n296), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n316), .A2(new_n661), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(new_n613), .A3(new_n570), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n776), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n664), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(new_n455), .ZN(G1340gat));
  NOR2_X1   g631(.A1(new_n830), .A2(new_n315), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(new_n457), .ZN(G1341gat));
  NOR2_X1   g633(.A1(new_n830), .A2(new_n734), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n465), .A2(KEYINPUT115), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n835), .B(new_n836), .ZN(G1342gat));
  OAI21_X1  g636(.A(G134gat), .B1(new_n830), .B2(new_n253), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT117), .ZN(new_n839));
  INV_X1    g638(.A(G134gat), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n253), .A2(new_n593), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n829), .A2(new_n840), .A3(new_n841), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n839), .A2(new_n846), .ZN(G1343gat));
  NOR2_X1   g646(.A1(new_n628), .A2(new_n566), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n828), .A2(new_n629), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n664), .A2(G141gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n776), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT119), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n828), .A2(new_n854), .A3(new_n629), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n776), .A2(new_n848), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n316), .A2(new_n661), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n823), .A2(new_n252), .A3(new_n824), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n661), .A2(new_n824), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n820), .A2(KEYINPUT118), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n660), .A2(new_n862), .A3(new_n314), .A4(new_n819), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n859), .B1(new_n864), .B2(new_n253), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n858), .B1(new_n865), .B2(new_n296), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n854), .B1(new_n866), .B2(new_n629), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n856), .A2(new_n857), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n661), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n382), .A2(new_n383), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n853), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n849), .B(KEYINPUT120), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n776), .A3(new_n850), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n872), .ZN(new_n876));
  OAI22_X1  g675(.A1(new_n871), .A2(new_n872), .B1(new_n873), .B2(new_n876), .ZN(G1344gat));
  AND2_X1   g676(.A1(new_n874), .A2(new_n776), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n357), .A3(new_n314), .ZN(new_n879));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n357), .C1(new_n868), .C2(new_n314), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  INV_X1    g680(.A(new_n857), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n866), .B2(new_n629), .ZN(new_n883));
  OAI211_X1 g682(.A(KEYINPUT57), .B(new_n629), .C1(new_n826), .C2(new_n827), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n314), .B(new_n882), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n881), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n879), .B1(new_n880), .B2(new_n887), .ZN(G1345gat));
  INV_X1    g687(.A(new_n868), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(new_n348), .A3(new_n734), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n878), .A2(new_n296), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n348), .ZN(G1346gat));
  OAI21_X1  g691(.A(G162gat), .B1(new_n889), .B2(new_n253), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n874), .A2(new_n349), .A3(new_n841), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1347gat));
  OAI21_X1  g694(.A(new_n566), .B1(new_n826), .B2(new_n827), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n504), .A2(new_n536), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G169gat), .B1(new_n899), .B2(new_n664), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n901), .A2(new_n740), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n570), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n905), .A2(G169gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n900), .B1(new_n906), .B2(new_n664), .ZN(G1348gat));
  INV_X1    g706(.A(new_n905), .ZN(new_n908));
  AOI21_X1  g707(.A(G176gat), .B1(new_n908), .B2(new_n314), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n899), .A2(new_n315), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(G176gat), .B2(new_n910), .ZN(G1349gat));
  OAI21_X1  g710(.A(G183gat), .B1(new_n899), .B2(new_n734), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n296), .B1(new_n439), .B2(new_n438), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n913), .B1(new_n908), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(KEYINPUT123), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT123), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n920), .B(new_n912), .C1(new_n905), .C2(new_n914), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n916), .A2(new_n918), .B1(new_n921), .B2(new_n917), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n899), .B2(new_n253), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n252), .A2(new_n427), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n905), .B2(new_n925), .ZN(G1351gat));
  NOR2_X1   g725(.A1(new_n606), .A2(new_n628), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n901), .A2(new_n740), .A3(new_n903), .A4(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(G197gat), .A3(new_n664), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT124), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n536), .A2(new_n613), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n711), .B(new_n931), .C1(new_n883), .C2(new_n885), .ZN(new_n932));
  OAI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n664), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(new_n933), .ZN(G1352gat));
  NOR3_X1   g733(.A1(new_n928), .A2(G204gat), .A3(new_n315), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT62), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n932), .A2(KEYINPUT125), .A3(new_n315), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT125), .B1(new_n932), .B2(new_n315), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(G204gat), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(G1353gat));
  NAND2_X1  g739(.A1(new_n866), .A2(new_n629), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n854), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n628), .B1(new_n942), .B2(new_n884), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n943), .A2(KEYINPUT126), .A3(new_n296), .A4(new_n931), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n932), .B2(new_n734), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n946), .A3(G211gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n948));
  NOR2_X1   g747(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n944), .A2(new_n946), .A3(G211gat), .A4(new_n949), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n904), .A2(new_n341), .A3(new_n296), .A4(new_n927), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(G1354gat));
  NOR4_X1   g753(.A1(new_n932), .A2(new_n340), .A3(new_n339), .A4(new_n253), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n904), .A2(new_n252), .A3(new_n927), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n327), .B2(new_n956), .ZN(G1355gat));
endmodule


