//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n627, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT65), .Z(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(G137), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n467), .A2(new_n463), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n458), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n459), .A2(new_n461), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(new_n463), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  NAND2_X1  g056(.A1(new_n462), .A2(new_n463), .ZN(new_n482));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT4), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n474), .A2(new_n485), .A3(G138), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n463), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n476), .A2(G126), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  AND2_X1   g068(.A1(KEYINPUT6), .A2(G651), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT6), .A2(G651), .ZN(new_n495));
  OAI21_X1  g070(.A(G543), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G50), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n498), .A2(KEYINPUT67), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(KEYINPUT67), .ZN(new_n500));
  INV_X1    g075(.A(new_n495), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n501), .A2(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n499), .A2(new_n500), .B1(G88), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT68), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n510), .B2(KEYINPUT68), .ZN(new_n514));
  OAI21_X1  g089(.A(G651), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n508), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n509), .A2(new_n518), .A3(G89), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n522), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n519), .A2(KEYINPUT70), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(KEYINPUT70), .B1(new_n519), .B2(new_n524), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n518), .B2(G543), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n528), .B(G543), .C1(new_n494), .C2(new_n495), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(G51), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n509), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n527), .A2(new_n535), .ZN(G168));
  NAND3_X1  g111(.A1(new_n509), .A2(new_n518), .A3(G90), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G651), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n496), .A2(KEYINPUT69), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n541), .B1(new_n542), .B2(new_n530), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n539), .ZN(new_n546));
  OAI21_X1  g121(.A(G43), .B1(new_n529), .B2(new_n531), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n509), .A2(new_n518), .A3(G81), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n542), .B2(new_n530), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT71), .B1(new_n553), .B2(new_n549), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n546), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  AND2_X1   g137(.A1(KEYINPUT5), .A2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(KEYINPUT5), .A2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n497), .A2(KEYINPUT9), .A3(G53), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n507), .A2(G91), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n496), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n573), .ZN(G299));
  OAI21_X1  g149(.A(KEYINPUT72), .B1(new_n540), .B2(new_n543), .ZN(new_n575));
  NAND2_X1  g150(.A1(G77), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G64), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n565), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n507), .B2(G90), .ZN(new_n579));
  OAI21_X1  g154(.A(G52), .B1(new_n529), .B2(new_n531), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G301));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n527), .B2(new_n535), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n542), .A2(new_n530), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G51), .B1(new_n509), .B2(new_n533), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n588), .B(KEYINPUT73), .C1(new_n526), .C2(new_n525), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G286));
  NAND2_X1  g166(.A1(new_n497), .A2(G49), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n507), .A2(G87), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  AOI22_X1  g170(.A1(G48), .A2(new_n497), .B1(new_n507), .B2(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n509), .A2(G61), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n597), .A2(new_n598), .B1(G73), .B2(G543), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n509), .A2(KEYINPUT74), .A3(G61), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n596), .B1(new_n601), .B2(new_n539), .ZN(G305));
  NAND2_X1  g177(.A1(new_n587), .A2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n565), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(new_n507), .B2(G85), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G290));
  XNOR2_X1  g183(.A(KEYINPUT75), .B(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n509), .A2(new_n518), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n507), .A2(G92), .A3(new_n609), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n565), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n613), .A2(new_n614), .B1(G651), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n587), .A2(G54), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n583), .ZN(G284));
  AOI21_X1  g197(.A(new_n621), .B1(G868), .B2(new_n583), .ZN(G321));
  NOR2_X1   g198(.A1(G299), .A2(G868), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n590), .B2(G868), .ZN(G297));
  AOI21_X1  g200(.A(new_n624), .B1(new_n590), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G860), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n620), .B1(G559), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT76), .ZN(G148));
  OR2_X1    g204(.A1(new_n620), .A2(G559), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n555), .B2(G868), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n474), .A2(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n474), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n476), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n463), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G2096), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n638), .A2(new_n639), .A3(new_n646), .ZN(G156));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT79), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT78), .B(G2438), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2430), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n650), .B(new_n651), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(new_n654), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n658), .A3(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2451), .B(G2454), .Z(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n662), .B(new_n663), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(new_n665), .B2(new_n668), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n665), .A2(new_n668), .ZN(new_n673));
  INV_X1    g248(.A(G14), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n648), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n648), .C1(new_n671), .C2(new_n670), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(G401));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT82), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2072), .B(G2078), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT83), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT18), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n681), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n681), .A2(new_n683), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n682), .B(KEYINPUT17), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n682), .B(KEYINPUT84), .Z(new_n691));
  OAI211_X1 g266(.A(new_n686), .B(new_n690), .C1(new_n687), .C2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(new_n645), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT85), .B(G2100), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n692), .B(G2096), .ZN(new_n696));
  INV_X1    g271(.A(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(G227));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1956), .B(G2474), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT86), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1961), .B(G1966), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n702), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT20), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n702), .B1(new_n704), .B2(new_n706), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n704), .A2(new_n706), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n708), .B(new_n711), .C1(new_n701), .C2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1991), .B(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G24), .ZN(new_n720));
  INV_X1    g295(.A(G290), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  INV_X1    g297(.A(G1986), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n474), .A2(G131), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT87), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n476), .A2(G119), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n463), .A2(G107), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G25), .B(new_n730), .S(G29), .Z(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n719), .A2(G23), .ZN(new_n734));
  INV_X1    g309(.A(G288), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n719), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT33), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1976), .ZN(new_n738));
  MUX2_X1   g313(.A(G6), .B(G305), .S(G16), .Z(new_n739));
  XOR2_X1   g314(.A(KEYINPUT32), .B(G1981), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n719), .A2(G22), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT88), .Z(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G303), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1971), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n738), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n724), .B(new_n733), .C1(new_n747), .C2(KEYINPUT34), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(KEYINPUT34), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G27), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G164), .B2(new_n755), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2078), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT26), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G129), .B2(new_n476), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n755), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n755), .B2(G32), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT93), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n766), .A2(new_n768), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT30), .B(G28), .ZN(new_n771));
  OR2_X1    g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  NAND2_X1  g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n771), .A2(new_n755), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n644), .B2(new_n755), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n758), .A2(new_n769), .A3(new_n770), .A4(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G34), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(KEYINPUT24), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(KEYINPUT24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n755), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G160), .B2(new_n755), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2084), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n719), .A2(G20), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT23), .ZN(new_n784));
  INV_X1    g359(.A(G299), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n719), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT95), .B(G1956), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n755), .A2(G35), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G162), .B2(new_n755), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT29), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2090), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n755), .A2(G33), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n462), .A2(G127), .ZN(new_n795));
  NAND2_X1  g370(.A1(G115), .A2(G2104), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n463), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G139), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n482), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT25), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n797), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n794), .B1(new_n802), .B2(new_n755), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2072), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n719), .A2(G5), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G171), .B2(new_n719), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1961), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n755), .A2(G26), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT28), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n474), .A2(G140), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n476), .A2(G128), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n463), .A2(G116), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n809), .B1(new_n814), .B2(G29), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT92), .B(G2067), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n804), .A2(new_n807), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n776), .A2(new_n789), .A3(new_n793), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G4), .A2(G16), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n618), .A2(new_n619), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(G16), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT91), .B(G1348), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n822), .B(new_n823), .Z(new_n824));
  OAI21_X1  g399(.A(new_n588), .B1(new_n526), .B2(new_n525), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n719), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT94), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G16), .B2(G21), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1966), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n719), .A2(G19), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n555), .B2(new_n719), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1341), .ZN(new_n834));
  NOR4_X1   g409(.A1(new_n819), .A2(new_n824), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n754), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(G311));
  AND2_X1   g413(.A1(new_n750), .A2(new_n751), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n754), .B(new_n835), .C1(new_n839), .C2(new_n752), .ZN(G150));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  INV_X1    g416(.A(G67), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n565), .B2(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n843), .A2(G651), .B1(new_n507), .B2(G93), .ZN(new_n844));
  OAI21_X1  g419(.A(G55), .B1(new_n529), .B2(new_n531), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT97), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n821), .A2(G559), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n851));
  XOR2_X1   g426(.A(new_n850), .B(new_n851), .Z(new_n852));
  INV_X1    g427(.A(new_n546), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n548), .B1(new_n547), .B2(new_n550), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n553), .A2(KEYINPUT71), .A3(new_n549), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n846), .ZN(new_n857));
  INV_X1    g432(.A(new_n846), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n555), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n852), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n627), .B1(new_n862), .B2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n849), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT98), .Z(G145));
  XNOR2_X1  g441(.A(new_n730), .B(new_n635), .ZN(new_n867));
  AOI22_X1  g442(.A1(G130), .A2(new_n476), .B1(new_n474), .B2(G142), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n869), .A2(KEYINPUT101), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n871), .A2(new_n463), .A3(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n463), .B2(G118), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n872), .B(new_n873), .C1(KEYINPUT101), .C2(new_n869), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n868), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n867), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n802), .B(new_n763), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n814), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n492), .A2(KEYINPUT99), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n487), .A2(new_n491), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n814), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n879), .B2(new_n884), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n877), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n644), .B(new_n480), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n471), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n877), .B2(new_n888), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  INV_X1    g469(.A(new_n887), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(new_n885), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n886), .A2(KEYINPUT102), .A3(new_n887), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n876), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n893), .B1(new_n898), .B2(KEYINPUT103), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n898), .A2(KEYINPUT103), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n892), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g477(.A(G303), .B(new_n721), .ZN(new_n903));
  XNOR2_X1  g478(.A(G305), .B(new_n735), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT42), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n821), .A2(G299), .ZN(new_n907));
  AOI21_X1  g482(.A(G299), .B1(new_n618), .B2(new_n619), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n620), .A2(new_n785), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n912), .B2(new_n908), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n907), .A2(new_n909), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(KEYINPUT104), .A3(new_n911), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n916), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n860), .B(new_n630), .ZN(new_n921));
  MUX2_X1   g496(.A(new_n919), .B(new_n920), .S(new_n921), .Z(new_n922));
  XNOR2_X1  g497(.A(new_n906), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(G868), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(G868), .B2(new_n858), .ZN(G295));
  OAI21_X1  g500(.A(new_n924), .B1(G868), .B2(new_n858), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  INV_X1    g502(.A(new_n905), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n586), .A2(G171), .A3(new_n589), .ZN(new_n929));
  NAND4_X1  g504(.A1(G168), .A2(KEYINPUT105), .A3(new_n575), .A4(new_n582), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n583), .B2(new_n825), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n860), .A2(new_n929), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n932), .A3(new_n930), .ZN(new_n934));
  AOI211_X1 g509(.A(new_n546), .B(new_n846), .C1(new_n554), .C2(new_n551), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n551), .A2(new_n554), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n858), .B1(new_n936), .B2(new_n853), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n910), .A2(new_n913), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n933), .A2(new_n939), .A3(KEYINPUT106), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n934), .A2(new_n938), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n920), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI211_X1 g523(.A(KEYINPUT107), .B(new_n920), .C1(new_n943), .C2(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n928), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n943), .A2(new_n918), .A3(new_n945), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n933), .A2(new_n939), .A3(new_n916), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n905), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(KEYINPUT43), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n953), .A2(new_n954), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n905), .B1(new_n951), .B2(new_n952), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT44), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n950), .A2(new_n957), .A3(new_n955), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n958), .B2(new_n959), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n927), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n956), .B2(new_n960), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n963), .B2(new_n964), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT108), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(G397));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n880), .A2(new_n973), .A3(new_n882), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n466), .A2(G40), .A3(new_n468), .A4(new_n470), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n978), .A2(KEYINPUT111), .A3(new_n979), .A4(new_n764), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(new_n982), .B2(new_n763), .ZN(new_n983));
  INV_X1    g558(.A(new_n978), .ZN(new_n984));
  INV_X1    g559(.A(G2067), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n814), .B(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(G1996), .B2(new_n763), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n980), .B(new_n983), .C1(new_n984), .C2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n989), .A2(KEYINPUT112), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(KEYINPUT112), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n730), .B(new_n732), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT113), .Z(new_n993));
  OAI211_X1 g568(.A(new_n990), .B(new_n991), .C1(new_n984), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n721), .A2(new_n723), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT110), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n723), .B2(new_n721), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n994), .B1(new_n978), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n735), .A2(G1976), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n492), .A2(new_n973), .ZN(new_n1000));
  OAI211_X1 g575(.A(G8), .B(new_n999), .C1(new_n1000), .C2(new_n977), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1001), .A2(KEYINPUT52), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n1002), .A2(KEYINPUT115), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(KEYINPUT115), .ZN(new_n1004));
  XNOR2_X1  g579(.A(G305), .B(G1981), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n1000), .B2(new_n977), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1003), .A2(new_n1004), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n735), .A2(G1976), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1001), .A2(KEYINPUT52), .A3(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT116), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g590(.A1(G303), .A2(G8), .B1(KEYINPUT114), .B2(KEYINPUT55), .ZN(new_n1016));
  NOR2_X1   g591(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n977), .B1(new_n1000), .B2(new_n975), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n880), .A2(KEYINPUT45), .A3(new_n973), .A4(new_n882), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1971), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1022));
  INV_X1    g597(.A(new_n977), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n492), .A2(new_n1024), .A3(new_n973), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(G2090), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1018), .B(G8), .C1(new_n1021), .C2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g603(.A(G1976), .B(G288), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G305), .A2(G1981), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI22_X1  g606(.A1(new_n1015), .A2(new_n1028), .B1(new_n1031), .B2(new_n1009), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1016), .B(new_n1017), .Z(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT119), .ZN(new_n1034));
  OAI21_X1  g609(.A(G8), .B1(new_n1027), .B2(new_n1021), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1026), .A2(G2084), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n977), .B1(new_n1000), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n975), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n492), .A2(new_n973), .A3(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(KEYINPUT118), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(KEYINPUT118), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1966), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1037), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1046), .A2(new_n1047), .A3(G286), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1036), .A2(new_n1014), .A3(new_n1011), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1032), .B1(new_n1049), .B2(KEYINPUT63), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1011), .A2(new_n1014), .A3(new_n1051), .A4(new_n1028), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(G2084), .B2(new_n1026), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1054), .B2(new_n825), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1046), .A2(G168), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT51), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1047), .B1(new_n1046), .B2(G168), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1052), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1063), .B2(G2078), .ZN(new_n1064));
  INV_X1    g639(.A(G1961), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1026), .A2(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n976), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G2078), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n977), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1020), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT126), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT126), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n976), .A2(new_n1075), .A3(new_n1020), .A4(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1067), .A2(new_n1077), .A3(G301), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1064), .B(new_n1066), .C1(new_n1044), .C2(new_n1071), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n583), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT127), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1067), .A2(new_n1077), .ZN(new_n1085));
  INV_X1    g660(.A(G171), .ZN(new_n1086));
  OAI221_X1 g661(.A(KEYINPUT54), .B1(new_n583), .B2(new_n1079), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT127), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1081), .A2(new_n1088), .A3(new_n1082), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1061), .A2(new_n1084), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1026), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1019), .A2(new_n1020), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(G299), .A2(KEYINPUT120), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT57), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1000), .A2(new_n977), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1026), .A2(new_n823), .B1(new_n985), .B2(new_n1100), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(new_n620), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1092), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1099), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1101), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n821), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT124), .B1(new_n1101), .B2(KEYINPUT60), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n620), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n555), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT121), .B(G1996), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1019), .A2(new_n1020), .A3(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT58), .B(G1341), .Z(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1000), .B2(new_n977), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1119), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1116), .A2(KEYINPUT61), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1115), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1099), .A2(KEYINPUT61), .A3(new_n1103), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT123), .Z(new_n1132));
  AOI21_X1  g707(.A(new_n1105), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1050), .B1(new_n1090), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1055), .A2(KEYINPUT51), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1054), .A2(new_n825), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1059), .B1(new_n1058), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT62), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1057), .A2(new_n1139), .A3(new_n1060), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1080), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1048), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1052), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n998), .B1(new_n1134), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n978), .B1(new_n763), .B2(new_n987), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n982), .A2(KEYINPUT46), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n982), .A2(KEYINPUT46), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT47), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n984), .A2(new_n996), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT48), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n994), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n732), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n730), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n990), .A2(new_n991), .A3(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n814), .A2(G2067), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n984), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1146), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g736(.A1(new_n695), .A2(new_n698), .A3(new_n456), .ZN(new_n1163));
  NOR2_X1   g737(.A1(new_n1163), .A2(G229), .ZN(new_n1164));
  OAI211_X1 g738(.A(new_n901), .B(new_n1164), .C1(new_n676), .C2(new_n678), .ZN(new_n1165));
  AOI21_X1  g739(.A(new_n1165), .B1(new_n964), .B2(new_n963), .ZN(G308));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1167), .A2(new_n965), .ZN(G225));
endmodule


