//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n208), .B1(G155gat), .B2(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(KEYINPUT76), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n207), .A2(new_n210), .A3(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n205), .A2(new_n206), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n220), .B(new_n214), .C1(new_n221), .C2(new_n209), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G197gat), .B(G204gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT72), .B(G211gat), .ZN(new_n225));
  INV_X1    g024(.A(G218gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n224), .B1(new_n227), .B2(KEYINPUT22), .ZN(new_n228));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(KEYINPUT73), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n230), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT29), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n223), .B1(new_n233), .B2(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n232), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n222), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT29), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n202), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n228), .A2(new_n229), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT29), .B1(new_n228), .B2(new_n229), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n244), .A2(new_n236), .B1(new_n217), .B2(new_n222), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n235), .A2(new_n239), .ZN(new_n246));
  INV_X1    g045(.A(new_n202), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G22gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(G22gat), .B1(new_n241), .B2(new_n248), .ZN(new_n252));
  XNOR2_X1  g051(.A(G78gat), .B(G106gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT31), .B(G50gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n256), .A2(KEYINPUT87), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(KEYINPUT87), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n251), .A2(new_n252), .ZN(new_n259));
  INV_X1    g058(.A(new_n255), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT88), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n262));
  AOI211_X1 g061(.A(new_n262), .B(new_n255), .C1(new_n251), .C2(new_n252), .ZN(new_n263));
  OAI22_X1  g062(.A1(new_n257), .A2(new_n258), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT23), .ZN(new_n266));
  INV_X1    g065(.A(G169gat), .ZN(new_n267));
  INV_X1    g066(.A(G176gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT23), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT25), .ZN(new_n273));
  INV_X1    g072(.A(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT24), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT24), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(G183gat), .A3(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(G183gat), .B2(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT64), .B(G190gat), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n282), .A2(new_n274), .B1(new_n276), .B2(new_n278), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT25), .B1(new_n283), .B2(new_n272), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n269), .A2(KEYINPUT26), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n265), .B1(new_n269), .B2(KEYINPUT26), .ZN(new_n288));
  OAI22_X1  g087(.A1(new_n287), .A2(new_n288), .B1(new_n274), .B2(new_n275), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT27), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT65), .B1(new_n290), .B2(G183gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT27), .B(G183gat), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n282), .B(new_n291), .C1(new_n292), .C2(KEYINPUT65), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n282), .A3(KEYINPUT28), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n289), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  INV_X1    g098(.A(G113gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(G120gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(G113gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n300), .A2(KEYINPUT67), .A3(G120gat), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n301), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G127gat), .ZN(new_n309));
  INV_X1    g108(.A(G127gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G134gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT1), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n300), .A2(G120gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n303), .A2(G113gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n309), .A2(new_n311), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n285), .A2(new_n298), .A3(KEYINPUT68), .A4(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n294), .A2(new_n293), .B1(new_n323), .B2(new_n292), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n284), .B(new_n281), .C1(new_n324), .C2(new_n289), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n320), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G227gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n325), .B2(new_n320), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT71), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT33), .ZN(new_n334));
  XNOR2_X1  g133(.A(G15gat), .B(G43gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT69), .ZN(new_n336));
  XNOR2_X1  g135(.A(G71gat), .B(G99gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n334), .B1(new_n338), .B2(KEYINPUT70), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(KEYINPUT70), .B2(new_n338), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT32), .ZN(new_n341));
  INV_X1    g140(.A(new_n329), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n331), .A2(new_n322), .A3(new_n326), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n342), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n334), .A2(KEYINPUT32), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n338), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT34), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n344), .A2(new_n348), .A3(KEYINPUT34), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n333), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n344), .A2(new_n348), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT34), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n355), .A2(KEYINPUT71), .A3(new_n332), .A4(new_n349), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n358));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n325), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n359), .B1(new_n285), .B2(new_n298), .ZN(new_n363));
  INV_X1    g162(.A(new_n235), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n281), .A2(new_n284), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n361), .B1(new_n366), .B2(new_n297), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n359), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n325), .A2(new_n360), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n235), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n358), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT75), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  OAI21_X1  g174(.A(new_n364), .B1(new_n362), .B2(new_n363), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n368), .A2(new_n235), .A3(new_n369), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT74), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n371), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n375), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n365), .A2(new_n370), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(KEYINPUT30), .A3(new_n380), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n379), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n264), .A2(new_n357), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(KEYINPUT35), .ZN(new_n389));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT0), .ZN(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(KEYINPUT84), .B(KEYINPUT6), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n217), .B2(new_n222), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n238), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n320), .A2(KEYINPUT77), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n314), .A2(new_n319), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n399), .A2(KEYINPUT79), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n400), .A2(new_n404), .A3(new_n402), .A4(new_n237), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n314), .A2(new_n319), .A3(new_n217), .A4(new_n222), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n412));
  AND3_X1   g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n410), .A2(KEYINPUT4), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n411), .B1(new_n410), .B2(new_n412), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n408), .A2(new_n409), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n402), .A3(new_n223), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT82), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n400), .A2(new_n421), .A3(new_n402), .A4(new_n223), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n410), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n409), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT5), .ZN(new_n427));
  INV_X1    g226(.A(new_n410), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n419), .B2(KEYINPUT82), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n409), .B1(new_n429), .B2(new_n422), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT83), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n418), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n412), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(KEYINPUT4), .B2(new_n428), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n408), .A2(new_n436), .A3(new_n431), .A4(new_n409), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n394), .B(new_n396), .C1(new_n433), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT85), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n426), .B1(new_n425), .B2(KEYINPUT5), .ZN(new_n441));
  AOI211_X1 g240(.A(KEYINPUT83), .B(new_n431), .C1(new_n423), .C2(new_n424), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n417), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n437), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n394), .A4(new_n396), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n394), .B1(new_n433), .B2(new_n438), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT90), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(KEYINPUT90), .A3(new_n394), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n443), .A2(new_n393), .A3(new_n437), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n395), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n389), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n452), .A3(new_n395), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n440), .A3(new_n446), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n457), .A2(new_n458), .A3(new_n387), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n457), .B2(new_n387), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n264), .A2(new_n357), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n455), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n384), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n375), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT37), .B1(new_n377), .B2(KEYINPUT92), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(new_n384), .B2(KEYINPUT92), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n381), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n371), .A2(KEYINPUT37), .A3(new_n378), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n375), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT93), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT93), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n475), .A3(new_n375), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n476), .A3(new_n466), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n471), .B1(new_n477), .B2(KEYINPUT38), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(new_n447), .A3(new_n453), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n429), .A2(new_n409), .A3(new_n422), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n435), .B1(new_n403), .B2(new_n407), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n480), .B(KEYINPUT39), .C1(new_n481), .C2(new_n409), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n408), .A2(new_n436), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n424), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT89), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT40), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n482), .A2(new_n485), .A3(new_n393), .A4(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n386), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n482), .A2(new_n485), .A3(new_n393), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n487), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n490), .A2(new_n450), .A3(new_n451), .A4(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n493), .A2(KEYINPUT91), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(KEYINPUT91), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n479), .B(new_n264), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n264), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n459), .B2(new_n460), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n357), .B(KEYINPUT36), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n464), .A2(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(G71gat), .A2(G78gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(G71gat), .A2(G78gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n502), .B(new_n503), .C1(KEYINPUT104), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n504), .ZN(new_n506));
  OR2_X1    g305(.A1(G57gat), .A2(G64gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(G57gat), .A2(G64gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n505), .B(new_n509), .Z(new_n510));
  INV_X1    g309(.A(KEYINPUT21), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G231gat), .A2(G233gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(G127gat), .B(G155gat), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT20), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n514), .B(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G183gat), .B(G211gat), .Z(new_n518));
  XOR2_X1   g317(.A(new_n517), .B(new_n518), .Z(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n250), .A2(G15gat), .ZN(new_n521));
  INV_X1    g320(.A(G15gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G22gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT99), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT99), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT16), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n525), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(G1gat), .B1(new_n525), .B2(new_n528), .ZN(new_n532));
  OAI211_X1 g331(.A(KEYINPUT100), .B(new_n520), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n526), .A2(new_n527), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n521), .A2(new_n523), .A3(new_n527), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n529), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n520), .A2(KEYINPUT100), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n525), .A2(new_n528), .A3(new_n530), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n520), .A2(KEYINPUT100), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n533), .A2(KEYINPUT101), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT101), .B1(new_n533), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n511), .B2(new_n510), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT105), .B(KEYINPUT19), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n519), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n519), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n540), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  INV_X1    g352(.A(G50gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(G43gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT97), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT15), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G43gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G50gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(G43gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT97), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT98), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(KEYINPUT98), .A3(new_n561), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT15), .ZN(new_n567));
  NAND2_X1  g366(.A1(G29gat), .A2(G36gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n567), .B(new_n568), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n571), .B1(KEYINPUT96), .B2(new_n569), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(KEYINPUT96), .B2(new_n569), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n568), .ZN(new_n577));
  INV_X1    g376(.A(new_n567), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n553), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n572), .B1(new_n564), .B2(new_n565), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n567), .B1(new_n576), .B2(new_n568), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT17), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n552), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT101), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n552), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n533), .A2(KEYINPUT101), .A3(new_n540), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n581), .A2(new_n582), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT102), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT102), .ZN(new_n595));
  AOI211_X1 g394(.A(new_n595), .B(new_n592), .C1(new_n589), .C2(new_n590), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n587), .B(KEYINPUT18), .C1(new_n594), .C2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT103), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n595), .B1(new_n543), .B2(new_n592), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n591), .A2(KEYINPUT102), .A3(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n602), .A2(KEYINPUT103), .A3(KEYINPUT18), .A4(new_n587), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n587), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT18), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n543), .A2(new_n592), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n594), .B2(new_n596), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n585), .B(KEYINPUT13), .Z(new_n609));
  AOI22_X1  g408(.A1(new_n605), .A2(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT94), .B(G197gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT11), .B(G169gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n604), .A2(new_n610), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(KEYINPUT95), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(new_n604), .B2(new_n610), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n580), .A2(new_n583), .ZN(new_n622));
  OR2_X1    g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT107), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT107), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n627), .A3(new_n624), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(KEYINPUT106), .A2(G85gat), .A3(G92gat), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT7), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(KEYINPUT106), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n624), .A2(KEYINPUT8), .ZN(new_n634));
  OR2_X1    g433(.A1(G85gat), .A2(G92gat), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n629), .A2(new_n636), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n622), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n593), .A2(new_n640), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n643));
  NAND2_X1  g442(.A1(G232gat), .A2(G233gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G190gat), .B(G218gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G134gat), .B(G162gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n643), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(KEYINPUT108), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n651), .A2(KEYINPUT108), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n648), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n648), .A2(new_n652), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G230gat), .A2(G233gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n510), .B1(new_n638), .B2(new_n639), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n629), .A2(new_n636), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n505), .B(new_n509), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n661), .A3(new_n637), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n640), .A2(KEYINPUT10), .A3(new_n661), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n658), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n657), .B1(new_n659), .B2(new_n662), .ZN(new_n667));
  XNOR2_X1  g466(.A(G120gat), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT109), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  OR3_X1    g470(.A1(new_n666), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT110), .Z(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n664), .B2(new_n665), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n671), .B1(new_n674), .B2(new_n667), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NOR4_X1   g475(.A1(new_n551), .A2(new_n621), .A3(new_n656), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n501), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n457), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(new_n529), .ZN(G1324gat));
  NAND3_X1  g479(.A1(new_n501), .A2(new_n386), .A3(new_n677), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT16), .B(G8gat), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(G8gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n684), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(G1325gat));
  OAI21_X1  g487(.A(G15gat), .B1(new_n678), .B2(new_n499), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n357), .A2(new_n522), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n678), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n678), .A2(new_n264), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  OR2_X1    g493(.A1(new_n654), .A2(new_n655), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n464), .B2(new_n500), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(KEYINPUT44), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n621), .A2(new_n550), .A3(new_n676), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701), .B2(new_n457), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n696), .A2(new_n700), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n457), .A2(G29gat), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n703), .A2(KEYINPUT111), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT111), .B1(new_n703), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(KEYINPUT45), .A3(new_n707), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n702), .A2(new_n710), .A3(new_n711), .ZN(G1328gat));
  OAI21_X1  g511(.A(G36gat), .B1(new_n701), .B2(new_n387), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n387), .A2(G36gat), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT46), .B1(new_n703), .B2(new_n715), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n703), .A2(KEYINPUT46), .A3(new_n715), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(G1329gat));
  INV_X1    g517(.A(new_n499), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n697), .A2(new_n719), .A3(new_n700), .A4(new_n698), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G43gat), .ZN(new_n721));
  INV_X1    g520(.A(new_n703), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n558), .A3(new_n357), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n721), .A2(KEYINPUT47), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1330gat));
  NAND4_X1  g527(.A1(new_n697), .A2(new_n497), .A3(new_n700), .A4(new_n698), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G50gat), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n264), .A2(G50gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT112), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n722), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n730), .A2(KEYINPUT48), .A3(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1331gat));
  NAND3_X1  g537(.A1(new_n621), .A2(new_n550), .A3(new_n695), .ZN(new_n739));
  INV_X1    g538(.A(new_n676), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT113), .B1(new_n501), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743));
  INV_X1    g542(.A(new_n741), .ZN(new_n744));
  AOI211_X1 g543(.A(new_n743), .B(new_n744), .C1(new_n464), .C2(new_n500), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n457), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g548(.A(new_n387), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT114), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n752), .B(new_n753), .Z(G1333gat));
  AND3_X1   g553(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n457), .A2(new_n387), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT86), .ZN(new_n757));
  INV_X1    g556(.A(new_n461), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n457), .A2(new_n458), .A3(new_n387), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n760), .A2(KEYINPUT35), .B1(new_n454), .B2(new_n389), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n741), .B1(new_n755), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n743), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n501), .A2(KEYINPUT113), .A3(new_n741), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(new_n357), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(G71gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n499), .A2(new_n766), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n746), .B2(new_n769), .ZN(new_n770));
  AND4_X1   g569(.A1(new_n768), .A2(new_n763), .A3(new_n764), .A4(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT50), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n774), .B(new_n767), .C1(new_n770), .C2(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n746), .A2(new_n497), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n551), .A2(new_n621), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT116), .Z(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n740), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n699), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n457), .ZN(new_n783));
  INV_X1    g582(.A(new_n780), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n696), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT51), .B1(new_n696), .B2(new_n784), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n457), .A2(G85gat), .A3(new_n740), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(G1336gat));
  NAND4_X1  g588(.A1(new_n697), .A2(new_n386), .A3(new_n698), .A4(new_n781), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G92gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n387), .A2(G92gat), .A3(new_n740), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n785), .B2(new_n786), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT52), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n791), .A2(new_n796), .A3(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n782), .B2(new_n499), .ZN(new_n799));
  INV_X1    g598(.A(G99gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n357), .A2(new_n800), .A3(new_n676), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n787), .B2(new_n801), .ZN(G1338gat));
  NAND4_X1  g601(.A1(new_n697), .A2(new_n497), .A3(new_n698), .A4(new_n781), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G106gat), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n264), .A2(G106gat), .A3(new_n740), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n785), .B2(new_n786), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n804), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(G1339gat));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n664), .A2(new_n665), .A3(new_n673), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n814), .A2(new_n666), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n664), .A2(new_n665), .ZN(new_n817));
  INV_X1    g616(.A(new_n673), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n671), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n813), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n666), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n664), .A2(new_n665), .A3(new_n673), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n671), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n674), .B2(new_n815), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n821), .A2(new_n672), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT117), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n821), .A2(new_n827), .A3(new_n830), .A4(new_n672), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n604), .A2(new_n610), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n618), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n604), .A2(new_n610), .A3(new_n616), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT118), .B1(new_n608), .B2(new_n609), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n602), .A2(new_n584), .ZN(new_n838));
  INV_X1    g637(.A(new_n585), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  INV_X1    g640(.A(new_n609), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n602), .A2(new_n841), .A3(new_n607), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n837), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n615), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(new_n835), .A3(new_n676), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n812), .B1(new_n836), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n829), .A2(new_n831), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n617), .B2(new_n620), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(new_n835), .A3(new_n676), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(KEYINPUT119), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n851), .A3(new_n695), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n656), .A2(new_n848), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n845), .A2(new_n835), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n550), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n621), .A2(new_n550), .A3(new_n695), .A4(new_n740), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(new_n457), .A3(new_n388), .ZN(new_n861));
  INV_X1    g660(.A(new_n621), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n676), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g665(.A1(new_n861), .A2(new_n550), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n310), .A2(KEYINPUT120), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n867), .B(new_n868), .ZN(G1342gat));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n861), .B(new_n656), .C1(new_n870), .C2(new_n308), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n308), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n871), .B(new_n872), .ZN(G1343gat));
  OAI21_X1  g672(.A(new_n850), .B1(new_n621), .B2(new_n828), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n695), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n856), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n859), .B1(new_n876), .B2(new_n551), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n877), .A2(new_n878), .A3(new_n264), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n849), .A2(new_n850), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n656), .B1(new_n880), .B2(new_n812), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n855), .B1(new_n881), .B2(new_n851), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n858), .B1(new_n882), .B2(new_n550), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n497), .ZN(new_n884));
  XOR2_X1   g683(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n885));
  AOI21_X1  g684(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n719), .A2(new_n457), .A3(new_n386), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n621), .A2(new_n203), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n886), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n860), .A2(new_n264), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n887), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n203), .B1(new_n894), .B2(new_n621), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(KEYINPUT58), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  INV_X1    g696(.A(new_n895), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n891), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(G1344gat));
  INV_X1    g699(.A(new_n894), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n204), .A3(new_n676), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G148gat), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n886), .A2(new_n888), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n676), .ZN(new_n906));
  INV_X1    g705(.A(new_n885), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n883), .A2(new_n497), .A3(new_n907), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n858), .B(KEYINPUT122), .Z(new_n909));
  OR3_X1    g708(.A1(new_n695), .A2(new_n854), .A3(new_n828), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n550), .B1(new_n875), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n497), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n878), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n676), .A3(new_n887), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n903), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n902), .B1(new_n906), .B2(new_n916), .ZN(G1345gat));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n211), .A3(new_n550), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n886), .A2(new_n551), .A3(new_n888), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n211), .ZN(G1346gat));
  NAND2_X1  g719(.A1(new_n656), .A2(new_n212), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n894), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n886), .A2(new_n695), .A3(new_n888), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n923), .A2(new_n924), .B1(new_n212), .B2(new_n925), .ZN(G1347gat));
  NAND2_X1  g725(.A1(new_n758), .A2(new_n386), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n457), .B(new_n928), .C1(new_n857), .C2(new_n859), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n267), .A3(new_n621), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n457), .B1(new_n857), .B2(new_n859), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(KEYINPUT124), .B(new_n457), .C1(new_n857), .C2(new_n859), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n862), .A3(new_n928), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n930), .B1(new_n936), .B2(new_n267), .ZN(G1348gat));
  OAI21_X1  g736(.A(G176gat), .B1(new_n929), .B2(new_n740), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n928), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n676), .A2(new_n268), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(G1349gat));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  OR3_X1    g741(.A1(new_n929), .A2(new_n942), .A3(new_n551), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n929), .B2(new_n551), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(G183gat), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n935), .A2(new_n292), .A3(new_n550), .A4(new_n928), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT60), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n929), .B2(new_n695), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n656), .A2(new_n282), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n939), .B2(new_n954), .ZN(G1351gat));
  NAND2_X1  g754(.A1(new_n499), .A2(new_n386), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(new_n747), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n958), .B1(new_n908), .B2(new_n913), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n621), .ZN(new_n961));
  INV_X1    g760(.A(new_n956), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n497), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n963), .B1(new_n933), .B2(new_n934), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n621), .A2(G197gat), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n965), .B1(new_n964), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n961), .B1(new_n967), .B2(new_n968), .ZN(G1352gat));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  INV_X1    g770(.A(new_n963), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n740), .A2(G204gat), .ZN(new_n973));
  AND4_X1   g772(.A1(new_n971), .A2(new_n935), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n971), .B1(new_n964), .B2(new_n973), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n935), .A2(new_n972), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n964), .A2(new_n971), .A3(new_n973), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT62), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n914), .A2(new_n676), .A3(new_n957), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G204gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n976), .A2(new_n980), .A3(new_n982), .ZN(G1353gat));
  NAND3_X1  g782(.A1(new_n964), .A2(new_n225), .A3(new_n550), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n959), .A2(new_n550), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1354gat));
  OAI21_X1  g787(.A(G218gat), .B1(new_n960), .B2(new_n695), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n964), .A2(new_n226), .A3(new_n656), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1355gat));
endmodule


