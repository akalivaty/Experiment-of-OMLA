

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752;

  XNOR2_X1 U372 ( .A(G143), .B(G128), .ZN(n497) );
  NAND2_X1 U373 ( .A1(n351), .A2(n363), .ZN(n365) );
  NAND2_X1 U374 ( .A1(n367), .A2(n368), .ZN(n351) );
  NOR2_X1 U375 ( .A1(n721), .A2(G902), .ZN(n440) );
  AND2_X4 U376 ( .A1(n365), .A2(n369), .ZN(n717) );
  OR2_X2 U377 ( .A1(n603), .A2(n385), .ZN(n384) );
  XNOR2_X2 U378 ( .A(n593), .B(n592), .ZN(n603) );
  XNOR2_X2 U379 ( .A(n567), .B(n423), .ZN(n681) );
  XNOR2_X2 U380 ( .A(n440), .B(n439), .ZN(n507) );
  XNOR2_X2 U381 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n449) );
  AND2_X1 U382 ( .A1(n639), .A2(n638), .ZN(n641) );
  INV_X1 U383 ( .A(n742), .ZN(n368) );
  XNOR2_X1 U384 ( .A(n515), .B(KEYINPUT32), .ZN(n625) );
  NOR2_X1 U385 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U386 ( .A1(n567), .A2(n527), .ZN(n574) );
  XNOR2_X1 U387 ( .A(n497), .B(KEYINPUT4), .ZN(n452) );
  INV_X1 U388 ( .A(G953), .ZN(n743) );
  INV_X1 U389 ( .A(G146), .ZN(n428) );
  NOR2_X1 U390 ( .A1(n726), .A2(KEYINPUT2), .ZN(n674) );
  NOR2_X2 U391 ( .A1(n645), .A2(n725), .ZN(n648) );
  XNOR2_X2 U392 ( .A(n534), .B(n475), .ZN(n529) );
  BUF_X1 U393 ( .A(n614), .Z(n726) );
  XNOR2_X2 U394 ( .A(n474), .B(KEYINPUT0), .ZN(n534) );
  NOR2_X2 U395 ( .A1(n570), .A2(n473), .ZN(n474) );
  AND2_X1 U396 ( .A1(n750), .A2(n372), .ZN(n382) );
  OR2_X1 U397 ( .A1(n617), .A2(G902), .ZN(n422) );
  NAND2_X1 U398 ( .A1(n368), .A2(n364), .ZN(n369) );
  AND2_X1 U399 ( .A1(n726), .A2(KEYINPUT2), .ZN(n364) );
  AND2_X1 U400 ( .A1(n383), .A2(n381), .ZN(n380) );
  AND2_X1 U401 ( .A1(n378), .A2(n376), .ZN(n375) );
  XNOR2_X1 U402 ( .A(n452), .B(n403), .ZN(n741) );
  XNOR2_X1 U403 ( .A(G104), .B(KEYINPUT75), .ZN(n415) );
  XNOR2_X1 U404 ( .A(n428), .B(n741), .ZN(n421) );
  XNOR2_X1 U405 ( .A(G110), .B(G107), .ZN(n454) );
  XNOR2_X1 U406 ( .A(n390), .B(KEYINPUT28), .ZN(n568) );
  NOR2_X1 U407 ( .A1(n562), .A2(n391), .ZN(n390) );
  INV_X1 U408 ( .A(KEYINPUT91), .ZN(n475) );
  NAND2_X1 U409 ( .A1(n679), .A2(n369), .ZN(n370) );
  XNOR2_X1 U410 ( .A(KEYINPUT77), .B(n678), .ZN(n679) );
  NOR2_X1 U411 ( .A1(n373), .A2(n372), .ZN(n371) );
  NAND2_X1 U412 ( .A1(n688), .A2(n392), .ZN(n391) );
  INV_X1 U413 ( .A(n566), .ZN(n392) );
  XNOR2_X1 U414 ( .A(KEYINPUT3), .B(G119), .ZN(n404) );
  XOR2_X1 U415 ( .A(G113), .B(G116), .Z(n405) );
  XNOR2_X1 U416 ( .A(G128), .B(G119), .ZN(n424) );
  XOR2_X1 U417 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n425) );
  XOR2_X1 U418 ( .A(G122), .B(G107), .Z(n494) );
  XNOR2_X1 U419 ( .A(G134), .B(G116), .ZN(n493) );
  XNOR2_X1 U420 ( .A(n394), .B(n393), .ZN(n502) );
  XNOR2_X1 U421 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n393) );
  XNOR2_X1 U422 ( .A(n395), .B(KEYINPUT67), .ZN(n394) );
  NAND2_X1 U423 ( .A1(n743), .A2(G234), .ZN(n395) );
  XNOR2_X1 U424 ( .A(n398), .B(n397), .ZN(n367) );
  INV_X1 U425 ( .A(KEYINPUT80), .ZN(n397) );
  INV_X1 U426 ( .A(G143), .ZN(n485) );
  XNOR2_X1 U427 ( .A(n421), .B(n420), .ZN(n617) );
  XNOR2_X1 U428 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U429 ( .A(n354), .B(n417), .ZN(n418) );
  NAND2_X1 U430 ( .A1(n665), .A2(KEYINPUT40), .ZN(n387) );
  BUF_X1 U431 ( .A(n563), .Z(n590) );
  INV_X1 U432 ( .A(KEYINPUT34), .ZN(n401) );
  INV_X1 U433 ( .A(n562), .ZN(n684) );
  AND2_X1 U434 ( .A1(n620), .A2(G953), .ZN(n725) );
  NAND2_X1 U435 ( .A1(n717), .A2(G210), .ZN(n637) );
  XNOR2_X1 U436 ( .A(n597), .B(n389), .ZN(n750) );
  XNOR2_X1 U437 ( .A(n598), .B(KEYINPUT114), .ZN(n389) );
  XNOR2_X1 U438 ( .A(n533), .B(KEYINPUT100), .ZN(n654) );
  AND2_X1 U439 ( .A1(n370), .A2(n352), .ZN(n716) );
  NOR2_X1 U440 ( .A1(n711), .A2(n360), .ZN(n352) );
  XOR2_X1 U441 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n353) );
  XOR2_X1 U442 ( .A(n406), .B(G101), .Z(n354) );
  XNOR2_X1 U443 ( .A(n426), .B(KEYINPUT71), .ZN(n355) );
  OR2_X1 U444 ( .A1(G902), .A2(n718), .ZN(n356) );
  AND2_X1 U445 ( .A1(n625), .A2(n624), .ZN(n357) );
  AND2_X1 U446 ( .A1(n388), .A2(n371), .ZN(n358) );
  XNOR2_X1 U447 ( .A(KEYINPUT76), .B(KEYINPUT35), .ZN(n359) );
  NAND2_X1 U448 ( .A1(n743), .A2(n714), .ZN(n360) );
  XOR2_X1 U449 ( .A(n632), .B(n636), .Z(n361) );
  XNOR2_X1 U450 ( .A(KEYINPUT46), .B(KEYINPUT81), .ZN(n599) );
  INV_X1 U451 ( .A(n599), .ZN(n372) );
  XOR2_X1 U452 ( .A(KEYINPUT70), .B(KEYINPUT48), .Z(n362) );
  OR2_X1 U453 ( .A1(n613), .A2(n675), .ZN(n363) );
  XNOR2_X1 U454 ( .A(n552), .B(KEYINPUT45), .ZN(n614) );
  NAND2_X1 U455 ( .A1(n551), .A2(n550), .ZN(n552) );
  INV_X1 U456 ( .A(n374), .ZN(n386) );
  NAND2_X1 U457 ( .A1(n388), .A2(n387), .ZN(n374) );
  NAND2_X1 U458 ( .A1(n358), .A2(n384), .ZN(n383) );
  INV_X1 U459 ( .A(n387), .ZN(n373) );
  NAND2_X1 U460 ( .A1(n382), .A2(n374), .ZN(n381) );
  NAND2_X1 U461 ( .A1(n386), .A2(n384), .ZN(n752) );
  NAND2_X1 U462 ( .A1(n380), .A2(n375), .ZN(n600) );
  NAND2_X1 U463 ( .A1(n377), .A2(n599), .ZN(n376) );
  INV_X1 U464 ( .A(n750), .ZN(n377) );
  NAND2_X1 U465 ( .A1(n379), .A2(n382), .ZN(n378) );
  INV_X1 U466 ( .A(n384), .ZN(n379) );
  OR2_X1 U467 ( .A1(n665), .A2(KEYINPUT40), .ZN(n385) );
  NAND2_X1 U468 ( .A1(n603), .A2(KEYINPUT40), .ZN(n388) );
  NAND2_X1 U469 ( .A1(n396), .A2(n612), .ZN(n742) );
  XNOR2_X1 U470 ( .A(n602), .B(n362), .ZN(n396) );
  NAND2_X1 U471 ( .A1(n614), .A2(n553), .ZN(n398) );
  XNOR2_X2 U472 ( .A(n399), .B(n359), .ZN(n521) );
  NAND2_X2 U473 ( .A1(n400), .A2(n584), .ZN(n399) );
  XNOR2_X2 U474 ( .A(n402), .B(n401), .ZN(n400) );
  NAND2_X1 U475 ( .A1(n529), .A2(n696), .ZN(n402) );
  XNOR2_X1 U476 ( .A(n427), .B(n355), .ZN(n434) );
  INV_X1 U477 ( .A(KEYINPUT66), .ZN(n506) );
  XNOR2_X1 U478 ( .A(n484), .B(n429), .ZN(n740) );
  BUF_X1 U479 ( .A(n696), .Z(n712) );
  XNOR2_X1 U480 ( .A(n617), .B(n616), .ZN(n618) );
  INV_X1 U481 ( .A(n725), .ZN(n638) );
  XNOR2_X1 U482 ( .A(G131), .B(G134), .ZN(n403) );
  XNOR2_X1 U483 ( .A(n405), .B(n404), .ZN(n733) );
  INV_X1 U484 ( .A(KEYINPUT65), .ZN(n406) );
  XNOR2_X1 U485 ( .A(n733), .B(n354), .ZN(n457) );
  XOR2_X1 U486 ( .A(KEYINPUT5), .B(G137), .Z(n408) );
  NOR2_X1 U487 ( .A1(G953), .A2(G237), .ZN(n478) );
  NAND2_X1 U488 ( .A1(n478), .A2(G210), .ZN(n407) );
  XNOR2_X1 U489 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U490 ( .A(n457), .B(n409), .ZN(n410) );
  XNOR2_X1 U491 ( .A(n421), .B(n410), .ZN(n642) );
  OR2_X1 U492 ( .A1(n642), .A2(G902), .ZN(n413) );
  INV_X1 U493 ( .A(KEYINPUT99), .ZN(n411) );
  XNOR2_X1 U494 ( .A(n411), .B(G472), .ZN(n412) );
  XNOR2_X2 U495 ( .A(n413), .B(n412), .ZN(n688) );
  INV_X1 U496 ( .A(KEYINPUT6), .ZN(n414) );
  XNOR2_X1 U497 ( .A(n688), .B(n414), .ZN(n560) );
  XOR2_X1 U498 ( .A(G137), .B(G140), .Z(n429) );
  XOR2_X1 U499 ( .A(n454), .B(n415), .Z(n416) );
  XNOR2_X1 U500 ( .A(n429), .B(n416), .ZN(n419) );
  NAND2_X1 U501 ( .A1(G227), .A2(n743), .ZN(n417) );
  XNOR2_X2 U502 ( .A(G469), .B(n422), .ZN(n567) );
  INV_X1 U503 ( .A(KEYINPUT1), .ZN(n423) );
  NAND2_X1 U504 ( .A1(n502), .A2(G221), .ZN(n427) );
  XNOR2_X1 U505 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X2 U506 ( .A(n428), .B(G125), .ZN(n450) );
  XNOR2_X2 U507 ( .A(n450), .B(n353), .ZN(n484) );
  XOR2_X1 U508 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n431) );
  XNOR2_X1 U509 ( .A(G110), .B(KEYINPUT94), .ZN(n430) );
  XNOR2_X1 U510 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U511 ( .A(n740), .B(n432), .ZN(n433) );
  XNOR2_X1 U512 ( .A(n434), .B(n433), .ZN(n721) );
  XOR2_X1 U513 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n436) );
  XNOR2_X1 U514 ( .A(G902), .B(KEYINPUT15), .ZN(n613) );
  NAND2_X1 U515 ( .A1(G234), .A2(n613), .ZN(n435) );
  XNOR2_X1 U516 ( .A(n436), .B(n435), .ZN(n441) );
  NAND2_X1 U517 ( .A1(G217), .A2(n441), .ZN(n438) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n437) );
  XNOR2_X1 U519 ( .A(n438), .B(n437), .ZN(n439) );
  NAND2_X1 U520 ( .A1(n441), .A2(G221), .ZN(n443) );
  INV_X1 U521 ( .A(KEYINPUT21), .ZN(n442) );
  XNOR2_X1 U522 ( .A(n443), .B(n442), .ZN(n683) );
  XNOR2_X1 U523 ( .A(n683), .B(KEYINPUT97), .ZN(n510) );
  NOR2_X2 U524 ( .A1(n507), .A2(n510), .ZN(n527) );
  INV_X1 U525 ( .A(n527), .ZN(n680) );
  NOR2_X1 U526 ( .A1(n681), .A2(n680), .ZN(n535) );
  NAND2_X1 U527 ( .A1(n560), .A2(n535), .ZN(n446) );
  INV_X1 U528 ( .A(KEYINPUT109), .ZN(n444) );
  XNOR2_X1 U529 ( .A(n444), .B(KEYINPUT33), .ZN(n445) );
  XNOR2_X1 U530 ( .A(n446), .B(n445), .ZN(n696) );
  INV_X1 U531 ( .A(G953), .ZN(n447) );
  NAND2_X1 U532 ( .A1(n447), .A2(G224), .ZN(n448) );
  XNOR2_X1 U533 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U534 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U535 ( .A(n453), .B(n452), .ZN(n456) );
  XNOR2_X1 U536 ( .A(G122), .B(G104), .ZN(n487) );
  XNOR2_X1 U537 ( .A(n487), .B(KEYINPUT16), .ZN(n455) );
  XNOR2_X1 U538 ( .A(n455), .B(n454), .ZN(n734) );
  XNOR2_X1 U539 ( .A(n456), .B(n734), .ZN(n459) );
  INV_X1 U540 ( .A(n457), .ZN(n458) );
  XNOR2_X1 U541 ( .A(n459), .B(n458), .ZN(n632) );
  INV_X1 U542 ( .A(n613), .ZN(n553) );
  OR2_X2 U543 ( .A1(n632), .A2(n553), .ZN(n463) );
  INV_X1 U544 ( .A(G902), .ZN(n490) );
  INV_X1 U545 ( .A(G237), .ZN(n460) );
  NAND2_X1 U546 ( .A1(n490), .A2(n460), .ZN(n464) );
  NAND2_X1 U547 ( .A1(n464), .A2(G210), .ZN(n461) );
  XNOR2_X1 U548 ( .A(n461), .B(KEYINPUT87), .ZN(n462) );
  XNOR2_X2 U549 ( .A(n463), .B(n462), .ZN(n563) );
  NAND2_X1 U550 ( .A1(n464), .A2(G214), .ZN(n578) );
  NAND2_X1 U551 ( .A1(n563), .A2(n578), .ZN(n466) );
  INV_X1 U552 ( .A(KEYINPUT19), .ZN(n465) );
  XNOR2_X1 U553 ( .A(n466), .B(n465), .ZN(n570) );
  NAND2_X1 U554 ( .A1(G234), .A2(G237), .ZN(n467) );
  XNOR2_X1 U555 ( .A(n467), .B(KEYINPUT14), .ZN(n471) );
  NAND2_X1 U556 ( .A1(G952), .A2(n471), .ZN(n468) );
  XNOR2_X1 U557 ( .A(KEYINPUT88), .B(n468), .ZN(n710) );
  NOR2_X1 U558 ( .A1(G953), .A2(n710), .ZN(n470) );
  INV_X1 U559 ( .A(KEYINPUT89), .ZN(n469) );
  XNOR2_X1 U560 ( .A(n470), .B(n469), .ZN(n557) );
  NAND2_X1 U561 ( .A1(G902), .A2(n471), .ZN(n554) );
  XOR2_X1 U562 ( .A(KEYINPUT90), .B(G898), .Z(n729) );
  NAND2_X1 U563 ( .A1(G953), .A2(n729), .ZN(n736) );
  NOR2_X1 U564 ( .A1(n554), .A2(n736), .ZN(n472) );
  NOR2_X1 U565 ( .A1(n557), .A2(n472), .ZN(n473) );
  XOR2_X1 U566 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n477) );
  XNOR2_X1 U567 ( .A(G113), .B(G140), .ZN(n476) );
  XNOR2_X1 U568 ( .A(n477), .B(n476), .ZN(n482) );
  XOR2_X1 U569 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n480) );
  NAND2_X1 U570 ( .A1(G214), .A2(n478), .ZN(n479) );
  XNOR2_X1 U571 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U572 ( .A(n482), .B(n481), .Z(n483) );
  XNOR2_X1 U573 ( .A(n484), .B(n483), .ZN(n489) );
  XNOR2_X1 U574 ( .A(n485), .B(G131), .ZN(n486) );
  XNOR2_X1 U575 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U576 ( .A(n489), .B(n488), .ZN(n627) );
  NAND2_X1 U577 ( .A1(n627), .A2(n490), .ZN(n492) );
  XOR2_X1 U578 ( .A(KEYINPUT13), .B(G475), .Z(n491) );
  XNOR2_X1 U579 ( .A(n492), .B(n491), .ZN(n542) );
  XNOR2_X1 U580 ( .A(KEYINPUT106), .B(G478), .ZN(n505) );
  XNOR2_X1 U581 ( .A(n494), .B(n493), .ZN(n501) );
  XOR2_X1 U582 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n496) );
  XNOR2_X1 U583 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n495) );
  XNOR2_X1 U584 ( .A(n496), .B(n495), .ZN(n499) );
  XOR2_X1 U585 ( .A(KEYINPUT103), .B(n497), .Z(n498) );
  XNOR2_X1 U586 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U587 ( .A(n501), .B(n500), .Z(n504) );
  NAND2_X1 U588 ( .A1(G217), .A2(n502), .ZN(n503) );
  XNOR2_X1 U589 ( .A(n504), .B(n503), .ZN(n718) );
  XNOR2_X1 U590 ( .A(n505), .B(n356), .ZN(n540) );
  AND2_X1 U591 ( .A1(n542), .A2(n540), .ZN(n584) );
  XNOR2_X1 U592 ( .A(n521), .B(n506), .ZN(n518) );
  INV_X1 U593 ( .A(n507), .ZN(n562) );
  INV_X1 U594 ( .A(n681), .ZN(n544) );
  NAND2_X1 U595 ( .A1(n684), .A2(n544), .ZN(n508) );
  XNOR2_X1 U596 ( .A(n508), .B(KEYINPUT108), .ZN(n509) );
  OR2_X1 U597 ( .A1(n509), .A2(n560), .ZN(n514) );
  OR2_X1 U598 ( .A1(n542), .A2(n540), .ZN(n594) );
  NOR2_X1 U599 ( .A1(n594), .A2(n510), .ZN(n511) );
  NAND2_X1 U600 ( .A1(n534), .A2(n511), .ZN(n513) );
  XNOR2_X1 U601 ( .A(KEYINPUT72), .B(KEYINPUT22), .ZN(n512) );
  XNOR2_X1 U602 ( .A(n513), .B(n512), .ZN(n548) );
  OR2_X1 U603 ( .A1(n514), .A2(n548), .ZN(n515) );
  AND2_X1 U604 ( .A1(n684), .A2(n681), .ZN(n516) );
  INV_X1 U605 ( .A(n688), .ZN(n531) );
  NAND2_X1 U606 ( .A1(n516), .A2(n531), .ZN(n517) );
  OR2_X1 U607 ( .A1(n548), .A2(n517), .ZN(n624) );
  NAND2_X1 U608 ( .A1(n518), .A2(n357), .ZN(n520) );
  INV_X1 U609 ( .A(KEYINPUT44), .ZN(n519) );
  NAND2_X1 U610 ( .A1(n520), .A2(n519), .ZN(n526) );
  AND2_X1 U611 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n522) );
  AND2_X1 U612 ( .A1(n624), .A2(n522), .ZN(n523) );
  NAND2_X1 U613 ( .A1(n625), .A2(n523), .ZN(n524) );
  OR2_X1 U614 ( .A1(n521), .A2(n524), .ZN(n525) );
  NAND2_X1 U615 ( .A1(n526), .A2(n525), .ZN(n551) );
  INV_X1 U616 ( .A(n574), .ZN(n528) );
  NAND2_X1 U617 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U618 ( .A(KEYINPUT98), .B(n530), .Z(n532) );
  NAND2_X1 U619 ( .A1(n532), .A2(n531), .ZN(n533) );
  BUF_X1 U620 ( .A(n534), .Z(n537) );
  NAND2_X1 U621 ( .A1(n688), .A2(n535), .ZN(n693) );
  INV_X1 U622 ( .A(n693), .ZN(n536) );
  NAND2_X1 U623 ( .A1(n537), .A2(n536), .ZN(n539) );
  INV_X1 U624 ( .A(KEYINPUT31), .ZN(n538) );
  XNOR2_X1 U625 ( .A(n539), .B(n538), .ZN(n667) );
  NAND2_X1 U626 ( .A1(n654), .A2(n667), .ZN(n543) );
  INV_X1 U627 ( .A(n540), .ZN(n541) );
  NAND2_X1 U628 ( .A1(n542), .A2(n541), .ZN(n665) );
  OR2_X1 U629 ( .A1(n542), .A2(n541), .ZN(n668) );
  INV_X1 U630 ( .A(n668), .ZN(n657) );
  XNOR2_X1 U631 ( .A(KEYINPUT107), .B(n657), .ZN(n604) );
  NAND2_X1 U632 ( .A1(n665), .A2(n604), .ZN(n701) );
  NAND2_X1 U633 ( .A1(n543), .A2(n701), .ZN(n549) );
  NOR2_X1 U634 ( .A1(n684), .A2(n544), .ZN(n546) );
  INV_X1 U635 ( .A(n560), .ZN(n545) );
  NAND2_X1 U636 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U637 ( .A1(n548), .A2(n547), .ZN(n649) );
  AND2_X1 U638 ( .A1(n549), .A2(n649), .ZN(n550) );
  OR2_X1 U639 ( .A1(n743), .A2(n554), .ZN(n555) );
  NOR2_X1 U640 ( .A1(G900), .A2(n555), .ZN(n556) );
  OR2_X1 U641 ( .A1(n557), .A2(n556), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n575), .A2(n683), .ZN(n566) );
  INV_X1 U643 ( .A(n578), .ZN(n697) );
  OR2_X1 U644 ( .A1(n566), .A2(n697), .ZN(n558) );
  NOR2_X1 U645 ( .A1(n665), .A2(n558), .ZN(n559) );
  NAND2_X1 U646 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U647 ( .A1(n562), .A2(n561), .ZN(n605) );
  NAND2_X1 U648 ( .A1(n605), .A2(n590), .ZN(n564) );
  XNOR2_X1 U649 ( .A(n564), .B(KEYINPUT36), .ZN(n565) );
  NOR2_X1 U650 ( .A1(n681), .A2(n565), .ZN(n671) );
  XOR2_X1 U651 ( .A(KEYINPUT82), .B(n671), .Z(n589) );
  NAND2_X1 U652 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U653 ( .A(KEYINPUT113), .B(n569), .ZN(n596) );
  INV_X1 U654 ( .A(n596), .ZN(n572) );
  BUF_X1 U655 ( .A(n570), .Z(n571) );
  NOR2_X1 U656 ( .A1(n572), .A2(n571), .ZN(n663) );
  NAND2_X1 U657 ( .A1(n663), .A2(n701), .ZN(n573) );
  XNOR2_X1 U658 ( .A(KEYINPUT47), .B(n573), .ZN(n587) );
  XNOR2_X1 U659 ( .A(n574), .B(KEYINPUT111), .ZN(n576) );
  NAND2_X1 U660 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U661 ( .A(KEYINPUT74), .B(n577), .ZN(n581) );
  NAND2_X1 U662 ( .A1(n688), .A2(n578), .ZN(n579) );
  XNOR2_X1 U663 ( .A(KEYINPUT30), .B(n579), .ZN(n580) );
  XNOR2_X1 U664 ( .A(n582), .B(KEYINPUT73), .ZN(n591) );
  INV_X1 U665 ( .A(n590), .ZN(n607) );
  NOR2_X1 U666 ( .A1(n591), .A2(n607), .ZN(n583) );
  XNOR2_X1 U667 ( .A(n583), .B(KEYINPUT112), .ZN(n585) );
  NAND2_X1 U668 ( .A1(n585), .A2(n584), .ZN(n661) );
  INV_X1 U669 ( .A(n661), .ZN(n586) );
  NOR2_X1 U670 ( .A1(n587), .A2(n586), .ZN(n588) );
  AND2_X1 U671 ( .A1(n589), .A2(n588), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n590), .B(KEYINPUT38), .ZN(n698) );
  NOR2_X1 U673 ( .A1(n591), .A2(n698), .ZN(n593) );
  XOR2_X1 U674 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n592) );
  XOR2_X1 U675 ( .A(KEYINPUT115), .B(KEYINPUT42), .Z(n598) );
  INV_X1 U676 ( .A(n594), .ZN(n700) );
  NOR2_X1 U677 ( .A1(n698), .A2(n697), .ZN(n702) );
  AND2_X1 U678 ( .A1(n700), .A2(n702), .ZN(n595) );
  XOR2_X1 U679 ( .A(KEYINPUT41), .B(n595), .Z(n713) );
  NAND2_X1 U680 ( .A1(n713), .A2(n596), .ZN(n597) );
  NAND2_X1 U681 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n673) );
  NAND2_X1 U683 ( .A1(n681), .A2(n605), .ZN(n606) );
  XNOR2_X1 U684 ( .A(n606), .B(KEYINPUT43), .ZN(n608) );
  AND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n610) );
  INV_X1 U686 ( .A(KEYINPUT110), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n610), .B(n609), .ZN(n751) );
  INV_X1 U688 ( .A(n751), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n673), .A2(n611), .ZN(n612) );
  INV_X1 U690 ( .A(KEYINPUT2), .ZN(n675) );
  NAND2_X1 U691 ( .A1(n717), .A2(G469), .ZN(n619) );
  XOR2_X1 U692 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n615) );
  XNOR2_X1 U693 ( .A(n615), .B(KEYINPUT58), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n619), .B(n618), .ZN(n621) );
  INV_X1 U695 ( .A(G952), .ZN(n620) );
  NOR2_X2 U696 ( .A1(n621), .A2(n725), .ZN(n623) );
  INV_X1 U697 ( .A(KEYINPUT125), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(G54) );
  XNOR2_X1 U699 ( .A(n624), .B(G110), .ZN(G12) );
  XNOR2_X1 U700 ( .A(n625), .B(G119), .ZN(G21) );
  XOR2_X1 U701 ( .A(G122), .B(n521), .Z(G24) );
  NAND2_X1 U702 ( .A1(n717), .A2(G475), .ZN(n629) );
  XNOR2_X1 U703 ( .A(KEYINPUT64), .B(KEYINPUT59), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n629), .B(n628), .ZN(n630) );
  NOR2_X2 U706 ( .A1(n630), .A2(n725), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U708 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n633), .B(KEYINPUT78), .ZN(n635) );
  XNOR2_X1 U710 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n637), .B(n361), .ZN(n639) );
  XOR2_X1 U713 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n640) );
  XNOR2_X1 U714 ( .A(n641), .B(n640), .ZN(G51) );
  NAND2_X1 U715 ( .A1(n717), .A2(G472), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n642), .B(KEYINPUT62), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U718 ( .A(KEYINPUT116), .B(KEYINPUT63), .ZN(n646) );
  XOR2_X1 U719 ( .A(n646), .B(KEYINPUT86), .Z(n647) );
  XNOR2_X1 U720 ( .A(n648), .B(n647), .ZN(G57) );
  XNOR2_X1 U721 ( .A(G101), .B(n649), .ZN(G3) );
  NOR2_X1 U722 ( .A1(n654), .A2(n665), .ZN(n651) );
  XNOR2_X1 U723 ( .A(G104), .B(KEYINPUT117), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(G6) );
  XOR2_X1 U725 ( .A(KEYINPUT26), .B(KEYINPUT118), .Z(n653) );
  XNOR2_X1 U726 ( .A(G107), .B(KEYINPUT27), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(n656) );
  NOR2_X1 U728 ( .A1(n654), .A2(n668), .ZN(n655) );
  XOR2_X1 U729 ( .A(n656), .B(n655), .Z(G9) );
  XOR2_X1 U730 ( .A(KEYINPUT29), .B(KEYINPUT119), .Z(n659) );
  NAND2_X1 U731 ( .A1(n663), .A2(n657), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n659), .B(n658), .ZN(n660) );
  XOR2_X1 U733 ( .A(G128), .B(n660), .Z(G30) );
  XNOR2_X1 U734 ( .A(G143), .B(n661), .ZN(G45) );
  INV_X1 U735 ( .A(n665), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U737 ( .A(G146), .B(n664), .ZN(G48) );
  NOR2_X1 U738 ( .A1(n665), .A2(n667), .ZN(n666) );
  XOR2_X1 U739 ( .A(G113), .B(n666), .Z(G15) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U741 ( .A(KEYINPUT120), .B(n669), .Z(n670) );
  XNOR2_X1 U742 ( .A(G116), .B(n670), .ZN(G18) );
  XNOR2_X1 U743 ( .A(G125), .B(n671), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n672), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U745 ( .A(G134), .B(n673), .Z(G36) );
  XNOR2_X1 U746 ( .A(n674), .B(KEYINPUT79), .ZN(n677) );
  NAND2_X1 U747 ( .A1(n675), .A2(n742), .ZN(n676) );
  NAND2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U750 ( .A(KEYINPUT50), .B(n682), .ZN(n691) );
  XOR2_X1 U751 ( .A(KEYINPUT121), .B(KEYINPUT49), .Z(n687) );
  INV_X1 U752 ( .A(n683), .ZN(n685) );
  NAND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U754 ( .A(n687), .B(n686), .ZN(n689) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U758 ( .A(KEYINPUT51), .B(n694), .Z(n695) );
  NAND2_X1 U759 ( .A1(n713), .A2(n695), .ZN(n707) );
  NAND2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U762 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U764 ( .A1(n712), .A2(n705), .ZN(n706) );
  NAND2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U766 ( .A(KEYINPUT52), .B(n708), .Z(n709) );
  NOR2_X1 U767 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U768 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U769 ( .A(KEYINPUT122), .B(KEYINPUT53), .ZN(n715) );
  XNOR2_X1 U770 ( .A(n716), .B(n715), .ZN(G75) );
  NAND2_X1 U771 ( .A1(n717), .A2(G478), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n725), .A2(n720), .ZN(G63) );
  NAND2_X1 U774 ( .A1(n717), .A2(G217), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n721), .B(KEYINPUT126), .ZN(n722) );
  XNOR2_X1 U776 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U777 ( .A1(n725), .A2(n724), .ZN(G66) );
  NAND2_X1 U778 ( .A1(n726), .A2(n743), .ZN(n732) );
  NAND2_X1 U779 ( .A1(G953), .A2(G224), .ZN(n727) );
  XOR2_X1 U780 ( .A(KEYINPUT61), .B(n727), .Z(n728) );
  NOR2_X1 U781 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U782 ( .A(n730), .B(KEYINPUT127), .ZN(n731) );
  NAND2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n739) );
  XNOR2_X1 U784 ( .A(n733), .B(G101), .ZN(n735) );
  XNOR2_X1 U785 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U787 ( .A(n739), .B(n738), .Z(G69) );
  XOR2_X1 U788 ( .A(n741), .B(n740), .Z(n745) );
  XNOR2_X1 U789 ( .A(n742), .B(n745), .ZN(n744) );
  NAND2_X1 U790 ( .A1(n744), .A2(n743), .ZN(n749) );
  XNOR2_X1 U791 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U792 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U793 ( .A1(n747), .A2(G953), .ZN(n748) );
  NAND2_X1 U794 ( .A1(n749), .A2(n748), .ZN(G72) );
  XNOR2_X1 U795 ( .A(G137), .B(n750), .ZN(G39) );
  XNOR2_X1 U796 ( .A(G140), .B(n751), .ZN(G42) );
  XNOR2_X1 U797 ( .A(n752), .B(G131), .ZN(G33) );
endmodule

