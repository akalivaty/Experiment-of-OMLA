//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT88), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G8gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n204), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  AND2_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n218));
  XNOR2_X1  g017(.A(G43gat), .B(G50gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT17), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n209), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n204), .B(new_n207), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n221), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT18), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n225), .A2(KEYINPUT18), .A3(new_n226), .A4(new_n229), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n209), .A2(new_n223), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n229), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n226), .B(KEYINPUT13), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G197gat), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT11), .B(G169gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT12), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n232), .A2(new_n243), .A3(new_n233), .A4(new_n237), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(KEYINPUT89), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT89), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n238), .A2(new_n248), .A3(new_n244), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT91), .ZN(new_n252));
  NAND2_X1  g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT7), .ZN(new_n254));
  XNOR2_X1  g053(.A(G99gat), .B(G106gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(G99gat), .A2(G106gat), .ZN(new_n256));
  INV_X1    g055(.A(G85gat), .ZN(new_n257));
  INV_X1    g056(.A(G92gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(KEYINPUT8), .A2(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n254), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n255), .B1(new_n254), .B2(new_n259), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(KEYINPUT90), .A2(G57gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(G64gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(G71gat), .A2(G78gat), .ZN(new_n265));
  OR2_X1    g064(.A1(G71gat), .A2(G78gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT9), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n270));
  AND2_X1   g069(.A1(G57gat), .A2(G64gat), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n265), .B(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n262), .A2(KEYINPUT10), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n262), .A2(new_n274), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n273), .B1(new_n260), .B2(new_n261), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n252), .B(new_n275), .C1(new_n278), .C2(KEYINPUT10), .ZN(new_n279));
  NAND2_X1  g078(.A1(G230gat), .A2(G233gat), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n275), .A2(new_n252), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n280), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G120gat), .B(G148gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT93), .ZN(new_n287));
  XNOR2_X1  g086(.A(G176gat), .B(G204gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n284), .A2(KEYINPUT92), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(new_n289), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(KEYINPUT92), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n282), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT21), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n273), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G231gat), .A2(G233gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G127gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n209), .B1(new_n297), .B2(new_n273), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(G155gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(G183gat), .B(G211gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n308), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI221_X1 g110(.A(new_n222), .B1(new_n260), .B2(new_n261), .C1(new_n223), .C2(new_n224), .ZN(new_n312));
  XNOR2_X1  g111(.A(G190gat), .B(G218gat), .ZN(new_n313));
  AND2_X1   g112(.A1(G232gat), .A2(G233gat), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n228), .A2(new_n262), .B1(KEYINPUT41), .B2(new_n314), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n313), .B1(new_n312), .B2(new_n315), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n314), .A2(KEYINPUT41), .ZN(new_n318));
  XNOR2_X1  g117(.A(G134gat), .B(G162gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OR3_X1    g120(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n316), .B2(new_n317), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n251), .A2(new_n296), .A3(new_n311), .A4(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n301), .A2(G134gat), .ZN(new_n328));
  INV_X1    g127(.A(G134gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G127gat), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n327), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT67), .B1(new_n301), .B2(G134gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n331), .A2(new_n332), .B1(KEYINPUT1), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G141gat), .B(G148gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(G155gat), .B2(G162gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G141gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G148gat), .ZN(new_n343));
  INV_X1    g142(.A(G148gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G141gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G155gat), .B(G162gat), .ZN(new_n347));
  INV_X1    g146(.A(G155gat), .ZN(new_n348));
  INV_X1    g147(.A(G162gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT2), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n329), .A2(G127gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n301), .A2(G134gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G120gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G113gat), .ZN(new_n356));
  INV_X1    g155(.A(G113gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G120gat), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT1), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n334), .A2(new_n341), .A3(new_n351), .A4(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n326), .B1(new_n361), .B2(KEYINPUT4), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT67), .B1(new_n352), .B2(new_n353), .ZN(new_n363));
  INV_X1    g162(.A(new_n332), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n359), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n328), .A2(new_n330), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n366), .A2(new_n333), .A3(KEYINPUT1), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n341), .A2(new_n351), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n368), .A2(KEYINPUT74), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n362), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n341), .A2(new_n351), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n341), .A2(new_n351), .A3(KEYINPUT73), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(KEYINPUT3), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n332), .B1(new_n366), .B2(KEYINPUT67), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n360), .B1(new_n381), .B2(new_n359), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n341), .A2(new_n351), .A3(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n375), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n373), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n361), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n390), .B2(new_n375), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n387), .A2(KEYINPUT75), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT75), .B1(new_n387), .B2(new_n391), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n370), .A2(new_n369), .A3(new_n334), .A4(new_n360), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n372), .A2(new_n394), .A3(KEYINPUT77), .ZN(new_n395));
  OR3_X1    g194(.A1(new_n361), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT5), .B(new_n375), .C1(new_n380), .C2(new_n385), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT78), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n396), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n341), .A2(new_n351), .A3(KEYINPUT73), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT73), .B1(new_n341), .B2(new_n351), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n401), .A2(new_n402), .A3(new_n383), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n382), .A2(new_n384), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n388), .B(new_n374), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT78), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n400), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n392), .A2(new_n393), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(G1gat), .B(G29gat), .Z(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n408), .A2(KEYINPUT6), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n387), .A2(new_n391), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT75), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n387), .A2(KEYINPUT75), .A3(new_n391), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n406), .B1(new_n400), .B2(new_n405), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n397), .A2(KEYINPUT78), .A3(new_n398), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n419), .A2(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n416), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n421), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n425), .B(new_n413), .C1(new_n393), .C2(new_n392), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n415), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT72), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT65), .ZN(new_n431));
  NAND2_X1  g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(G169gat), .A2(G176gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n432), .B1(new_n433), .B2(KEYINPUT23), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT23), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n435), .A2(G169gat), .A3(G176gat), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n431), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT24), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n438), .A2(G183gat), .A3(G190gat), .ZN(new_n439));
  INV_X1    g238(.A(G183gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G190gat), .ZN(new_n441));
  INV_X1    g240(.A(G190gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G183gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n439), .B1(new_n444), .B2(KEYINPUT24), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n433), .A2(KEYINPUT23), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n435), .B1(G169gat), .B2(G176gat), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n446), .A2(KEYINPUT65), .A3(new_n447), .A4(new_n432), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n437), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n450));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n436), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n438), .B1(new_n441), .B2(new_n443), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT25), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n452), .A2(new_n453), .A3(new_n439), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n449), .A2(new_n450), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n433), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n456));
  INV_X1    g255(.A(G169gat), .ZN(new_n457));
  INV_X1    g256(.A(G176gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n456), .A2(new_n461), .A3(KEYINPUT66), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT27), .B(G183gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT28), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n442), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n440), .A2(KEYINPUT27), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G183gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n471), .A3(new_n442), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT28), .ZN(new_n473));
  AND4_X1   g272(.A1(new_n464), .A2(new_n465), .A3(new_n468), .A4(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n430), .B1(new_n455), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G226gat), .ZN(new_n476));
  INV_X1    g275(.A(G233gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n449), .A2(new_n450), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n454), .A2(new_n451), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n465), .A2(new_n473), .A3(new_n468), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n464), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n481), .B1(new_n487), .B2(new_n478), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n481), .B(new_n478), .C1(new_n455), .C2(new_n474), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n480), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G211gat), .A2(G218gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT22), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(G197gat), .A2(G204gat), .ZN(new_n495));
  AND2_X1   g294(.A1(G197gat), .A2(G204gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G211gat), .ZN(new_n498));
  INV_X1    g297(.A(G218gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n492), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n492), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(new_n494), .C1(new_n495), .C2(new_n496), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n491), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n478), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n480), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  XOR2_X1   g307(.A(G8gat), .B(G36gat), .Z(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT70), .ZN(new_n510));
  XNOR2_X1  g309(.A(G64gat), .B(G92gat), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n510), .B(new_n511), .Z(new_n512));
  NAND4_X1  g311(.A1(new_n506), .A2(KEYINPUT30), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n512), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n482), .A2(new_n483), .B1(new_n464), .B2(new_n485), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT69), .B1(new_n515), .B2(new_n479), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n489), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n504), .B1(new_n517), .B2(new_n480), .ZN(new_n518));
  INV_X1    g317(.A(new_n508), .ZN(new_n519));
  OAI211_X1 g318(.A(KEYINPUT71), .B(new_n514), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n516), .A2(new_n489), .B1(new_n479), .B2(new_n475), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n508), .B1(new_n522), .B2(new_n504), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT71), .B1(new_n523), .B2(new_n514), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n429), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n514), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT71), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n528), .A2(KEYINPUT72), .A3(new_n513), .A4(new_n520), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n508), .B(new_n512), .C1(new_n522), .C2(new_n504), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n428), .A2(new_n525), .A3(new_n529), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT79), .ZN(new_n534));
  INV_X1    g333(.A(new_n532), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n408), .A2(new_n414), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(new_n416), .A3(new_n426), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n535), .B1(new_n537), .B2(new_n415), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT79), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n538), .A2(new_n539), .A3(new_n525), .A4(new_n529), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n541));
  NAND2_X1  g340(.A1(G228gat), .A2(G233gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n504), .B1(new_n384), .B2(new_n430), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT3), .B1(new_n504), .B2(new_n430), .ZN(new_n544));
  OAI22_X1  g343(.A1(new_n543), .A2(KEYINPUT80), .B1(new_n544), .B2(new_n370), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n384), .A2(new_n430), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n546), .A2(KEYINPUT80), .A3(new_n505), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n542), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT81), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT81), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n550), .B(new_n542), .C1(new_n545), .C2(new_n547), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n544), .A2(new_n401), .A3(new_n402), .ZN(new_n553));
  NOR3_X1   g352(.A1(new_n553), .A2(new_n542), .A3(new_n543), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(KEYINPUT31), .B(G50gat), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G78gat), .B(G106gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G22gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n557), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n552), .A2(new_n561), .A3(new_n555), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n560), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n561), .B1(new_n552), .B2(new_n555), .ZN(new_n565));
  AOI211_X1 g364(.A(new_n557), .B(new_n554), .C1(new_n549), .C2(new_n551), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n484), .A2(new_n486), .A3(new_n382), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n368), .B1(new_n455), .B2(new_n474), .ZN(new_n571));
  INV_X1    g370(.A(G227gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(new_n477), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT68), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n570), .A2(new_n571), .A3(new_n576), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n570), .A2(new_n571), .ZN(new_n581));
  INV_X1    g380(.A(new_n573), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT34), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT34), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G15gat), .B(G43gat), .Z(new_n588));
  XNOR2_X1  g387(.A(G71gat), .B(G99gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n580), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n578), .A2(KEYINPUT32), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n585), .B1(new_n581), .B2(new_n582), .ZN(new_n594));
  AOI211_X1 g393(.A(KEYINPUT34), .B(new_n573), .C1(new_n570), .C2(new_n571), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT33), .B1(new_n575), .B2(new_n577), .ZN(new_n597));
  INV_X1    g396(.A(new_n590), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n591), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n593), .B1(new_n591), .B2(new_n599), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n541), .B1(new_n569), .B2(new_n602), .ZN(new_n603));
  NOR4_X1   g402(.A1(new_n568), .A2(new_n600), .A3(new_n601), .A4(KEYINPUT86), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n534), .B(new_n540), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT35), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT84), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n415), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n408), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n414), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n537), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n528), .A2(new_n513), .A3(new_n520), .A4(new_n532), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT85), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT85), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n610), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n602), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n618), .A2(KEYINPUT35), .A3(new_n568), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n606), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n534), .A2(new_n540), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n568), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT37), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n512), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n523), .B2(new_n514), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n506), .B2(new_n508), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT38), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n608), .A2(new_n628), .A3(new_n609), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n480), .A2(new_n507), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n624), .B1(new_n630), .B2(new_n505), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n491), .A2(new_n504), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT38), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n512), .B1(new_n506), .B2(new_n508), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n625), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n537), .A2(new_n530), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n569), .B1(new_n629), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT83), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n380), .A2(new_n385), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n395), .A2(new_n396), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n375), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n390), .A2(new_n375), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n640), .A2(new_n643), .A3(new_n375), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n413), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT82), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT82), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n651), .A3(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n645), .A2(KEYINPUT40), .A3(new_n413), .A4(new_n646), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n423), .B2(new_n413), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AND4_X1   g455(.A1(new_n638), .A2(new_n611), .A3(new_n653), .A4(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n650), .B2(new_n652), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n638), .B1(new_n658), .B2(new_n611), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n637), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT36), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n600), .B2(new_n601), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n591), .A2(new_n599), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n592), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n591), .A2(new_n593), .A3(new_n599), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(KEYINPUT36), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n623), .A2(new_n660), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n325), .B1(new_n621), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n428), .B(KEYINPUT94), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n611), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT16), .B(G8gat), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT95), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n674), .A2(G8gat), .ZN(new_n681));
  OAI22_X1  g480(.A1(new_n681), .A2(new_n675), .B1(new_n674), .B2(new_n676), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n679), .B1(new_n680), .B2(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(KEYINPUT96), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n600), .A2(new_n601), .A3(new_n661), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT36), .B1(new_n664), .B2(new_n665), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n662), .A2(new_n666), .A3(KEYINPUT96), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT97), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n669), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n618), .A2(G15gat), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n691), .A2(G15gat), .B1(new_n669), .B2(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT98), .Z(G1326gat));
  NAND2_X1  g493(.A1(new_n669), .A2(new_n568), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT99), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  AOI21_X1  g497(.A(new_n324), .B1(new_n621), .B2(new_n668), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n250), .A2(new_n311), .A3(new_n295), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(G29gat), .A3(new_n670), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT45), .Z(new_n703));
  INV_X1    g502(.A(new_n324), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n569), .B1(new_n534), .B2(new_n540), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n637), .A2(new_n657), .A3(new_n659), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n706), .A2(new_n707), .A3(new_n689), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n605), .A2(KEYINPUT35), .B1(new_n617), .B2(new_n619), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n704), .B(new_n705), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n699), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n700), .B(KEYINPUT100), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n714), .B2(new_n670), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n703), .A2(new_n715), .ZN(G1328gat));
  AND2_X1   g515(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n701), .A2(G36gat), .A3(new_n612), .ZN(new_n720));
  MUX2_X1   g519(.A(new_n719), .B(new_n717), .S(new_n720), .Z(new_n721));
  OAI21_X1  g520(.A(G36gat), .B1(new_n714), .B2(new_n612), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1329gat));
  NOR3_X1   g522(.A1(new_n701), .A2(G43gat), .A3(new_n618), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n712), .A2(new_n713), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n690), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n726), .B2(G43gat), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(G43gat), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n725), .B2(new_n689), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n727), .A2(KEYINPUT47), .B1(new_n729), .B2(new_n731), .ZN(G1330gat));
  INV_X1    g531(.A(G50gat), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n725), .B2(new_n568), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n701), .A2(G50gat), .A3(new_n569), .ZN(new_n736));
  OR3_X1    g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(KEYINPUT104), .ZN(new_n738));
  OAI21_X1  g537(.A(G50gat), .B1(new_n714), .B2(new_n569), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT103), .B(KEYINPUT48), .Z(new_n743));
  OAI21_X1  g542(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(G1331gat));
  NAND3_X1  g543(.A1(new_n250), .A2(new_n311), .A3(new_n324), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n687), .A2(new_n688), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n623), .A2(new_n660), .A3(new_n746), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n296), .B(new_n745), .C1(new_n621), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n671), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT105), .B(G57gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1332gat));
  OR2_X1    g550(.A1(new_n611), .A2(KEYINPUT106), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n611), .A2(KEYINPUT106), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n748), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT107), .Z(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1333gat));
  NAND2_X1  g559(.A1(new_n748), .A2(new_n690), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n618), .A2(G71gat), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n761), .A2(G71gat), .B1(new_n748), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n568), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n251), .A2(new_n311), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n296), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n712), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n670), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n704), .B(new_n767), .C1(new_n708), .C2(new_n709), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n621), .A2(new_n747), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n704), .A4(new_n767), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n671), .A2(new_n257), .A3(new_n295), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n771), .B1(new_n778), .B2(new_n779), .ZN(G1336gat));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n776), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n755), .A2(G92gat), .A3(new_n296), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n712), .A2(new_n611), .A3(new_n769), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n786), .A2(KEYINPUT109), .B1(new_n787), .B2(G92gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n785), .ZN(new_n789));
  AOI211_X1 g588(.A(KEYINPUT109), .B(new_n789), .C1(new_n783), .C2(new_n776), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n781), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G92gat), .B1(new_n770), .B2(new_n755), .ZN(new_n793));
  XOR2_X1   g592(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n777), .B2(new_n785), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT111), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n799));
  INV_X1    g598(.A(new_n769), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n623), .A2(new_n660), .A3(new_n667), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n704), .B1(new_n801), .B2(new_n709), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT44), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n800), .B1(new_n803), .B2(new_n710), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n258), .B1(new_n804), .B2(new_n611), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n784), .B2(new_n785), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n805), .A2(new_n790), .A3(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n799), .B(new_n796), .C1(new_n808), .C2(new_n781), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n798), .A2(new_n809), .ZN(G1337gat));
  INV_X1    g609(.A(G99gat), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n777), .A2(new_n811), .A3(new_n602), .A4(new_n295), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n804), .A2(new_n690), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n813), .B2(new_n811), .ZN(G1338gat));
  OAI21_X1  g613(.A(G106gat), .B1(new_n770), .B2(new_n569), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n569), .A2(G106gat), .A3(new_n296), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT53), .B1(new_n777), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n784), .A2(new_n816), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n820), .A2(KEYINPUT112), .A3(KEYINPUT53), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT112), .B1(new_n820), .B2(KEYINPUT53), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(G1339gat));
  INV_X1    g622(.A(new_n311), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n235), .A2(new_n236), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n226), .B1(new_n225), .B2(new_n229), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n242), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n322), .A2(new_n246), .A3(new_n323), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n279), .A2(new_n281), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n283), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(KEYINPUT54), .A3(new_n282), .ZN(new_n832));
  XNOR2_X1  g631(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n279), .A2(new_n281), .A3(new_n280), .A4(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n289), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n835), .A3(KEYINPUT55), .ZN(new_n836));
  INV_X1    g635(.A(new_n294), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n835), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n829), .A2(KEYINPUT114), .A3(new_n836), .A4(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n839), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n294), .A3(new_n836), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n844), .B2(new_n828), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n247), .A2(new_n840), .A3(new_n249), .A4(new_n836), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n246), .A2(new_n827), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n295), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n704), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n824), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n745), .A2(new_n295), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT115), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n851), .A2(new_n856), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n670), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n603), .A2(new_n604), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n859), .A2(new_n860), .A3(new_n755), .ZN(new_n861));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n251), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n858), .A2(new_n568), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(new_n671), .A3(new_n602), .A4(new_n755), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n357), .A3(new_n250), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n862), .A2(new_n865), .ZN(G1340gat));
  AOI21_X1  g665(.A(G120gat), .B1(new_n861), .B2(new_n295), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n864), .A2(new_n355), .A3(new_n296), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  NAND3_X1  g668(.A1(new_n861), .A2(new_n301), .A3(new_n311), .ZN(new_n870));
  OAI21_X1  g669(.A(G127gat), .B1(new_n864), .B2(new_n824), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  NOR2_X1   g671(.A1(new_n611), .A2(new_n324), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n859), .A2(new_n329), .A3(new_n860), .A4(new_n873), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n864), .B2(new_n324), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  NOR3_X1   g677(.A1(new_n689), .A2(new_n670), .A3(new_n754), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n855), .A2(new_n568), .A3(new_n857), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n569), .A2(new_n882), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n844), .A2(KEYINPUT117), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n840), .B2(new_n836), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n885), .A2(new_n250), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n849), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n324), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n846), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n311), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n884), .B1(new_n892), .B2(new_n852), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(KEYINPUT118), .B(new_n884), .C1(new_n892), .C2(new_n852), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n883), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n251), .B(new_n879), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G141gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n690), .A2(new_n569), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n859), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n902), .A2(new_n342), .A3(new_n251), .A4(new_n755), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT58), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n900), .B(new_n903), .C1(new_n905), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1344gat));
  NAND2_X1  g709(.A1(new_n902), .A2(new_n755), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(G148gat), .A3(new_n296), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT120), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n879), .B1(new_n897), .B2(new_n898), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n914), .B(G148gat), .C1(new_n915), .C2(new_n296), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n829), .A2(new_n836), .A3(new_n840), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n311), .B1(new_n890), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n852), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(KEYINPUT57), .A3(new_n569), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(KEYINPUT57), .B2(new_n880), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n295), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n344), .B1(new_n922), .B2(new_n879), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n916), .B1(new_n923), .B2(new_n914), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n913), .A2(new_n924), .ZN(G1345gat));
  OAI21_X1  g724(.A(G155gat), .B1(new_n915), .B2(new_n824), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n902), .A2(new_n348), .A3(new_n311), .A4(new_n755), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(KEYINPUT121), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1346gat));
  OAI21_X1  g731(.A(G162gat), .B1(new_n915), .B2(new_n324), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n902), .A2(new_n349), .A3(new_n873), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1347gat));
  NAND4_X1  g734(.A1(new_n863), .A2(new_n670), .A3(new_n611), .A4(new_n602), .ZN(new_n936));
  OAI21_X1  g735(.A(G169gat), .B1(new_n936), .B2(new_n250), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT123), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n858), .A2(new_n671), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n860), .A2(new_n754), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT122), .Z(new_n941));
  AND2_X1   g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n457), .A3(new_n251), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n938), .A2(new_n943), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n936), .B2(new_n296), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n942), .A2(new_n458), .A3(new_n295), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1349gat));
  OAI21_X1  g746(.A(G183gat), .B1(new_n936), .B2(new_n824), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n466), .A3(new_n311), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n942), .A2(new_n442), .A3(new_n704), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n936), .A2(new_n324), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n954), .A4(G190gat), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n442), .B1(new_n957), .B2(KEYINPUT61), .ZN(new_n958));
  AOI22_X1  g757(.A1(new_n953), .A2(new_n958), .B1(KEYINPUT124), .B2(new_n954), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n952), .B1(new_n956), .B2(new_n959), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n690), .A2(new_n671), .A3(new_n612), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n921), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(G197gat), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n962), .A2(new_n963), .A3(new_n250), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n939), .A2(new_n754), .A3(new_n901), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(G197gat), .B1(new_n966), .B2(new_n251), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n964), .A2(new_n967), .ZN(G1352gat));
  NAND2_X1  g767(.A1(new_n922), .A2(new_n961), .ZN(new_n969));
  XNOR2_X1  g768(.A(KEYINPUT125), .B(G204gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n965), .A2(new_n296), .A3(new_n970), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1353gat));
  NAND3_X1  g773(.A1(new_n966), .A2(new_n498), .A3(new_n311), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n921), .A2(new_n311), .A3(new_n961), .ZN(new_n977));
  AND4_X1   g776(.A1(new_n976), .A2(new_n977), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(G211gat), .B1(new_n976), .B2(KEYINPUT63), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AOI22_X1  g779(.A1(new_n977), .A2(new_n980), .B1(new_n976), .B2(KEYINPUT63), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n975), .B1(new_n978), .B2(new_n981), .ZN(G1354gat));
  OAI21_X1  g781(.A(new_n499), .B1(new_n965), .B2(new_n324), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT127), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n962), .A2(new_n499), .A3(new_n324), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n984), .A2(new_n985), .ZN(G1355gat));
endmodule


