//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT64), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(new_n188), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n191), .A2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n189), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n187), .A2(new_n198), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n194), .A2(new_n197), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  OAI22_X1  g021(.A1(new_n198), .A2(new_n199), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n190), .A2(new_n192), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n205), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G224), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G953), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n205), .B(new_n212), .C1(new_n214), .C2(G953), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G113), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G119), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT65), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G116), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n225), .A2(G119), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n223), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n220), .A2(new_n222), .ZN(new_n233));
  INV_X1    g047(.A(new_n230), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT65), .B(G116), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n233), .B(new_n234), .C1(new_n235), .C2(new_n224), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n231), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n235), .B2(new_n224), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT66), .A3(new_n223), .ZN(new_n239));
  INV_X1    g053(.A(G104), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT3), .B1(new_n240), .B2(G107), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n242));
  INV_X1    g056(.A(G107), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(G104), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(G107), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G101), .ZN(new_n247));
  INV_X1    g061(.A(G101), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n241), .A2(new_n244), .A3(new_n248), .A4(new_n245), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n251), .A3(G101), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n237), .A2(new_n239), .A3(new_n250), .A4(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n234), .B(new_n254), .C1(new_n235), .C2(new_n224), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT88), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT88), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n219), .B1(new_n260), .B2(new_n230), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n243), .A2(G104), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n240), .A2(G107), .ZN(new_n264));
  OAI21_X1  g078(.A(G101), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n249), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n249), .B2(new_n265), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n236), .B(new_n262), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n253), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(G110), .B(G122), .Z(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n273));
  INV_X1    g087(.A(new_n271), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n253), .A2(new_n274), .A3(new_n269), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT6), .A4(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n253), .A2(new_n274), .A3(new_n269), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n274), .B1(new_n253), .B2(new_n269), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT89), .B1(new_n278), .B2(new_n279), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n218), .B(new_n276), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT90), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n273), .B1(new_n272), .B2(KEYINPUT6), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n272), .A2(KEYINPUT6), .A3(new_n275), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT90), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n218), .A4(new_n276), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n261), .B1(new_n238), .B2(new_n256), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n290), .B(new_n236), .C1(new_n267), .C2(new_n268), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT91), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n249), .A2(new_n265), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT83), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n249), .A2(new_n265), .A3(new_n266), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(KEYINPUT91), .A3(new_n236), .A4(new_n290), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n262), .A2(new_n236), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n294), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(new_n271), .B(KEYINPUT8), .Z(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n216), .B(new_n217), .C1(KEYINPUT7), .C2(new_n215), .ZN(new_n304));
  OR3_X1    g118(.A1(new_n213), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n303), .A2(new_n275), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n289), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n308), .B1(new_n283), .B2(new_n288), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n311), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(KEYINPUT92), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G214), .B1(G237), .B2(G902), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n314), .A2(KEYINPUT92), .A3(new_n311), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G475), .ZN(new_n321));
  NOR2_X1   g135(.A1(KEYINPUT93), .A2(G143), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(G237), .A2(G953), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(G214), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(G214), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n322), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G131), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT17), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT95), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(G125), .A2(G140), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(G125), .A2(G140), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT16), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(new_n189), .ZN(new_n338));
  AOI21_X1  g152(.A(G146), .B1(new_n335), .B2(new_n336), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G131), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n325), .A2(new_n327), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n329), .A2(new_n330), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT95), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n328), .A2(new_n344), .A3(KEYINPUT17), .A4(G131), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n331), .A2(new_n340), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G113), .B(G122), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(new_n240), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n328), .A2(KEYINPUT18), .A3(G131), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n333), .B2(new_n334), .ZN(new_n351));
  INV_X1    g165(.A(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n204), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT78), .A3(new_n332), .ZN(new_n354));
  AOI21_X1  g168(.A(G146), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n332), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(new_n189), .ZN(new_n357));
  AND2_X1   g171(.A1(KEYINPUT18), .A2(G131), .ZN(new_n358));
  OAI221_X1 g172(.A(new_n349), .B1(new_n355), .B2(new_n357), .C1(new_n328), .C2(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n346), .A2(new_n348), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n348), .B1(new_n346), .B2(new_n359), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n321), .B1(new_n362), .B2(new_n307), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT19), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n365), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n356), .A2(new_n366), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n351), .A2(new_n354), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n366), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n189), .B(new_n367), .C1(new_n370), .C2(new_n365), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n338), .B1(new_n329), .B2(new_n342), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n348), .B1(new_n373), .B2(new_n359), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n321), .B(new_n307), .C1(new_n360), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT20), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT96), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(KEYINPUT20), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n375), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n364), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G952), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(G953), .ZN(new_n383));
  INV_X1    g197(.A(G234), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G953), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT74), .B(G902), .Z(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI211_X1 g204(.A(new_n388), .B(new_n390), .C1(G234), .C2(G237), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT21), .B(G898), .Z(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n387), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT98), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT15), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G478), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G128), .B(G143), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT13), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n191), .A2(G128), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n400), .B(G134), .C1(KEYINPUT13), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G134), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n226), .A2(new_n228), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G122), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n225), .A2(G122), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n243), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G122), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n226), .B2(new_n228), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n411), .A2(G107), .A3(new_n407), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n402), .B(new_n404), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n414), .B(new_n408), .C1(new_n235), .C2(new_n410), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(G107), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n406), .A2(new_n243), .A3(new_n408), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n399), .B(new_n403), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT9), .B(G234), .ZN(new_n421));
  INV_X1    g235(.A(G217), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n421), .A2(new_n422), .A3(G953), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n413), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n413), .B2(new_n420), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n390), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT97), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n398), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n427), .ZN(new_n430));
  OAI211_X1 g244(.A(KEYINPUT97), .B(new_n390), .C1(new_n424), .C2(new_n425), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n395), .B(new_n429), .C1(new_n432), .C2(new_n397), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n397), .B1(new_n430), .B2(new_n431), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT98), .B1(new_n434), .B2(new_n428), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n381), .A2(new_n394), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G221), .ZN(new_n438));
  INV_X1    g252(.A(new_n421), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(new_n307), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT11), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n403), .B2(G137), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n403), .A2(G137), .ZN(new_n443));
  INV_X1    g257(.A(G137), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT11), .A3(G134), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G131), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n442), .A2(new_n445), .A3(new_n341), .A4(new_n443), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT10), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n249), .A2(new_n265), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n203), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n203), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n297), .A2(KEYINPUT10), .A3(new_n203), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT67), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n206), .A2(new_n207), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n210), .B(new_n459), .C1(new_n460), .C2(new_n195), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n208), .B2(new_n210), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n250), .B(new_n252), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n450), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n456), .A2(new_n450), .A3(new_n464), .A4(new_n457), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n388), .A2(G227), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(G140), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT81), .B(G110), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n203), .A2(new_n452), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT82), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n203), .A2(new_n452), .A3(new_n453), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n297), .B2(new_n203), .ZN(new_n478));
  INV_X1    g292(.A(new_n203), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n479), .A2(new_n295), .A3(KEYINPUT85), .A4(new_n296), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n449), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT12), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n481), .A2(new_n482), .A3(new_n485), .A4(new_n449), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n466), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n470), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n472), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G469), .B1(new_n489), .B2(G902), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n471), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n466), .A2(KEYINPUT87), .A3(new_n470), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n492), .A2(new_n484), .A3(new_n486), .A4(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n466), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n488), .B1(new_n465), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT86), .A2(G469), .ZN(new_n498));
  OR2_X1    g312(.A1(KEYINPUT86), .A2(G469), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n497), .A2(new_n390), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n440), .B1(new_n490), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n437), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n320), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n369), .A2(new_n189), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n224), .A2(G128), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n224), .A2(G128), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(KEYINPUT77), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(KEYINPUT77), .B2(new_n505), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT24), .B(G110), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n506), .A2(KEYINPUT23), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(KEYINPUT23), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n505), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(G110), .ZN(new_n514));
  OAI221_X1 g328(.A(new_n504), .B1(new_n189), .B2(new_n337), .C1(new_n510), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(G110), .ZN(new_n516));
  OAI221_X1 g330(.A(new_n516), .B1(new_n508), .B2(new_n509), .C1(new_n339), .C2(new_n338), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n438), .A2(new_n384), .A3(G953), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n519), .B(new_n520), .Z(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n515), .A2(new_n517), .A3(new_n521), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n422), .B1(new_n390), .B2(G234), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(G902), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT80), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AND4_X1   g342(.A1(KEYINPUT80), .A2(new_n523), .A3(new_n524), .A4(new_n527), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n523), .A2(new_n524), .ZN(new_n531));
  OAI22_X1  g345(.A1(new_n531), .A2(new_n389), .B1(KEYINPUT79), .B2(KEYINPUT25), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n526), .A2(KEYINPUT76), .ZN(new_n533));
  NOR2_X1   g347(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n523), .A2(new_n390), .A3(new_n534), .A4(new_n524), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n526), .A2(KEYINPUT76), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n532), .A2(new_n533), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n324), .A2(G210), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT29), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n237), .A2(new_n239), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n449), .B1(new_n462), .B2(new_n463), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n444), .A2(G134), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n403), .A2(G137), .ZN(new_n550));
  OAI21_X1  g364(.A(G131), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n448), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n203), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT28), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT73), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n548), .A2(new_n553), .ZN(new_n558));
  INV_X1    g372(.A(new_n547), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(KEYINPUT71), .A3(new_n554), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n547), .A2(new_n548), .A3(new_n562), .A4(new_n553), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(KEYINPUT28), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT72), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n561), .A2(new_n563), .A3(KEYINPUT72), .A4(KEYINPUT28), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n546), .B(new_n557), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n540), .B1(new_n568), .B2(new_n389), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n557), .B1(new_n566), .B2(new_n567), .ZN(new_n570));
  INV_X1    g384(.A(new_n546), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(KEYINPUT75), .A3(new_n390), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT30), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n203), .A2(new_n552), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n447), .A2(new_n448), .B1(new_n208), .B2(new_n210), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n548), .A2(KEYINPUT30), .A3(new_n553), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n559), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n554), .ZN(new_n580));
  INV_X1    g394(.A(new_n545), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT29), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT69), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n559), .B(new_n583), .C1(new_n575), .C2(new_n576), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n554), .A2(KEYINPUT69), .ZN(new_n585));
  INV_X1    g399(.A(new_n576), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n547), .B1(new_n553), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n584), .B(KEYINPUT28), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n556), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n582), .B1(new_n589), .B2(new_n581), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n569), .A2(new_n573), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NOR2_X1   g406(.A1(G472), .A2(G902), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT70), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n579), .A2(new_n545), .A3(new_n554), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT31), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT31), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n579), .A2(new_n597), .A3(new_n545), .A4(new_n554), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n589), .A2(new_n581), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n594), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n598), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n545), .B1(new_n588), .B2(new_n556), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT70), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n593), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT32), .ZN(new_n606));
  INV_X1    g420(.A(new_n593), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n600), .A2(new_n594), .A3(new_n598), .A4(new_n596), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT70), .B1(new_n602), .B2(new_n603), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT32), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n539), .B1(new_n592), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n503), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  NAND2_X1  g430(.A1(new_n490), .A2(new_n500), .ZN(new_n617));
  INV_X1    g431(.A(new_n440), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(G472), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n389), .B1(new_n608), .B2(new_n609), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n605), .B(new_n538), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n311), .B1(new_n289), .B2(new_n309), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n312), .B(new_n308), .C1(new_n283), .C2(new_n288), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n317), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n424), .A2(new_n425), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT33), .Z(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(G478), .A3(new_n390), .ZN(new_n629));
  INV_X1    g443(.A(new_n426), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n629), .B1(G478), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n381), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n626), .A2(new_n632), .A3(new_n394), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n638));
  INV_X1    g452(.A(new_n394), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n375), .A2(KEYINPUT20), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n363), .B1(new_n640), .B2(new_n378), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n436), .A2(new_n638), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n642), .B(new_n317), .C1(new_n624), .C2(new_n625), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n436), .A2(new_n639), .A3(new_n641), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n644), .A2(KEYINPUT99), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n637), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n317), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n313), .B2(new_n315), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n644), .A2(KEYINPUT99), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(KEYINPUT100), .A3(new_n649), .A4(new_n642), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n623), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  OAI21_X1  g468(.A(new_n605), .B1(new_n620), .B2(new_n621), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n518), .B(KEYINPUT101), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n527), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n537), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n503), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  AOI22_X1  g479(.A1(G472), .A2(new_n591), .B1(new_n606), .B2(new_n612), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n666), .A2(new_n619), .A3(new_n661), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n387), .B1(new_n391), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n436), .A2(new_n641), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n667), .A2(new_n648), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NAND2_X1  g488(.A1(new_n580), .A2(new_n545), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n307), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n545), .B1(new_n561), .B2(new_n563), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n610), .A2(new_n611), .ZN(new_n679));
  AOI211_X1 g493(.A(KEYINPUT32), .B(new_n607), .C1(new_n608), .C2(new_n609), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n613), .A2(KEYINPUT102), .A3(new_n678), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT38), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT92), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n624), .A2(new_n625), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n687), .B1(new_n689), .B2(new_n318), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n316), .A2(KEYINPUT38), .A3(new_n319), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n686), .A2(new_n692), .A3(new_n660), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n669), .B(KEYINPUT39), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n619), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT103), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n695), .B(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n381), .A2(new_n317), .A3(new_n436), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n693), .A2(new_n697), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  INV_X1    g519(.A(new_n631), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n378), .A2(new_n377), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n640), .ZN(new_n708));
  INV_X1    g522(.A(new_n380), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n363), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n648), .A2(new_n711), .A3(new_n670), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n648), .A2(KEYINPUT104), .A3(new_n711), .A4(new_n670), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n667), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NAND2_X1  g532(.A1(new_n592), .A2(new_n613), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n497), .A2(new_n390), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n618), .A3(new_n500), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n719), .A2(new_n633), .A3(new_n538), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NOR3_X1   g540(.A1(new_n666), .A2(new_n539), .A3(new_n722), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n651), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  NOR2_X1   g543(.A1(new_n722), .A2(new_n626), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n719), .A2(new_n437), .A3(new_n730), .A4(new_n660), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  NOR2_X1   g546(.A1(new_n624), .A2(new_n625), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n702), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n599), .B1(new_n570), .B2(new_n545), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n593), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n538), .B(new_n736), .C1(new_n620), .C2(new_n621), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n734), .A2(new_n738), .A3(new_n639), .A4(new_n723), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  OAI21_X1  g554(.A(new_n736), .B1(new_n621), .B2(new_n620), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(new_n661), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n381), .A2(new_n631), .A3(new_n670), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n730), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  AOI21_X1  g561(.A(new_n647), .B1(new_n316), .B2(new_n319), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n501), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n614), .A3(new_n745), .A4(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n614), .A2(new_n501), .A3(new_n745), .A4(new_n748), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(KEYINPUT106), .B(G131), .Z(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G33));
  NAND3_X1  g572(.A1(new_n750), .A2(new_n614), .A3(new_n672), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  XOR2_X1   g574(.A(new_n489), .B(KEYINPUT45), .Z(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(G469), .ZN(new_n762));
  NAND2_X1  g576(.A1(G469), .A2(G902), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n765), .B(G469), .C1(new_n761), .C2(G902), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n500), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n618), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n694), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n710), .A2(new_n631), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n710), .A2(KEYINPUT43), .A3(new_n631), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n655), .A3(new_n660), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT44), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n748), .B(KEYINPUT107), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n769), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n768), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n767), .A2(KEYINPUT47), .A3(new_n618), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n744), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n666), .A3(new_n539), .A4(new_n748), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NOR2_X1   g599(.A1(G952), .A2(G953), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n689), .A2(new_n647), .A3(new_n318), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n434), .A2(new_n428), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n632), .B1(new_n788), .B2(new_n381), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n787), .A2(new_n623), .A3(new_n639), .A4(new_n789), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n724), .A2(new_n790), .A3(new_n731), .A4(new_n739), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n503), .B1(new_n614), .B2(new_n662), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n641), .A2(new_n788), .A3(new_n670), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT109), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n719), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n741), .A2(new_n744), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n750), .B(new_n660), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n791), .A2(new_n728), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n752), .A2(new_n755), .A3(new_n759), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n619), .A2(new_n669), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n685), .A2(new_n661), .A3(new_n734), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n717), .A2(new_n673), .A3(new_n803), .A4(new_n746), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n666), .A2(new_n619), .A3(new_n626), .A4(new_n661), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n672), .A2(new_n807), .B1(new_n716), .B2(new_n667), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(KEYINPUT52), .A3(new_n746), .A4(new_n803), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n801), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n798), .B2(new_n799), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n806), .A2(new_n809), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n728), .A2(new_n792), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n790), .A2(new_n724), .A3(new_n731), .A4(new_n739), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n796), .B1(new_n719), .B2(new_n794), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n816), .A2(new_n661), .A3(new_n749), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n799), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT110), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n812), .A2(new_n813), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AOI221_X4 g637(.A(KEYINPUT54), .B1(new_n800), .B2(new_n810), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n798), .A2(new_n811), .A3(new_n799), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT110), .B1(new_n818), .B2(new_n819), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n813), .A4(new_n822), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n821), .A2(new_n801), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n812), .A2(new_n820), .A3(new_n813), .A4(new_n822), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n824), .B1(new_n833), .B2(KEYINPUT54), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n683), .A2(new_n684), .A3(new_n723), .A4(new_n748), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n539), .A2(new_n386), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n835), .A2(new_n381), .A3(new_n631), .A4(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n748), .A2(new_n723), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n386), .B1(new_n772), .B2(new_n773), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n840), .A3(new_n743), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT113), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n647), .A3(new_n738), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n690), .A2(new_n691), .A3(new_n723), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT50), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n686), .A2(new_n706), .A3(new_n839), .A4(new_n836), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n848), .B(new_n841), .C1(new_n849), .C2(new_n381), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n843), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n721), .A2(new_n500), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n440), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n781), .A2(new_n782), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n840), .A2(new_n738), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n777), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n843), .A2(new_n847), .A3(KEYINPUT114), .A4(new_n850), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n853), .A2(KEYINPUT51), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n730), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT115), .Z(new_n863));
  INV_X1    g677(.A(KEYINPUT48), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n839), .A2(new_n840), .ZN(new_n865));
  INV_X1    g679(.A(new_n614), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT48), .A4(new_n614), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n686), .A2(new_n711), .A3(new_n839), .A4(new_n836), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n867), .A2(new_n383), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n838), .A2(new_n842), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n859), .A2(new_n871), .A3(new_n847), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n861), .A2(new_n863), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n786), .B1(new_n834), .B2(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n854), .A2(KEYINPUT108), .A3(KEYINPUT49), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n770), .B(new_n878), .C1(KEYINPUT108), .C2(KEYINPUT49), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n854), .B1(KEYINPUT108), .B2(KEYINPUT49), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n538), .A2(new_n880), .A3(new_n317), .A4(new_n618), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n692), .A3(new_n686), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT116), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n875), .B(new_n824), .C1(KEYINPUT54), .C2(new_n833), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n885), .B(new_n882), .C1(new_n886), .C2(new_n786), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(G75));
  NAND2_X1  g702(.A1(new_n286), .A2(new_n276), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n218), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT55), .Z(new_n891));
  NAND2_X1  g705(.A1(new_n821), .A2(new_n823), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n810), .A2(new_n800), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n390), .B(new_n311), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT117), .B1(new_n894), .B2(KEYINPUT56), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n893), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n389), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n896), .B(new_n897), .C1(new_n899), .C2(new_n311), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n891), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n891), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n382), .A2(G953), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT118), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(G51));
  XNOR2_X1  g720(.A(new_n898), .B(KEYINPUT54), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n763), .B(KEYINPUT57), .Z(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n497), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n899), .A2(new_n762), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(G54));
  INV_X1    g726(.A(KEYINPUT58), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n899), .A2(new_n913), .A3(new_n321), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n360), .A2(new_n374), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n905), .B1(new_n916), .B2(new_n917), .ZN(G60));
  XNOR2_X1  g732(.A(new_n628), .B(KEYINPUT119), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n834), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n919), .ZN(new_n923));
  INV_X1    g737(.A(new_n921), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n907), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n922), .A2(new_n925), .A3(new_n904), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT120), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT60), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n898), .A2(new_n658), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n525), .B1(new_n898), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n905), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g747(.A(G953), .B1(new_n393), .B2(new_n214), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n814), .A2(new_n815), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(G953), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n889), .B1(G898), .B2(new_n388), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G69));
  NAND3_X1  g752(.A1(new_n717), .A2(new_n673), .A3(new_n746), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n808), .A2(KEYINPUT122), .A3(new_n746), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n769), .A2(new_n614), .A3(new_n734), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n784), .A2(new_n941), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n799), .B(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n946), .A2(new_n778), .ZN(new_n947));
  AOI21_X1  g761(.A(G953), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n577), .A2(new_n578), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT121), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n367), .B1(new_n370), .B2(new_n365), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(G227), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n953), .B2(new_n668), .ZN(new_n954));
  AND2_X1   g768(.A1(KEYINPUT124), .A2(G900), .ZN(new_n955));
  NOR2_X1   g769(.A1(KEYINPUT124), .A2(G900), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n948), .A2(new_n952), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n704), .A2(new_n941), .A3(new_n942), .A4(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n960), .A2(new_n778), .ZN(new_n961));
  AND4_X1   g775(.A1(new_n614), .A2(new_n695), .A3(new_n748), .A4(new_n789), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n941), .A2(new_n704), .A3(new_n942), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(KEYINPUT62), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n961), .A2(new_n784), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n954), .B1(new_n965), .B2(G953), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n958), .B1(new_n966), .B2(new_n952), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT125), .ZN(G72));
  NAND4_X1  g782(.A1(new_n961), .A2(new_n784), .A3(new_n964), .A4(new_n935), .ZN(new_n969));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  AOI21_X1  g785(.A(new_n675), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n904), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n580), .A2(new_n545), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n944), .A2(new_n935), .A3(new_n947), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n971), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n675), .A3(new_n971), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT127), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n833), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n975), .A2(new_n979), .A3(new_n982), .ZN(G57));
endmodule


