

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U324 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U325 ( .A(KEYINPUT99), .B(KEYINPUT37), .ZN(n472) );
  XOR2_X1 U326 ( .A(n463), .B(KEYINPUT28), .Z(n531) );
  XNOR2_X1 U327 ( .A(n345), .B(n445), .ZN(n517) );
  INV_X1 U328 ( .A(G197GAT), .ZN(n330) );
  XNOR2_X1 U329 ( .A(n331), .B(n330), .ZN(n333) );
  XNOR2_X1 U330 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n415) );
  XNOR2_X1 U331 ( .A(n333), .B(n332), .ZN(n431) );
  XNOR2_X1 U332 ( .A(n336), .B(n373), .ZN(n337) );
  XNOR2_X1 U333 ( .A(KEYINPUT98), .B(KEYINPUT36), .ZN(n387) );
  XNOR2_X1 U334 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U335 ( .A(n338), .B(n337), .ZN(n340) );
  XNOR2_X1 U336 ( .A(n564), .B(n387), .ZN(n585) );
  XNOR2_X1 U337 ( .A(n435), .B(n434), .ZN(n450) );
  XNOR2_X1 U338 ( .A(n381), .B(n380), .ZN(n386) );
  XNOR2_X1 U339 ( .A(n473), .B(n472), .ZN(n514) );
  INV_X1 U340 ( .A(G169GAT), .ZN(n451) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n475) );
  XOR2_X1 U342 ( .A(n449), .B(n448), .Z(n533) );
  XNOR2_X1 U343 ( .A(n451), .B(KEYINPUT120), .ZN(n452) );
  XNOR2_X1 U344 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U345 ( .A(n453), .B(n452), .ZN(G1348GAT) );
  XNOR2_X1 U346 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT69), .B(G15GAT), .Z(n293) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(G113GAT), .ZN(n292) );
  XNOR2_X1 U349 ( .A(n293), .B(n292), .ZN(n310) );
  XOR2_X1 U350 ( .A(G197GAT), .B(G141GAT), .Z(n295) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(G22GAT), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n297) );
  XOR2_X1 U353 ( .A(G50GAT), .B(G36GAT), .Z(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n306) );
  XNOR2_X1 U355 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n298), .B(KEYINPUT29), .ZN(n299) );
  XOR2_X1 U357 ( .A(n299), .B(KEYINPUT66), .Z(n304) );
  XOR2_X1 U358 ( .A(G29GAT), .B(KEYINPUT67), .Z(n301) );
  XNOR2_X1 U359 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n375) );
  XNOR2_X1 U361 ( .A(G1GAT), .B(G8GAT), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n302), .B(KEYINPUT68), .ZN(n351) );
  XNOR2_X1 U363 ( .A(n375), .B(n351), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n306), .B(n305), .ZN(n308) );
  NAND2_X1 U366 ( .A1(G229GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n570) );
  XOR2_X1 U369 ( .A(KEYINPUT1), .B(KEYINPUT89), .Z(n312) );
  XNOR2_X1 U370 ( .A(G1GAT), .B(KEYINPUT90), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n329) );
  XOR2_X1 U372 ( .A(KEYINPUT77), .B(G162GAT), .Z(n314) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(G134GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U375 ( .A(G155GAT), .B(G148GAT), .Z(n316) );
  XNOR2_X1 U376 ( .A(G127GAT), .B(G120GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U378 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U379 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n320) );
  NAND2_X1 U380 ( .A1(G225GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U382 ( .A(KEYINPUT5), .B(n321), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U384 ( .A(G85GAT), .B(G57GAT), .Z(n390) );
  XOR2_X1 U385 ( .A(n324), .B(n390), .Z(n327) );
  XOR2_X1 U386 ( .A(G113GAT), .B(KEYINPUT0), .Z(n444) );
  XNOR2_X1 U387 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n325), .B(KEYINPUT2), .ZN(n428) );
  XNOR2_X1 U389 ( .A(n444), .B(n428), .ZN(n326) );
  XNOR2_X1 U390 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n515) );
  XNOR2_X1 U392 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n331) );
  XOR2_X1 U393 ( .A(KEYINPUT87), .B(G218GAT), .Z(n332) );
  XNOR2_X1 U394 ( .A(G8GAT), .B(n431), .ZN(n338) );
  XOR2_X1 U395 ( .A(G64GAT), .B(G92GAT), .Z(n335) );
  XNOR2_X1 U396 ( .A(G176GAT), .B(G204GAT), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n400) );
  XOR2_X1 U398 ( .A(KEYINPUT91), .B(n400), .Z(n336) );
  XOR2_X1 U399 ( .A(G36GAT), .B(G190GAT), .Z(n373) );
  AND2_X1 U400 ( .A1(G226GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n345) );
  XNOR2_X1 U402 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n341), .B(KEYINPUT83), .ZN(n342) );
  XOR2_X1 U404 ( .A(n342), .B(KEYINPUT18), .Z(n344) );
  XNOR2_X1 U405 ( .A(G169GAT), .B(G183GAT), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n445) );
  XOR2_X1 U407 ( .A(KEYINPUT117), .B(n517), .Z(n414) );
  XOR2_X1 U408 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n389) );
  XOR2_X1 U409 ( .A(G64GAT), .B(G57GAT), .Z(n347) );
  XNOR2_X1 U410 ( .A(G211GAT), .B(G78GAT), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U412 ( .A(n348), .B(G71GAT), .Z(n350) );
  XOR2_X1 U413 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XNOR2_X1 U414 ( .A(G183GAT), .B(n442), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n355) );
  XOR2_X1 U416 ( .A(G22GAT), .B(G155GAT), .Z(n420) );
  XOR2_X1 U417 ( .A(n420), .B(n351), .Z(n353) );
  NAND2_X1 U418 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U420 ( .A(n355), .B(n354), .Z(n363) );
  XOR2_X1 U421 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n357) );
  XNOR2_X1 U422 ( .A(KEYINPUT13), .B(KEYINPUT80), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n359) );
  XNOR2_X1 U425 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n582) );
  INV_X1 U429 ( .A(KEYINPUT77), .ZN(n364) );
  NAND2_X1 U430 ( .A1(G92GAT), .A2(n364), .ZN(n367) );
  INV_X1 U431 ( .A(G92GAT), .ZN(n365) );
  NAND2_X1 U432 ( .A1(n365), .A2(KEYINPUT77), .ZN(n366) );
  NAND2_X1 U433 ( .A1(n367), .A2(n366), .ZN(n369) );
  XNOR2_X1 U434 ( .A(G106GAT), .B(G85GAT), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n370), .B(G218GAT), .ZN(n372) );
  XOR2_X1 U437 ( .A(G43GAT), .B(G134GAT), .Z(n439) );
  XOR2_X1 U438 ( .A(n439), .B(G99GAT), .Z(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n374) );
  XOR2_X1 U440 ( .A(n374), .B(n373), .Z(n381) );
  XOR2_X1 U441 ( .A(G50GAT), .B(G162GAT), .Z(n421) );
  XNOR2_X1 U442 ( .A(n375), .B(n421), .ZN(n379) );
  XOR2_X1 U443 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n377) );
  NAND2_X1 U444 ( .A1(G232GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U445 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U446 ( .A(KEYINPUT75), .B(KEYINPUT64), .Z(n383) );
  XNOR2_X1 U447 ( .A(KEYINPUT9), .B(KEYINPUT74), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U449 ( .A(n384), .B(KEYINPUT76), .Z(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n564) );
  NOR2_X1 U451 ( .A1(n582), .A2(n585), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n405) );
  XNOR2_X1 U453 ( .A(n390), .B(KEYINPUT70), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n391), .B(KEYINPUT72), .ZN(n404) );
  XNOR2_X1 U455 ( .A(G106GAT), .B(G78GAT), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n392), .B(G148GAT), .ZN(n430) );
  XOR2_X1 U457 ( .A(n430), .B(KEYINPUT71), .Z(n394) );
  NAND2_X1 U458 ( .A1(G230GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U460 ( .A(KEYINPUT32), .B(KEYINPUT13), .Z(n396) );
  XNOR2_X1 U461 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U463 ( .A(n398), .B(n397), .Z(n402) );
  XNOR2_X1 U464 ( .A(G99GAT), .B(G71GAT), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n399), .B(G120GAT), .ZN(n438) );
  XNOR2_X1 U466 ( .A(n438), .B(n400), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n576) );
  NOR2_X1 U469 ( .A1(n405), .A2(n576), .ZN(n406) );
  NAND2_X1 U470 ( .A1(n406), .A2(n570), .ZN(n412) );
  NAND2_X1 U471 ( .A1(n564), .A2(n582), .ZN(n409) );
  XNOR2_X1 U472 ( .A(KEYINPUT41), .B(n576), .ZN(n547) );
  NOR2_X1 U473 ( .A1(n547), .A2(n570), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n407), .B(KEYINPUT46), .ZN(n408) );
  NOR2_X1 U475 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n410), .B(KEYINPUT47), .ZN(n411) );
  NAND2_X1 U477 ( .A1(n412), .A2(n411), .ZN(n413) );
  XNOR2_X1 U478 ( .A(KEYINPUT48), .B(n413), .ZN(n526) );
  NAND2_X1 U479 ( .A1(n414), .A2(n526), .ZN(n416) );
  NOR2_X1 U480 ( .A1(n515), .A2(n417), .ZN(n569) );
  XOR2_X1 U481 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n419) );
  XNOR2_X1 U482 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n425) );
  XOR2_X1 U484 ( .A(G204GAT), .B(KEYINPUT23), .Z(n423) );
  XNOR2_X1 U485 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U487 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U490 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n463) );
  NAND2_X1 U493 ( .A1(n569), .A2(n463), .ZN(n435) );
  XOR2_X1 U494 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n434) );
  XOR2_X1 U495 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n437) );
  XNOR2_X1 U496 ( .A(G190GAT), .B(G176GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n449) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U501 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n448) );
  NAND2_X1 U504 ( .A1(n450), .A2(n533), .ZN(n563) );
  NOR2_X1 U505 ( .A1(n570), .A2(n563), .ZN(n453) );
  NOR2_X1 U506 ( .A1(n576), .A2(n570), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(KEYINPUT73), .ZN(n485) );
  NAND2_X1 U508 ( .A1(n517), .A2(n533), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n455), .A2(n463), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n456), .B(KEYINPUT25), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT95), .B(n457), .Z(n461) );
  NOR2_X1 U512 ( .A1(n533), .A2(n463), .ZN(n458) );
  XOR2_X1 U513 ( .A(KEYINPUT26), .B(n458), .Z(n459) );
  XOR2_X1 U514 ( .A(KEYINPUT94), .B(n459), .Z(n568) );
  XNOR2_X1 U515 ( .A(n517), .B(KEYINPUT27), .ZN(n464) );
  AND2_X1 U516 ( .A1(n568), .A2(n464), .ZN(n460) );
  NOR2_X1 U517 ( .A1(n461), .A2(n460), .ZN(n462) );
  NOR2_X1 U518 ( .A1(n515), .A2(n462), .ZN(n470) );
  NAND2_X1 U519 ( .A1(n464), .A2(n515), .ZN(n527) );
  NOR2_X1 U520 ( .A1(n531), .A2(n527), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT92), .B(n465), .Z(n467) );
  XOR2_X1 U522 ( .A(n533), .B(KEYINPUT85), .Z(n466) );
  OR2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U524 ( .A(KEYINPUT93), .B(n468), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n470), .A2(n469), .ZN(n483) );
  NOR2_X1 U526 ( .A1(n585), .A2(n483), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n582), .A2(n471), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n485), .A2(n514), .ZN(n474) );
  XNOR2_X1 U529 ( .A(n474), .B(KEYINPUT38), .ZN(n499) );
  NAND2_X1 U530 ( .A1(n533), .A2(n499), .ZN(n478) );
  XOR2_X1 U531 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n476) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n487) );
  INV_X1 U533 ( .A(n582), .ZN(n479) );
  NAND2_X1 U534 ( .A1(n479), .A2(n564), .ZN(n480) );
  XNOR2_X1 U535 ( .A(n480), .B(KEYINPUT16), .ZN(n481) );
  XNOR2_X1 U536 ( .A(n481), .B(KEYINPUT82), .ZN(n482) );
  NOR2_X1 U537 ( .A1(n483), .A2(n482), .ZN(n484) );
  XOR2_X1 U538 ( .A(KEYINPUT96), .B(n484), .Z(n502) );
  NOR2_X1 U539 ( .A1(n502), .A2(n485), .ZN(n492) );
  NAND2_X1 U540 ( .A1(n492), .A2(n515), .ZN(n486) );
  XNOR2_X1 U541 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U542 ( .A1(n517), .A2(n492), .ZN(n488) );
  XNOR2_X1 U543 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U545 ( .A1(n492), .A2(n533), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U547 ( .A(G15GAT), .B(n491), .Z(G1326GAT) );
  NAND2_X1 U548 ( .A1(n492), .A2(n531), .ZN(n493) );
  XNOR2_X1 U549 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U550 ( .A1(n515), .A2(n499), .ZN(n495) );
  XOR2_X1 U551 ( .A(KEYINPUT39), .B(KEYINPUT100), .Z(n494) );
  XNOR2_X1 U552 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(n496), .ZN(G1328GAT) );
  XOR2_X1 U554 ( .A(G36GAT), .B(KEYINPUT101), .Z(n498) );
  NAND2_X1 U555 ( .A1(n499), .A2(n517), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n499), .A2(n531), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n504) );
  XNOR2_X1 U560 ( .A(n547), .B(KEYINPUT104), .ZN(n556) );
  INV_X1 U561 ( .A(n556), .ZN(n501) );
  NAND2_X1 U562 ( .A1(n501), .A2(n570), .ZN(n513) );
  NOR2_X1 U563 ( .A1(n502), .A2(n513), .ZN(n509) );
  NAND2_X1 U564 ( .A1(n509), .A2(n515), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  XOR2_X1 U567 ( .A(G64GAT), .B(KEYINPUT105), .Z(n507) );
  NAND2_X1 U568 ( .A1(n509), .A2(n517), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1333GAT) );
  NAND2_X1 U570 ( .A1(n509), .A2(n533), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U573 ( .A1(n509), .A2(n531), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U576 ( .A1(n514), .A2(n513), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n522), .A2(n515), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n517), .A2(n522), .ZN(n518) );
  XNOR2_X1 U580 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n520) );
  NAND2_X1 U582 ( .A1(n522), .A2(n533), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n524) );
  NAND2_X1 U586 ( .A1(n522), .A2(n531), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  INV_X1 U589 ( .A(n526), .ZN(n528) );
  NOR2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U591 ( .A(KEYINPUT111), .B(n529), .Z(n545) );
  INV_X1 U592 ( .A(n545), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n540) );
  NOR2_X1 U595 ( .A1(n570), .A2(n540), .ZN(n534) );
  XOR2_X1 U596 ( .A(n534), .B(KEYINPUT112), .Z(n535) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  NOR2_X1 U598 ( .A1(n556), .A2(n540), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NOR2_X1 U601 ( .A1(n582), .A2(n540), .ZN(n538) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(n538), .Z(n539) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  NOR2_X1 U604 ( .A1(n540), .A2(n564), .ZN(n544) );
  XOR2_X1 U605 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n542) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n568), .A2(n545), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n570), .A2(n553), .ZN(n546) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n547), .A2(n553), .ZN(n549) );
  XNOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n582), .A2(n553), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT115), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n564), .A2(n553), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT116), .B(n554), .Z(n555) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  NOR2_X1 U622 ( .A1(n563), .A2(n556), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n558) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(KEYINPUT56), .B(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n582), .A2(n563), .ZN(n562) );
  XOR2_X1 U629 ( .A(G183GAT), .B(n562), .Z(G1350GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n584) );
  NOR2_X1 U635 ( .A1(n570), .A2(n584), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(KEYINPUT124), .B(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  INV_X1 U641 ( .A(n576), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n584), .A2(n577), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n579) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n584), .ZN(n583) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

