

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  NOR2_X1 U322 ( .A1(n429), .A2(n428), .ZN(n430) );
  OR2_X1 U323 ( .A1(n450), .A2(n503), .ZN(n451) );
  XOR2_X1 U324 ( .A(n393), .B(n425), .Z(n547) );
  XOR2_X1 U325 ( .A(n392), .B(n391), .Z(n425) );
  XNOR2_X1 U326 ( .A(n430), .B(KEYINPUT48), .ZN(n539) );
  XNOR2_X1 U327 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n394) );
  XNOR2_X1 U328 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U329 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U330 ( .A(n385), .B(n384), .ZN(n390) );
  XNOR2_X1 U331 ( .A(n366), .B(n365), .ZN(n367) );
  INV_X1 U332 ( .A(n539), .ZN(n540) );
  XNOR2_X1 U333 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U334 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U335 ( .A(n451), .B(KEYINPUT123), .ZN(n562) );
  XOR2_X1 U336 ( .A(n449), .B(n448), .Z(n523) );
  XNOR2_X1 U337 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n452) );
  XOR2_X1 U338 ( .A(G106GAT), .B(KEYINPUT77), .Z(n291) );
  NAND2_X1 U339 ( .A1(G232GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U340 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U341 ( .A(G134GAT), .B(n292), .ZN(n304) );
  XOR2_X1 U342 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n294) );
  XNOR2_X1 U343 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U345 ( .A(G36GAT), .B(G190GAT), .Z(n347) );
  XOR2_X1 U346 ( .A(n295), .B(n347), .Z(n299) );
  XOR2_X1 U347 ( .A(G29GAT), .B(G43GAT), .Z(n297) );
  XNOR2_X1 U348 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n368) );
  XOR2_X1 U350 ( .A(G50GAT), .B(G162GAT), .Z(n326) );
  XNOR2_X1 U351 ( .A(n368), .B(n326), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U353 ( .A(n300), .B(KEYINPUT78), .Z(n302) );
  XOR2_X1 U354 ( .A(G99GAT), .B(G85GAT), .Z(n378) );
  XNOR2_X1 U355 ( .A(G218GAT), .B(n378), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U357 ( .A(n304), .B(n303), .Z(n551) );
  XOR2_X1 U358 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n306) );
  XNOR2_X1 U359 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n324) );
  XOR2_X1 U361 ( .A(G85GAT), .B(G162GAT), .Z(n308) );
  XNOR2_X1 U362 ( .A(G29GAT), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U364 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n310) );
  XNOR2_X1 U365 ( .A(G1GAT), .B(G148GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U367 ( .A(n312), .B(n311), .Z(n322) );
  XOR2_X1 U368 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n314) );
  XNOR2_X1 U369 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U371 ( .A(G141GAT), .B(n315), .Z(n339) );
  XOR2_X1 U372 ( .A(G120GAT), .B(KEYINPUT0), .Z(n317) );
  XNOR2_X1 U373 ( .A(G113GAT), .B(G134GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n441) );
  XOR2_X1 U375 ( .A(G57GAT), .B(n441), .Z(n319) );
  NAND2_X1 U376 ( .A1(G225GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n339), .B(n320), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n495) );
  XOR2_X1 U381 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n328) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(G78GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n325), .B(G148GAT), .ZN(n388) );
  XNOR2_X1 U384 ( .A(n326), .B(n388), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U386 ( .A(KEYINPUT23), .B(G204GAT), .Z(n330) );
  NAND2_X1 U387 ( .A1(G228GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U389 ( .A(n332), .B(n331), .Z(n337) );
  XOR2_X1 U390 ( .A(KEYINPUT21), .B(G218GAT), .Z(n334) );
  XNOR2_X1 U391 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U393 ( .A(G197GAT), .B(n335), .Z(n355) );
  XNOR2_X1 U394 ( .A(G22GAT), .B(n355), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n463) );
  NAND2_X1 U397 ( .A1(n495), .A2(n463), .ZN(n432) );
  XOR2_X1 U398 ( .A(KEYINPUT97), .B(KEYINPUT94), .Z(n341) );
  XNOR2_X1 U399 ( .A(KEYINPUT79), .B(KEYINPUT95), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U401 ( .A(n342), .B(KEYINPUT93), .Z(n344) );
  XOR2_X1 U402 ( .A(G169GAT), .B(G8GAT), .Z(n358) );
  XNOR2_X1 U403 ( .A(n358), .B(KEYINPUT96), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n351) );
  XOR2_X1 U405 ( .A(G183GAT), .B(KEYINPUT18), .Z(n346) );
  XNOR2_X1 U406 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n439) );
  XOR2_X1 U408 ( .A(n347), .B(n439), .Z(n349) );
  NAND2_X1 U409 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U411 ( .A(n351), .B(n350), .Z(n357) );
  XOR2_X1 U412 ( .A(G92GAT), .B(G64GAT), .Z(n353) );
  XNOR2_X1 U413 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U415 ( .A(G204GAT), .B(n354), .Z(n392) );
  XNOR2_X1 U416 ( .A(n355), .B(n392), .ZN(n356) );
  XOR2_X1 U417 ( .A(n357), .B(n356), .Z(n513) );
  INV_X1 U418 ( .A(n513), .ZN(n501) );
  XOR2_X1 U419 ( .A(G36GAT), .B(G50GAT), .Z(n360) );
  XOR2_X1 U420 ( .A(G22GAT), .B(G1GAT), .Z(n403) );
  XNOR2_X1 U421 ( .A(n358), .B(n403), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n366) );
  XOR2_X1 U423 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n362) );
  XNOR2_X1 U424 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n364) );
  AND2_X1 U426 ( .A1(G229GAT), .A2(G233GAT), .ZN(n363) );
  XOR2_X1 U427 ( .A(n367), .B(KEYINPUT30), .Z(n374) );
  XNOR2_X1 U428 ( .A(n368), .B(KEYINPUT69), .ZN(n372) );
  XOR2_X1 U429 ( .A(G197GAT), .B(G141GAT), .Z(n370) );
  XNOR2_X1 U430 ( .A(G15GAT), .B(G113GAT), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n370), .B(n369), .ZN(n371) );
  INV_X1 U432 ( .A(n375), .ZN(n568) );
  XNOR2_X1 U433 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n393) );
  XOR2_X1 U434 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n377) );
  XNOR2_X1 U435 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n385) );
  XOR2_X1 U438 ( .A(KEYINPUT76), .B(KEYINPUT73), .Z(n381) );
  XNOR2_X1 U439 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n383) );
  AND2_X1 U441 ( .A1(G230GAT), .A2(G233GAT), .ZN(n382) );
  XOR2_X1 U442 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n387) );
  XNOR2_X1 U443 ( .A(G71GAT), .B(G57GAT), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n398) );
  XOR2_X1 U445 ( .A(n388), .B(n398), .Z(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n391) );
  NAND2_X1 U447 ( .A1(n568), .A2(n547), .ZN(n395) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n418) );
  XOR2_X1 U449 ( .A(G78GAT), .B(G211GAT), .Z(n397) );
  XNOR2_X1 U450 ( .A(G183GAT), .B(G155GAT), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n402) );
  XOR2_X1 U452 ( .A(n398), .B(KEYINPUT12), .Z(n400) );
  NAND2_X1 U453 ( .A1(G231GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U455 ( .A(n402), .B(n401), .Z(n405) );
  XOR2_X1 U456 ( .A(G15GAT), .B(G127GAT), .Z(n444) );
  XNOR2_X1 U457 ( .A(n403), .B(n444), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U459 ( .A(KEYINPUT85), .B(KEYINPUT79), .Z(n407) );
  XNOR2_X1 U460 ( .A(G8GAT), .B(G64GAT), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U462 ( .A(n409), .B(n408), .Z(n417) );
  XOR2_X1 U463 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n411) );
  XNOR2_X1 U464 ( .A(KEYINPUT83), .B(KEYINPUT14), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U466 ( .A(KEYINPUT82), .B(KEYINPUT86), .Z(n413) );
  XNOR2_X1 U467 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n575) );
  NOR2_X1 U471 ( .A1(n418), .A2(n575), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n419), .B(KEYINPUT112), .ZN(n420) );
  INV_X1 U473 ( .A(n551), .ZN(n455) );
  NAND2_X1 U474 ( .A1(n420), .A2(n455), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n421), .B(KEYINPUT47), .ZN(n429) );
  XOR2_X1 U476 ( .A(KEYINPUT36), .B(n455), .Z(n577) );
  NAND2_X1 U477 ( .A1(n577), .A2(n575), .ZN(n424) );
  XOR2_X1 U478 ( .A(KEYINPUT113), .B(KEYINPUT45), .Z(n422) );
  XNOR2_X1 U479 ( .A(KEYINPUT65), .B(n422), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n426) );
  INV_X1 U481 ( .A(n425), .ZN(n454) );
  NAND2_X1 U482 ( .A1(n426), .A2(n454), .ZN(n427) );
  NOR2_X1 U483 ( .A1(n427), .A2(n568), .ZN(n428) );
  NOR2_X1 U484 ( .A1(n501), .A2(n539), .ZN(n431) );
  XOR2_X1 U485 ( .A(KEYINPUT54), .B(n431), .Z(n564) );
  OR2_X1 U486 ( .A1(n432), .A2(n564), .ZN(n434) );
  XOR2_X1 U487 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n450) );
  XOR2_X1 U489 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n436) );
  XNOR2_X1 U490 ( .A(G99GAT), .B(G176GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n449) );
  XOR2_X1 U492 ( .A(KEYINPUT20), .B(G71GAT), .Z(n438) );
  NAND2_X1 U493 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n443) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U498 ( .A(n445), .B(n444), .Z(n447) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(G190GAT), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  INV_X1 U501 ( .A(n523), .ZN(n503) );
  NAND2_X1 U502 ( .A1(n551), .A2(n562), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XNOR2_X1 U504 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n472) );
  INV_X1 U505 ( .A(n495), .ZN(n565) );
  NAND2_X1 U506 ( .A1(n568), .A2(n454), .ZN(n482) );
  NAND2_X1 U507 ( .A1(n455), .A2(n575), .ZN(n456) );
  XOR2_X1 U508 ( .A(KEYINPUT16), .B(n456), .Z(n470) );
  XOR2_X1 U509 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n457) );
  XOR2_X1 U510 ( .A(n463), .B(n457), .Z(n506) );
  INV_X1 U511 ( .A(n506), .ZN(n517) );
  XNOR2_X1 U512 ( .A(n513), .B(KEYINPUT27), .ZN(n461) );
  NAND2_X1 U513 ( .A1(n565), .A2(n461), .ZN(n537) );
  NOR2_X1 U514 ( .A1(n517), .A2(n537), .ZN(n522) );
  NAND2_X1 U515 ( .A1(n522), .A2(n503), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n458), .B(KEYINPUT98), .ZN(n469) );
  NOR2_X1 U517 ( .A1(n523), .A2(n463), .ZN(n460) );
  XNOR2_X1 U518 ( .A(KEYINPUT99), .B(KEYINPUT26), .ZN(n459) );
  XOR2_X1 U519 ( .A(n460), .B(n459), .Z(n567) );
  NAND2_X1 U520 ( .A1(n567), .A2(n461), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n523), .A2(n513), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n467), .A2(n495), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n479) );
  NAND2_X1 U527 ( .A1(n470), .A2(n479), .ZN(n493) );
  NOR2_X1 U528 ( .A1(n482), .A2(n493), .ZN(n476) );
  NAND2_X1 U529 ( .A1(n565), .A2(n476), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U531 ( .A1(n513), .A2(n476), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U534 ( .A1(n476), .A2(n523), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  NAND2_X1 U536 ( .A1(n476), .A2(n517), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(KEYINPUT100), .ZN(n478) );
  XNOR2_X1 U538 ( .A(G22GAT), .B(n478), .ZN(G1327GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n486) );
  NAND2_X1 U540 ( .A1(n577), .A2(n479), .ZN(n480) );
  NOR2_X1 U541 ( .A1(n480), .A2(n575), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(KEYINPUT37), .ZN(n510) );
  NOR2_X1 U543 ( .A1(n510), .A2(n482), .ZN(n483) );
  XOR2_X1 U544 ( .A(KEYINPUT101), .B(n483), .Z(n484) );
  XNOR2_X1 U545 ( .A(KEYINPUT38), .B(n484), .ZN(n491) );
  NAND2_X1 U546 ( .A1(n565), .A2(n491), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(n487), .ZN(G1328GAT) );
  NAND2_X1 U549 ( .A1(n491), .A2(n513), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U551 ( .A1(n491), .A2(n523), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(KEYINPUT40), .ZN(n490) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  NAND2_X1 U554 ( .A1(n491), .A2(n517), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n492), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U556 ( .A(KEYINPUT104), .B(n547), .ZN(n559) );
  NAND2_X1 U557 ( .A1(n559), .A2(n375), .ZN(n509) );
  NOR2_X1 U558 ( .A1(n493), .A2(n509), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n494), .B(KEYINPUT105), .ZN(n505) );
  NOR2_X1 U560 ( .A1(n495), .A2(n505), .ZN(n500) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n497) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U564 ( .A(KEYINPUT103), .B(n498), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n501), .A2(n505), .ZN(n502) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n502), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n503), .A2(n505), .ZN(n504) );
  XOR2_X1 U569 ( .A(G71GAT), .B(n504), .Z(G1334GAT) );
  NOR2_X1 U570 ( .A1(n506), .A2(n505), .ZN(n508) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  XNOR2_X1 U573 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n512) );
  NOR2_X1 U574 ( .A1(n510), .A2(n509), .ZN(n518) );
  NAND2_X1 U575 ( .A1(n565), .A2(n518), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n518), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U579 ( .A(G99GAT), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U580 ( .A1(n518), .A2(n523), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1338GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n520) );
  NAND2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U585 ( .A(G106GAT), .B(n521), .Z(G1339GAT) );
  NAND2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U587 ( .A1(n524), .A2(n539), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n525), .B(KEYINPUT114), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n568), .A2(n532), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U592 ( .A1(n559), .A2(n532), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n530) );
  NAND2_X1 U595 ( .A1(n575), .A2(n532), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U599 ( .A1(n532), .A2(n551), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT116), .Z(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  INV_X1 U603 ( .A(n567), .ZN(n538) );
  NOR2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n541) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT118), .B(n542), .Z(n552) );
  NAND2_X1 U607 ( .A1(n552), .A2(n568), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n543), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT119), .B(n546), .Z(n549) );
  NAND2_X1 U613 ( .A1(n552), .A2(n547), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n552), .A2(n575), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U617 ( .A(G162GAT), .B(KEYINPUT121), .Z(n554) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n562), .A2(n568), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(n558), .Z(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n562), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n575), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n578) );
  NAND2_X1 U633 ( .A1(n578), .A2(n568), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n578), .A2(n425), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n578), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

