

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594;

  NOR2_X1 U326 ( .A1(n470), .A2(n469), .ZN(n485) );
  XNOR2_X1 U327 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U328 ( .A(n365), .B(n364), .Z(n294) );
  XNOR2_X1 U329 ( .A(n415), .B(KEYINPUT109), .ZN(n416) );
  XNOR2_X1 U330 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U331 ( .A(KEYINPUT21), .B(G197GAT), .Z(n356) );
  XNOR2_X1 U332 ( .A(n371), .B(n370), .ZN(n372) );
  INV_X1 U333 ( .A(KEYINPUT37), .ZN(n473) );
  XNOR2_X1 U334 ( .A(n373), .B(n372), .ZN(n375) );
  XNOR2_X1 U335 ( .A(n473), .B(KEYINPUT100), .ZN(n474) );
  XNOR2_X1 U336 ( .A(n339), .B(n338), .ZN(n343) );
  XNOR2_X1 U337 ( .A(n475), .B(n474), .ZN(n519) );
  XOR2_X1 U338 ( .A(n466), .B(KEYINPUT28), .Z(n527) );
  XNOR2_X1 U339 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U340 ( .A(n478), .B(KEYINPUT39), .ZN(n479) );
  XNOR2_X1 U341 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n480), .B(n479), .ZN(G1328GAT) );
  XNOR2_X1 U343 ( .A(G85GAT), .B(KEYINPUT72), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n295), .B(G99GAT), .ZN(n367) );
  XOR2_X1 U345 ( .A(G162GAT), .B(G50GAT), .Z(n333) );
  XOR2_X1 U346 ( .A(n367), .B(n333), .Z(n297) );
  NAND2_X1 U347 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n311) );
  XOR2_X1 U349 ( .A(KEYINPUT75), .B(KEYINPUT9), .Z(n299) );
  XNOR2_X1 U350 ( .A(KEYINPUT10), .B(KEYINPUT64), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U352 ( .A(G92GAT), .B(G106GAT), .Z(n301) );
  XNOR2_X1 U353 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U355 ( .A(n303), .B(n302), .Z(n309) );
  XOR2_X1 U356 ( .A(G36GAT), .B(G190GAT), .Z(n305) );
  XNOR2_X1 U357 ( .A(G218GAT), .B(KEYINPUT76), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n350) );
  XOR2_X1 U359 ( .A(G43GAT), .B(KEYINPUT7), .Z(n307) );
  XNOR2_X1 U360 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n382) );
  XNOR2_X1 U362 ( .A(n350), .B(n382), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n544) );
  INV_X1 U365 ( .A(n544), .ZN(n561) );
  NAND2_X1 U366 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XOR2_X1 U367 ( .A(G127GAT), .B(G15GAT), .Z(n401) );
  XNOR2_X1 U368 ( .A(n312), .B(n401), .ZN(n326) );
  XOR2_X1 U369 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n314) );
  XNOR2_X1 U370 ( .A(G71GAT), .B(G176GAT), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U372 ( .A(G183GAT), .B(G99GAT), .Z(n316) );
  XNOR2_X1 U373 ( .A(G190GAT), .B(G43GAT), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U375 ( .A(n318), .B(n317), .Z(n324) );
  XOR2_X1 U376 ( .A(G113GAT), .B(G120GAT), .Z(n320) );
  XNOR2_X1 U377 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n444) );
  XOR2_X1 U379 ( .A(G169GAT), .B(KEYINPUT19), .Z(n322) );
  XNOR2_X1 U380 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n345) );
  XNOR2_X1 U382 ( .A(n444), .B(n345), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U384 ( .A(n326), .B(n325), .Z(n494) );
  XOR2_X1 U385 ( .A(KEYINPUT23), .B(n356), .Z(n328) );
  XOR2_X1 U386 ( .A(G155GAT), .B(G22GAT), .Z(n397) );
  XNOR2_X1 U387 ( .A(G218GAT), .B(n397), .ZN(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U389 ( .A(KEYINPUT85), .B(G204GAT), .Z(n330) );
  NAND2_X1 U390 ( .A1(G228GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n339) );
  XOR2_X1 U393 ( .A(n333), .B(G211GAT), .Z(n337) );
  XOR2_X1 U394 ( .A(KEYINPUT84), .B(KEYINPUT24), .Z(n335) );
  XNOR2_X1 U395 ( .A(KEYINPUT83), .B(KEYINPUT22), .ZN(n334) );
  XOR2_X1 U396 ( .A(n335), .B(n334), .Z(n336) );
  XNOR2_X1 U397 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n340), .B(KEYINPUT2), .ZN(n443) );
  XNOR2_X1 U399 ( .A(G148GAT), .B(G106GAT), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n341), .B(G78GAT), .ZN(n366) );
  XNOR2_X1 U401 ( .A(n443), .B(n366), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n466) );
  XNOR2_X1 U403 ( .A(G183GAT), .B(G211GAT), .ZN(n344) );
  XOR2_X1 U404 ( .A(n344), .B(G8GAT), .Z(n395) );
  XNOR2_X1 U405 ( .A(n395), .B(n345), .ZN(n361) );
  XOR2_X1 U406 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n355) );
  XOR2_X1 U407 ( .A(KEYINPUT73), .B(G176GAT), .Z(n347) );
  XNOR2_X1 U408 ( .A(G92GAT), .B(G204GAT), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n348), .B(G64GAT), .ZN(n374) );
  INV_X1 U411 ( .A(n374), .ZN(n349) );
  NAND2_X1 U412 ( .A1(n350), .A2(n349), .ZN(n353) );
  INV_X1 U413 ( .A(n350), .ZN(n351) );
  NAND2_X1 U414 ( .A1(n351), .A2(n374), .ZN(n352) );
  NAND2_X1 U415 ( .A1(n353), .A2(n352), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n359) );
  AND2_X1 U418 ( .A1(G226GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n460) );
  INV_X1 U421 ( .A(n460), .ZN(n523) );
  XOR2_X1 U422 ( .A(KEYINPUT13), .B(KEYINPUT69), .Z(n363) );
  XNOR2_X1 U423 ( .A(G57GAT), .B(G71GAT), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n396) );
  XOR2_X1 U425 ( .A(KEYINPUT71), .B(n396), .Z(n365) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n294), .B(n366), .ZN(n373) );
  XNOR2_X1 U428 ( .A(G120GAT), .B(n367), .ZN(n371) );
  XOR2_X1 U429 ( .A(KEYINPUT31), .B(KEYINPUT70), .Z(n369) );
  XNOR2_X1 U430 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n582) );
  XNOR2_X1 U433 ( .A(KEYINPUT41), .B(n582), .ZN(n564) );
  XOR2_X1 U434 ( .A(G1GAT), .B(KEYINPUT67), .Z(n398) );
  XOR2_X1 U435 ( .A(G169GAT), .B(G50GAT), .Z(n377) );
  XNOR2_X1 U436 ( .A(G113GAT), .B(G36GAT), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U438 ( .A(n398), .B(n378), .Z(n380) );
  NAND2_X1 U439 ( .A1(G229GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U441 ( .A(n381), .B(KEYINPUT65), .Z(n384) );
  XNOR2_X1 U442 ( .A(n382), .B(KEYINPUT66), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n392) );
  XOR2_X1 U444 ( .A(G197GAT), .B(G22GAT), .Z(n386) );
  XNOR2_X1 U445 ( .A(G141GAT), .B(G15GAT), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U447 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n388) );
  XNOR2_X1 U448 ( .A(G8GAT), .B(KEYINPUT68), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U450 ( .A(n390), .B(n389), .Z(n391) );
  XOR2_X1 U451 ( .A(n392), .B(n391), .Z(n578) );
  INV_X1 U452 ( .A(n578), .ZN(n551) );
  NOR2_X1 U453 ( .A1(n564), .A2(n551), .ZN(n394) );
  XOR2_X1 U454 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n414) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n412) );
  XOR2_X1 U457 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U458 ( .A1(G231GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U460 ( .A(n402), .B(n401), .Z(n410) );
  XOR2_X1 U461 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n404) );
  XNOR2_X1 U462 ( .A(G78GAT), .B(G64GAT), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U464 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n406) );
  XNOR2_X1 U465 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U469 ( .A(n412), .B(n411), .Z(n558) );
  XNOR2_X1 U470 ( .A(KEYINPUT107), .B(n558), .ZN(n571) );
  NOR2_X1 U471 ( .A1(n571), .A2(n544), .ZN(n413) );
  NAND2_X1 U472 ( .A1(n414), .A2(n413), .ZN(n417) );
  INV_X1 U473 ( .A(KEYINPUT47), .ZN(n415) );
  XOR2_X1 U474 ( .A(KEYINPUT36), .B(n544), .Z(n591) );
  NOR2_X1 U475 ( .A1(n558), .A2(n591), .ZN(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT45), .B(KEYINPUT110), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  NAND2_X1 U478 ( .A1(n420), .A2(n551), .ZN(n421) );
  NOR2_X1 U479 ( .A1(n582), .A2(n421), .ZN(n422) );
  NOR2_X1 U480 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U481 ( .A(KEYINPUT48), .B(n424), .ZN(n530) );
  NOR2_X1 U482 ( .A1(n523), .A2(n530), .ZN(n427) );
  XOR2_X1 U483 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n425) );
  XNOR2_X1 U484 ( .A(KEYINPUT54), .B(n425), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n447) );
  XOR2_X1 U486 ( .A(G127GAT), .B(G85GAT), .Z(n429) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(G162GAT), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U489 ( .A(KEYINPUT5), .B(G57GAT), .Z(n431) );
  XNOR2_X1 U490 ( .A(G155GAT), .B(G148GAT), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U492 ( .A(n433), .B(n432), .Z(n438) );
  XOR2_X1 U493 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n435) );
  NAND2_X1 U494 ( .A1(G225GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U495 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U496 ( .A(KEYINPUT87), .B(n436), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U498 ( .A(G1GAT), .B(KEYINPUT88), .Z(n440) );
  XNOR2_X1 U499 ( .A(KEYINPUT86), .B(KEYINPUT4), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U501 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U503 ( .A(n446), .B(n445), .Z(n521) );
  NAND2_X1 U504 ( .A1(n447), .A2(n521), .ZN(n576) );
  NOR2_X1 U505 ( .A1(n466), .A2(n576), .ZN(n448) );
  XOR2_X1 U506 ( .A(KEYINPUT55), .B(n448), .Z(n449) );
  NAND2_X1 U507 ( .A1(n494), .A2(n449), .ZN(n570) );
  NOR2_X1 U508 ( .A1(n561), .A2(n570), .ZN(n452) );
  INV_X1 U509 ( .A(KEYINPUT58), .ZN(n450) );
  NOR2_X1 U510 ( .A1(n551), .A2(n570), .ZN(n455) );
  INV_X1 U511 ( .A(G169GAT), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n453), .B(KEYINPUT120), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n455), .B(n454), .ZN(G1348GAT) );
  XNOR2_X1 U514 ( .A(KEYINPUT101), .B(KEYINPUT38), .ZN(n477) );
  NOR2_X1 U515 ( .A1(n582), .A2(n551), .ZN(n456) );
  XNOR2_X1 U516 ( .A(KEYINPUT74), .B(n456), .ZN(n487) );
  INV_X1 U517 ( .A(n521), .ZN(n489) );
  INV_X1 U518 ( .A(n494), .ZN(n531) );
  NOR2_X1 U519 ( .A1(n523), .A2(n531), .ZN(n457) );
  NOR2_X1 U520 ( .A1(n466), .A2(n457), .ZN(n458) );
  XNOR2_X1 U521 ( .A(n458), .B(KEYINPUT93), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n459), .B(KEYINPUT25), .ZN(n463) );
  XOR2_X1 U523 ( .A(n460), .B(KEYINPUT27), .Z(n465) );
  NAND2_X1 U524 ( .A1(n531), .A2(n466), .ZN(n461) );
  XOR2_X1 U525 ( .A(n461), .B(KEYINPUT26), .Z(n549) );
  INV_X1 U526 ( .A(n549), .ZN(n577) );
  NOR2_X1 U527 ( .A1(n465), .A2(n577), .ZN(n462) );
  NOR2_X1 U528 ( .A1(n463), .A2(n462), .ZN(n464) );
  NOR2_X1 U529 ( .A1(n489), .A2(n464), .ZN(n470) );
  OR2_X1 U530 ( .A1(n521), .A2(n465), .ZN(n548) );
  INV_X1 U531 ( .A(n527), .ZN(n499) );
  NOR2_X1 U532 ( .A1(n548), .A2(n499), .ZN(n532) );
  XNOR2_X1 U533 ( .A(KEYINPUT91), .B(n532), .ZN(n467) );
  NOR2_X1 U534 ( .A1(n494), .A2(n467), .ZN(n468) );
  XNOR2_X1 U535 ( .A(n468), .B(KEYINPUT92), .ZN(n469) );
  INV_X1 U536 ( .A(n558), .ZN(n586) );
  NOR2_X1 U537 ( .A1(n485), .A2(n586), .ZN(n471) );
  XNOR2_X1 U538 ( .A(n471), .B(KEYINPUT99), .ZN(n472) );
  NOR2_X1 U539 ( .A1(n591), .A2(n472), .ZN(n475) );
  AND2_X1 U540 ( .A1(n487), .A2(n519), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(n507) );
  NOR2_X1 U542 ( .A1(n521), .A2(n507), .ZN(n480) );
  XNOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n478) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n482) );
  NAND2_X1 U545 ( .A1(n561), .A2(n586), .ZN(n481) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n483), .B(KEYINPUT80), .ZN(n484) );
  NOR2_X1 U548 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U549 ( .A(KEYINPUT94), .B(n486), .ZN(n510) );
  NAND2_X1 U550 ( .A1(n510), .A2(n487), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n488), .B(KEYINPUT95), .ZN(n498) );
  NAND2_X1 U552 ( .A1(n498), .A2(n489), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n490), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n460), .A2(n498), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n492), .B(KEYINPUT96), .ZN(n493) );
  XNOR2_X1 U557 ( .A(G8GAT), .B(n493), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U559 ( .A1(n498), .A2(n494), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U561 ( .A(G15GAT), .B(n497), .Z(G1326GAT) );
  NAND2_X1 U562 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT98), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G22GAT), .B(n501), .ZN(G1327GAT) );
  NOR2_X1 U565 ( .A1(n523), .A2(n507), .ZN(n502) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n504) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n506) );
  NOR2_X1 U570 ( .A1(n507), .A2(n531), .ZN(n505) );
  XOR2_X1 U571 ( .A(n506), .B(n505), .Z(G1330GAT) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n509) );
  NOR2_X1 U573 ( .A1(n527), .A2(n507), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  NOR2_X1 U575 ( .A1(n578), .A2(n564), .ZN(n520) );
  NAND2_X1 U576 ( .A1(n520), .A2(n510), .ZN(n516) );
  NOR2_X1 U577 ( .A1(n521), .A2(n516), .ZN(n511) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U579 ( .A(KEYINPUT42), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U580 ( .A1(n523), .A2(n516), .ZN(n513) );
  XOR2_X1 U581 ( .A(KEYINPUT106), .B(n513), .Z(n514) );
  XNOR2_X1 U582 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U583 ( .A1(n531), .A2(n516), .ZN(n515) );
  XOR2_X1 U584 ( .A(G71GAT), .B(n515), .Z(G1334GAT) );
  NOR2_X1 U585 ( .A1(n527), .A2(n516), .ZN(n518) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n520), .A2(n519), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n521), .A2(n526), .ZN(n522) );
  XOR2_X1 U590 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U591 ( .A1(n523), .A2(n526), .ZN(n524) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n531), .A2(n526), .ZN(n525) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U595 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT111), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n545), .A2(n578), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT112), .Z(n538) );
  INV_X1 U604 ( .A(n564), .ZN(n536) );
  NAND2_X1 U605 ( .A1(n545), .A2(n536), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n540) );
  XOR2_X1 U607 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n542) );
  NAND2_X1 U610 ( .A1(n545), .A2(n571), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U616 ( .A1(n548), .A2(n530), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n551), .A2(n560), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n557) );
  NOR2_X1 U624 ( .A1(n564), .A2(n560), .ZN(n556) );
  XOR2_X1 U625 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U626 ( .A1(n558), .A2(n560), .ZN(n559) );
  XOR2_X1 U627 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NOR2_X1 U631 ( .A1(n570), .A2(n564), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n566) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(KEYINPUT56), .B(n567), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n574) );
  INV_X1 U638 ( .A(n570), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G183GAT), .B(n575), .ZN(G1350GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n589) );
  NAND2_X1 U644 ( .A1(n589), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n589), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT126), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
  INV_X1 U654 ( .A(n589), .ZN(n590) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

