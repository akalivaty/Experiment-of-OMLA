

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XOR2_X1 U324 ( .A(n329), .B(n328), .Z(n292) );
  XNOR2_X1 U325 ( .A(n330), .B(n292), .ZN(n331) );
  XNOR2_X1 U326 ( .A(n378), .B(KEYINPUT48), .ZN(n379) );
  XNOR2_X1 U327 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U328 ( .A(n380), .B(n379), .ZN(n544) );
  XNOR2_X1 U329 ( .A(KEYINPUT125), .B(n456), .ZN(n588) );
  XNOR2_X1 U330 ( .A(n458), .B(G218GAT), .ZN(n459) );
  XNOR2_X1 U331 ( .A(n460), .B(n459), .ZN(G1355GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT11), .B(G92GAT), .Z(n294) );
  XNOR2_X1 U333 ( .A(G134GAT), .B(G106GAT), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n310) );
  XOR2_X1 U335 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n296) );
  NAND2_X1 U336 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U338 ( .A(n297), .B(KEYINPUT66), .Z(n302) );
  XOR2_X1 U339 ( .A(G29GAT), .B(G43GAT), .Z(n299) );
  XNOR2_X1 U340 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n299), .B(n298), .ZN(n343) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .ZN(n300) );
  XNOR2_X1 U343 ( .A(n300), .B(KEYINPUT81), .ZN(n385) );
  XNOR2_X1 U344 ( .A(n343), .B(n385), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U346 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n304) );
  XOR2_X1 U347 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G85GAT), .Z(n327) );
  XNOR2_X1 U349 ( .A(n419), .B(n327), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n306), .B(n305), .Z(n308) );
  XNOR2_X1 U352 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U354 ( .A(n310), .B(n309), .ZN(n559) );
  XNOR2_X1 U355 ( .A(KEYINPUT36), .B(n559), .ZN(n485) );
  XOR2_X1 U356 ( .A(G92GAT), .B(G64GAT), .Z(n312) );
  XNOR2_X1 U357 ( .A(G204GAT), .B(KEYINPUT78), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U359 ( .A(G176GAT), .B(n313), .Z(n386) );
  XOR2_X1 U360 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n315) );
  NAND2_X1 U361 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n317) );
  INV_X1 U363 ( .A(KEYINPUT74), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n326) );
  INV_X1 U365 ( .A(KEYINPUT72), .ZN(n318) );
  NAND2_X1 U366 ( .A1(KEYINPUT13), .A2(n318), .ZN(n321) );
  INV_X1 U367 ( .A(KEYINPUT13), .ZN(n319) );
  NAND2_X1 U368 ( .A1(n319), .A2(KEYINPUT72), .ZN(n320) );
  NAND2_X1 U369 ( .A1(n321), .A2(n320), .ZN(n323) );
  XNOR2_X1 U370 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n354) );
  XNOR2_X1 U372 ( .A(G106GAT), .B(G78GAT), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n324), .B(G148GAT), .ZN(n418) );
  XNOR2_X1 U374 ( .A(n354), .B(n418), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n332) );
  XOR2_X1 U376 ( .A(G120GAT), .B(G71GAT), .Z(n440) );
  XNOR2_X1 U377 ( .A(n440), .B(n327), .ZN(n330) );
  XOR2_X1 U378 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n329) );
  XNOR2_X1 U379 ( .A(KEYINPUT77), .B(KEYINPUT31), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n386), .B(n333), .ZN(n584) );
  XOR2_X1 U381 ( .A(KEYINPUT41), .B(n584), .Z(n569) );
  INV_X1 U382 ( .A(n569), .ZN(n549) );
  XOR2_X1 U383 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n335) );
  XNOR2_X1 U384 ( .A(G22GAT), .B(G15GAT), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U386 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n337) );
  XNOR2_X1 U387 ( .A(KEYINPUT67), .B(KEYINPUT71), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n350) );
  XOR2_X1 U390 ( .A(G197GAT), .B(G141GAT), .Z(n341) );
  XNOR2_X1 U391 ( .A(G50GAT), .B(G36GAT), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U393 ( .A(G169GAT), .B(G8GAT), .Z(n390) );
  XOR2_X1 U394 ( .A(n342), .B(n390), .Z(n348) );
  XOR2_X1 U395 ( .A(n343), .B(KEYINPUT70), .Z(n345) );
  NAND2_X1 U396 ( .A1(G229GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U398 ( .A(G113GAT), .B(G1GAT), .Z(n410) );
  XNOR2_X1 U399 ( .A(n346), .B(n410), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n580) );
  INV_X1 U402 ( .A(n580), .ZN(n547) );
  NOR2_X1 U403 ( .A1(n549), .A2(n547), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n351), .B(KEYINPUT46), .ZN(n369) );
  XOR2_X1 U405 ( .A(G22GAT), .B(G155GAT), .Z(n423) );
  XOR2_X1 U406 ( .A(G78GAT), .B(n423), .Z(n353) );
  XOR2_X1 U407 ( .A(G15GAT), .B(G127GAT), .Z(n441) );
  XNOR2_X1 U408 ( .A(n441), .B(G211GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U410 ( .A(n354), .B(KEYINPUT82), .Z(n356) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U413 ( .A(n358), .B(n357), .Z(n360) );
  XNOR2_X1 U414 ( .A(G183GAT), .B(G71GAT), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n368) );
  XOR2_X1 U416 ( .A(KEYINPUT15), .B(G64GAT), .Z(n362) );
  XNOR2_X1 U417 ( .A(G1GAT), .B(G8GAT), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U419 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n364) );
  XNOR2_X1 U420 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U422 ( .A(n366), .B(n365), .Z(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n589) );
  NOR2_X1 U424 ( .A1(n369), .A2(n589), .ZN(n370) );
  NAND2_X1 U425 ( .A1(n370), .A2(n559), .ZN(n371) );
  XNOR2_X1 U426 ( .A(n371), .B(KEYINPUT47), .ZN(n377) );
  INV_X1 U427 ( .A(n589), .ZN(n555) );
  NOR2_X1 U428 ( .A1(n485), .A2(n555), .ZN(n372) );
  XNOR2_X1 U429 ( .A(KEYINPUT45), .B(n372), .ZN(n374) );
  INV_X1 U430 ( .A(n584), .ZN(n373) );
  NAND2_X1 U431 ( .A1(n374), .A2(n373), .ZN(n375) );
  NOR2_X1 U432 ( .A1(n375), .A2(n580), .ZN(n376) );
  NOR2_X1 U433 ( .A1(n377), .A2(n376), .ZN(n380) );
  XOR2_X1 U434 ( .A(KEYINPUT64), .B(KEYINPUT113), .Z(n378) );
  XOR2_X1 U435 ( .A(G183GAT), .B(KEYINPUT17), .Z(n382) );
  XNOR2_X1 U436 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n446) );
  XOR2_X1 U438 ( .A(G211GAT), .B(KEYINPUT21), .Z(n384) );
  XNOR2_X1 U439 ( .A(G197GAT), .B(G218GAT), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n430) );
  XNOR2_X1 U441 ( .A(n446), .B(n430), .ZN(n394) );
  XOR2_X1 U442 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n388) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U445 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U446 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n518) );
  NOR2_X1 U449 ( .A1(n544), .A2(n518), .ZN(n396) );
  INV_X1 U450 ( .A(KEYINPUT54), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n417) );
  XOR2_X1 U452 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n398) );
  XNOR2_X1 U453 ( .A(G120GAT), .B(G57GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n416) );
  XOR2_X1 U455 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n400) );
  XNOR2_X1 U456 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n406) );
  XOR2_X1 U458 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n402) );
  XNOR2_X1 U459 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n431) );
  XOR2_X1 U461 ( .A(G134GAT), .B(KEYINPUT0), .Z(n445) );
  XOR2_X1 U462 ( .A(n431), .B(n445), .Z(n404) );
  NAND2_X1 U463 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n414) );
  XOR2_X1 U466 ( .A(G85GAT), .B(G148GAT), .Z(n408) );
  XNOR2_X1 U467 ( .A(G127GAT), .B(G162GAT), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U469 ( .A(n409), .B(G155GAT), .Z(n412) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(n410), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n491) );
  NOR2_X1 U474 ( .A1(n417), .A2(n491), .ZN(n563) );
  XOR2_X1 U475 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U476 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U478 ( .A(n422), .B(G204GAT), .Z(n425) );
  XNOR2_X1 U479 ( .A(n423), .B(KEYINPUT90), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U481 ( .A(KEYINPUT92), .B(KEYINPUT22), .Z(n427) );
  XNOR2_X1 U482 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U484 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n564) );
  XOR2_X1 U487 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n435) );
  XNOR2_X1 U488 ( .A(G169GAT), .B(KEYINPUT89), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U490 ( .A(G176GAT), .B(KEYINPUT87), .Z(n437) );
  XNOR2_X1 U491 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n453) );
  XOR2_X1 U494 ( .A(G190GAT), .B(n440), .Z(n443) );
  XNOR2_X1 U495 ( .A(G113GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U497 ( .A(n444), .B(G99GAT), .Z(n451) );
  XOR2_X1 U498 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U501 ( .A(G43GAT), .B(n449), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n453), .B(n452), .ZN(n567) );
  INV_X1 U504 ( .A(n567), .ZN(n528) );
  NOR2_X1 U505 ( .A1(n564), .A2(n528), .ZN(n455) );
  XNOR2_X1 U506 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n546) );
  NAND2_X1 U508 ( .A1(n563), .A2(n546), .ZN(n456) );
  INV_X1 U509 ( .A(n588), .ZN(n457) );
  NOR2_X1 U510 ( .A1(n485), .A2(n457), .ZN(n460) );
  XNOR2_X1 U511 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n458) );
  INV_X1 U512 ( .A(n491), .ZN(n515) );
  NOR2_X1 U513 ( .A1(n547), .A2(n584), .ZN(n488) );
  INV_X1 U514 ( .A(n559), .ZN(n577) );
  NOR2_X1 U515 ( .A1(n577), .A2(n555), .ZN(n461) );
  XNOR2_X1 U516 ( .A(KEYINPUT16), .B(n461), .ZN(n473) );
  INV_X1 U517 ( .A(n518), .ZN(n494) );
  NAND2_X1 U518 ( .A1(n528), .A2(n494), .ZN(n462) );
  NAND2_X1 U519 ( .A1(n462), .A2(n564), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n463), .B(KEYINPUT99), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n464), .B(KEYINPUT25), .ZN(n466) );
  XOR2_X1 U522 ( .A(n518), .B(KEYINPUT27), .Z(n469) );
  NAND2_X1 U523 ( .A1(n469), .A2(n546), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n515), .A2(n467), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n468), .B(KEYINPUT100), .ZN(n472) );
  XOR2_X1 U527 ( .A(n564), .B(KEYINPUT28), .Z(n499) );
  NAND2_X1 U528 ( .A1(n469), .A2(n491), .ZN(n543) );
  NOR2_X1 U529 ( .A1(n499), .A2(n543), .ZN(n529) );
  XOR2_X1 U530 ( .A(n529), .B(KEYINPUT97), .Z(n470) );
  NAND2_X1 U531 ( .A1(n470), .A2(n567), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n483) );
  NAND2_X1 U533 ( .A1(n473), .A2(n483), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT101), .ZN(n504) );
  NAND2_X1 U535 ( .A1(n488), .A2(n504), .ZN(n480) );
  NOR2_X1 U536 ( .A1(n515), .A2(n480), .ZN(n475) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n475), .Z(n476) );
  XNOR2_X1 U538 ( .A(KEYINPUT34), .B(n476), .ZN(G1324GAT) );
  NOR2_X1 U539 ( .A1(n518), .A2(n480), .ZN(n477) );
  XOR2_X1 U540 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  NOR2_X1 U541 ( .A1(n567), .A2(n480), .ZN(n479) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U543 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  INV_X1 U544 ( .A(n499), .ZN(n524) );
  NOR2_X1 U545 ( .A1(n524), .A2(n480), .ZN(n481) );
  XOR2_X1 U546 ( .A(KEYINPUT102), .B(n481), .Z(n482) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  XOR2_X1 U549 ( .A(KEYINPUT104), .B(KEYINPUT38), .Z(n490) );
  NAND2_X1 U550 ( .A1(n555), .A2(n483), .ZN(n484) );
  NOR2_X1 U551 ( .A1(n485), .A2(n484), .ZN(n487) );
  XNOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n487), .B(n486), .ZN(n514) );
  NAND2_X1 U554 ( .A1(n488), .A2(n514), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n490), .B(n489), .ZN(n500) );
  NAND2_X1 U556 ( .A1(n500), .A2(n491), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n494), .A2(n500), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n497) );
  NAND2_X1 U561 ( .A1(n500), .A2(n528), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(KEYINPUT106), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n502), .ZN(G1331GAT) );
  NAND2_X1 U567 ( .A1(n569), .A2(n547), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(KEYINPUT107), .ZN(n513) );
  NAND2_X1 U569 ( .A1(n504), .A2(n513), .ZN(n510) );
  NOR2_X1 U570 ( .A1(n515), .A2(n510), .ZN(n505) );
  XOR2_X1 U571 ( .A(n505), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U573 ( .A1(n518), .A2(n510), .ZN(n507) );
  XOR2_X1 U574 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U575 ( .A1(n567), .A2(n510), .ZN(n508) );
  XOR2_X1 U576 ( .A(KEYINPUT108), .B(n508), .Z(n509) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(n509), .ZN(G1334GAT) );
  NOR2_X1 U578 ( .A1(n524), .A2(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n515), .A2(n523), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U585 ( .A1(n518), .A2(n523), .ZN(n519) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(n519), .Z(n520) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  NOR2_X1 U588 ( .A1(n567), .A2(n523), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1338GAT) );
  NOR2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n526) );
  XNOR2_X1 U592 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n527), .Z(G1339GAT) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U596 ( .A1(n544), .A2(n530), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n539), .A2(n580), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n531), .B(KEYINPUT114), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n534) );
  NAND2_X1 U601 ( .A1(n539), .A2(n569), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n537) );
  NAND2_X1 U605 ( .A1(n539), .A2(n589), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n538), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U609 ( .A1(n539), .A2(n577), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n542), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n558) );
  NOR2_X1 U614 ( .A1(n547), .A2(n558), .ZN(n548) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n548), .Z(G1344GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n558), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(KEYINPUT53), .B(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n558), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT120), .B(n556), .Z(n557) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(n562), .ZN(G1347GAT) );
  AND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT55), .B(n565), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n576), .A2(n580), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT57), .Z(n571) );
  NAND2_X1 U635 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  NAND2_X1 U639 ( .A1(n589), .A2(n576), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT124), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G183GAT), .B(n575), .ZN(G1350GAT) );
  XNOR2_X1 U642 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1351GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  NAND2_X1 U646 ( .A1(n588), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n588), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(n587), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
endmodule

