

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751;

  AND2_X1 U364 ( .A1(n382), .A2(n381), .ZN(n387) );
  AND2_X1 U365 ( .A1(n359), .A2(n747), .ZN(n377) );
  INV_X1 U366 ( .A(n612), .ZN(n410) );
  XNOR2_X1 U367 ( .A(G110), .B(G104), .ZN(n483) );
  INV_X1 U368 ( .A(KEYINPUT70), .ZN(n513) );
  INV_X1 U369 ( .A(G119), .ZN(n512) );
  XNOR2_X2 U370 ( .A(n558), .B(n552), .ZN(n587) );
  AND2_X4 U371 ( .A1(n343), .A2(n657), .ZN(n712) );
  NAND2_X1 U372 ( .A1(n387), .A2(n388), .ZN(n343) );
  XOR2_X1 U373 ( .A(KEYINPUT96), .B(n506), .Z(n661) );
  XNOR2_X1 U374 ( .A(n593), .B(n592), .ZN(n690) );
  XNOR2_X1 U375 ( .A(n557), .B(KEYINPUT1), .ZN(n589) );
  INV_X1 U376 ( .A(G953), .ZN(n738) );
  NOR2_X2 U377 ( .A1(n397), .A2(n572), .ZN(n573) );
  NOR2_X2 U378 ( .A1(n560), .A2(n410), .ZN(n544) );
  XNOR2_X2 U379 ( .A(n400), .B(KEYINPUT32), .ZN(n747) );
  XNOR2_X2 U380 ( .A(n591), .B(n590), .ZN(n606) );
  OR2_X2 U381 ( .A1(n701), .A2(G902), .ZN(n445) );
  XNOR2_X2 U382 ( .A(n396), .B(G131), .ZN(n486) );
  XNOR2_X2 U383 ( .A(n436), .B(KEYINPUT64), .ZN(n533) );
  XNOR2_X2 U384 ( .A(G143), .B(G128), .ZN(n436) );
  NOR2_X1 U385 ( .A1(n675), .A2(n674), .ZN(n679) );
  INV_X4 U386 ( .A(KEYINPUT69), .ZN(n396) );
  AND2_X1 U387 ( .A1(n360), .A2(n352), .ZN(n388) );
  NAND2_X1 U388 ( .A1(n393), .A2(n615), .ZN(n418) );
  AND2_X1 U389 ( .A1(n631), .A2(n614), .ZN(n615) );
  NOR2_X1 U390 ( .A1(n650), .A2(n750), .ZN(n570) );
  AND2_X1 U391 ( .A1(n411), .A2(n410), .ZN(n636) );
  XNOR2_X1 U392 ( .A(n542), .B(KEYINPUT40), .ZN(n749) );
  XNOR2_X1 U393 ( .A(n599), .B(n598), .ZN(n603) );
  NOR2_X1 U394 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U395 ( .A(n356), .B(KEYINPUT41), .ZN(n673) );
  NAND2_X1 U396 ( .A1(n679), .A2(n676), .ZN(n356) );
  NOR2_X2 U397 ( .A1(n368), .A2(n609), .ZN(n565) );
  XNOR2_X1 U398 ( .A(n564), .B(KEYINPUT38), .ZN(n675) );
  OR2_X1 U399 ( .A1(n527), .A2(n577), .ZN(n368) );
  OR2_X1 U400 ( .A1(n424), .A2(n660), .ZN(n560) );
  XNOR2_X1 U401 ( .A(n365), .B(n364), .ZN(n711) );
  NAND2_X1 U402 ( .A1(n369), .A2(KEYINPUT79), .ZN(n372) );
  XNOR2_X2 U403 ( .A(n344), .B(n345), .ZN(n581) );
  NOR2_X1 U404 ( .A1(n696), .A2(n616), .ZN(n344) );
  XOR2_X1 U405 ( .A(n540), .B(n539), .Z(n345) );
  XNOR2_X2 U406 ( .A(n533), .B(n462), .ZN(n485) );
  XNOR2_X1 U407 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n451) );
  XNOR2_X1 U408 ( .A(n505), .B(n504), .ZN(n506) );
  NAND2_X1 U409 ( .A1(n639), .A2(KEYINPUT44), .ZN(n446) );
  XNOR2_X1 U410 ( .A(n461), .B(n373), .ZN(n498) );
  NAND2_X1 U411 ( .A1(n372), .A2(n371), .ZN(n373) );
  NAND2_X1 U412 ( .A1(n370), .A2(G234), .ZN(n371) );
  XNOR2_X1 U413 ( .A(n429), .B(n428), .ZN(n733) );
  XNOR2_X1 U414 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n428) );
  XNOR2_X1 U415 ( .A(n430), .B(G140), .ZN(n429) );
  INV_X1 U416 ( .A(G125), .ZN(n430) );
  INV_X1 U417 ( .A(G134), .ZN(n462) );
  XNOR2_X1 U418 ( .A(n613), .B(n402), .ZN(n401) );
  INV_X1 U419 ( .A(KEYINPUT100), .ZN(n402) );
  NOR2_X1 U420 ( .A1(n647), .A2(n636), .ZN(n613) );
  INV_X1 U421 ( .A(KEYINPUT76), .ZN(n590) );
  XNOR2_X1 U422 ( .A(n733), .B(n427), .ZN(n502) );
  INV_X1 U423 ( .A(G146), .ZN(n427) );
  NAND2_X1 U424 ( .A1(n386), .A2(KEYINPUT80), .ZN(n385) );
  BUF_X1 U425 ( .A(n690), .Z(n404) );
  NAND2_X1 U426 ( .A1(n712), .A2(G475), .ZN(n435) );
  INV_X1 U427 ( .A(KEYINPUT101), .ZN(n399) );
  XOR2_X1 U428 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n475) );
  NOR2_X1 U429 ( .A1(G953), .A2(G237), .ZN(n520) );
  XNOR2_X1 U430 ( .A(n519), .B(n518), .ZN(n528) );
  XNOR2_X1 U431 ( .A(n517), .B(n516), .ZN(n519) );
  INV_X1 U432 ( .A(KEYINPUT3), .ZN(n516) );
  XNOR2_X1 U433 ( .A(n486), .B(n395), .ZN(n487) );
  INV_X1 U434 ( .A(G137), .ZN(n395) );
  XOR2_X1 U435 ( .A(KEYINPUT4), .B(G146), .Z(n534) );
  XNOR2_X1 U436 ( .A(n420), .B(n532), .ZN(n536) );
  XNOR2_X1 U437 ( .A(n533), .B(n421), .ZN(n420) );
  INV_X1 U438 ( .A(KEYINPUT18), .ZN(n530) );
  NAND2_X1 U439 ( .A1(n375), .A2(n447), .ZN(n374) );
  OR2_X1 U440 ( .A1(n646), .A2(n644), .ZN(n550) );
  AND2_X1 U441 ( .A1(n660), .A2(n661), .ZN(n665) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n726) );
  XNOR2_X1 U443 ( .A(n380), .B(G107), .ZN(n378) );
  INV_X1 U444 ( .A(KEYINPUT88), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n528), .B(n450), .ZN(n725) );
  XNOR2_X1 U446 ( .A(G122), .B(KEYINPUT16), .ZN(n450) );
  XOR2_X1 U447 ( .A(KEYINPUT95), .B(G110), .Z(n501) );
  XNOR2_X1 U448 ( .A(G128), .B(G137), .ZN(n500) );
  XNOR2_X1 U449 ( .A(G119), .B(KEYINPUT71), .ZN(n496) );
  XOR2_X1 U450 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n497) );
  INV_X1 U451 ( .A(KEYINPUT117), .ZN(n458) );
  XNOR2_X1 U452 ( .A(n355), .B(n409), .ZN(n622) );
  XNOR2_X1 U453 ( .A(n465), .B(n468), .ZN(n409) );
  XNOR2_X1 U454 ( .A(n485), .B(n469), .ZN(n355) );
  XNOR2_X1 U455 ( .A(G143), .B(G113), .ZN(n472) );
  BUF_X1 U456 ( .A(n673), .Z(n403) );
  XNOR2_X1 U457 ( .A(n366), .B(n351), .ZN(n541) );
  NAND2_X1 U458 ( .A1(n565), .A2(n367), .ZN(n366) );
  INV_X1 U459 ( .A(n675), .ZN(n367) );
  XNOR2_X1 U460 ( .A(KEYINPUT107), .B(KEYINPUT33), .ZN(n592) );
  NAND2_X1 U461 ( .A1(n606), .A2(n600), .ZN(n593) );
  XNOR2_X1 U462 ( .A(n597), .B(KEYINPUT22), .ZN(n598) );
  NAND2_X1 U463 ( .A1(n557), .A2(n665), .ZN(n609) );
  XOR2_X1 U464 ( .A(KEYINPUT86), .B(n623), .Z(n710) );
  INV_X1 U465 ( .A(KEYINPUT47), .ZN(n407) );
  NAND2_X1 U466 ( .A1(n515), .A2(n514), .ZN(n517) );
  NOR2_X1 U467 ( .A1(G953), .A2(KEYINPUT79), .ZN(n370) );
  NAND2_X1 U468 ( .A1(n738), .A2(G234), .ZN(n369) );
  INV_X1 U469 ( .A(KEYINPUT17), .ZN(n421) );
  INV_X1 U470 ( .A(KEYINPUT44), .ZN(n447) );
  OR2_X1 U471 ( .A1(G237), .A2(G902), .ZN(n538) );
  XOR2_X1 U472 ( .A(G101), .B(KEYINPUT5), .Z(n522) );
  INV_X1 U473 ( .A(G101), .ZN(n484) );
  XOR2_X1 U474 ( .A(KEYINPUT7), .B(G122), .Z(n464) );
  XNOR2_X1 U475 ( .A(G116), .B(G107), .ZN(n463) );
  XNOR2_X1 U476 ( .A(KEYINPUT103), .B(KEYINPUT102), .ZN(n466) );
  XOR2_X1 U477 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n467) );
  XNOR2_X1 U478 ( .A(n476), .B(n398), .ZN(n477) );
  XOR2_X1 U479 ( .A(G122), .B(G104), .Z(n473) );
  INV_X1 U480 ( .A(n653), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n358), .B(n349), .ZN(n507) );
  XNOR2_X1 U482 ( .A(KEYINPUT92), .B(KEYINPUT14), .ZN(n358) );
  NOR2_X1 U483 ( .A1(n567), .A2(n566), .ZN(n676) );
  XNOR2_X1 U484 ( .A(n736), .B(n490), .ZN(n394) );
  XNOR2_X1 U485 ( .A(n449), .B(n537), .ZN(n696) );
  XNOR2_X1 U486 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U487 ( .A(n725), .B(n529), .ZN(n449) );
  INV_X1 U488 ( .A(KEYINPUT45), .ZN(n417) );
  XNOR2_X1 U489 ( .A(n526), .B(n406), .ZN(n527) );
  INV_X1 U490 ( .A(KEYINPUT30), .ZN(n406) );
  XNOR2_X1 U491 ( .A(n482), .B(n481), .ZN(n546) );
  INV_X1 U492 ( .A(KEYINPUT13), .ZN(n480) );
  NAND2_X1 U493 ( .A1(n712), .A2(G472), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n460), .B(n347), .ZN(n364) );
  XNOR2_X1 U495 ( .A(n502), .B(n499), .ZN(n365) );
  NAND2_X1 U496 ( .A1(n459), .A2(n457), .ZN(n456) );
  NAND2_X1 U497 ( .A1(n622), .A2(n458), .ZN(n457) );
  NAND2_X1 U498 ( .A1(n621), .A2(KEYINPUT117), .ZN(n459) );
  NAND2_X1 U499 ( .A1(n712), .A2(G478), .ZN(n620) );
  NAND2_X1 U500 ( .A1(n455), .A2(n454), .ZN(n453) );
  NAND2_X1 U501 ( .A1(n622), .A2(KEYINPUT117), .ZN(n454) );
  NAND2_X1 U502 ( .A1(n621), .A2(n458), .ZN(n455) );
  INV_X1 U503 ( .A(n403), .ZN(n689) );
  INV_X1 U504 ( .A(n553), .ZN(n415) );
  AND2_X1 U505 ( .A1(n664), .A2(n413), .ZN(n412) );
  INV_X1 U506 ( .A(n660), .ZN(n413) );
  XNOR2_X1 U507 ( .A(n608), .B(n607), .ZN(n647) );
  NOR2_X1 U508 ( .A1(n546), .A2(n566), .ZN(n644) );
  NOR2_X1 U509 ( .A1(n610), .A2(n609), .ZN(n611) );
  INV_X1 U510 ( .A(KEYINPUT60), .ZN(n432) );
  INV_X1 U511 ( .A(KEYINPUT56), .ZN(n422) );
  XNOR2_X1 U512 ( .A(n726), .B(n451), .ZN(n529) );
  XOR2_X1 U513 ( .A(n495), .B(n494), .Z(n346) );
  XOR2_X1 U514 ( .A(n497), .B(n496), .Z(n347) );
  AND2_X1 U515 ( .A1(n745), .A2(n447), .ZN(n348) );
  AND2_X1 U516 ( .A1(G234), .A2(G237), .ZN(n349) );
  XNOR2_X1 U517 ( .A(n550), .B(KEYINPUT106), .ZN(n678) );
  AND2_X1 U518 ( .A1(n419), .A2(n654), .ZN(n350) );
  XOR2_X1 U519 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n351) );
  INV_X1 U520 ( .A(KEYINPUT80), .ZN(n389) );
  XNOR2_X1 U521 ( .A(n394), .B(n529), .ZN(n701) );
  NAND2_X1 U522 ( .A1(KEYINPUT2), .A2(n616), .ZN(n352) );
  INV_X1 U523 ( .A(n492), .ZN(n386) );
  AND2_X1 U524 ( .A1(n456), .A2(n710), .ZN(n353) );
  AND2_X1 U525 ( .A1(n453), .A2(n710), .ZN(n354) );
  INV_X1 U526 ( .A(KEYINPUT34), .ZN(n444) );
  NAND2_X1 U527 ( .A1(G210), .A2(n712), .ZN(n699) );
  NOR2_X2 U528 ( .A1(n603), .A2(n600), .ZN(n414) );
  NAND2_X1 U529 ( .A1(n748), .A2(n749), .ZN(n549) );
  XNOR2_X2 U530 ( .A(n547), .B(n548), .ZN(n748) );
  INV_X1 U531 ( .A(n443), .ZN(n610) );
  XNOR2_X2 U532 ( .A(n588), .B(KEYINPUT0), .ZN(n443) );
  NAND2_X1 U533 ( .A1(n401), .A2(n678), .ZN(n614) );
  NAND2_X1 U534 ( .A1(n362), .A2(n386), .ZN(n361) );
  XNOR2_X1 U535 ( .A(n357), .B(KEYINPUT93), .ZN(n509) );
  NAND2_X1 U536 ( .A1(n508), .A2(G902), .ZN(n357) );
  INV_X1 U537 ( .A(n577), .ZN(n425) );
  NAND2_X1 U538 ( .A1(n589), .A2(n665), .ZN(n591) );
  NOR2_X1 U539 ( .A1(n745), .A2(n446), .ZN(n359) );
  NAND2_X1 U540 ( .A1(n361), .A2(n389), .ZN(n360) );
  INV_X1 U541 ( .A(n737), .ZN(n362) );
  XNOR2_X2 U542 ( .A(n363), .B(n346), .ZN(n660) );
  NOR2_X1 U543 ( .A1(n711), .A2(G902), .ZN(n363) );
  NAND2_X1 U544 ( .A1(n376), .A2(n374), .ZN(n393) );
  NAND2_X1 U545 ( .A1(n747), .A2(n639), .ZN(n375) );
  NOR2_X1 U546 ( .A1(n377), .A2(n348), .ZN(n376) );
  XNOR2_X1 U547 ( .A(n483), .B(n484), .ZN(n379) );
  AND2_X1 U548 ( .A1(n414), .A2(n563), .ZN(n605) );
  NAND2_X1 U549 ( .A1(n443), .A2(n596), .ZN(n599) );
  NAND2_X1 U550 ( .A1(n610), .A2(KEYINPUT34), .ZN(n440) );
  NAND2_X1 U551 ( .A1(n443), .A2(n444), .ZN(n442) );
  NAND2_X1 U552 ( .A1(n721), .A2(n389), .ZN(n381) );
  NAND2_X1 U553 ( .A1(n384), .A2(n383), .ZN(n382) );
  NOR2_X1 U554 ( .A1(n737), .A2(n385), .ZN(n383) );
  INV_X1 U555 ( .A(n721), .ZN(n384) );
  NOR2_X1 U556 ( .A1(n721), .A2(n737), .ZN(n655) );
  XNOR2_X1 U557 ( .A(n390), .B(KEYINPUT118), .ZN(G63) );
  NAND2_X1 U558 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U559 ( .A1(n620), .A2(n354), .ZN(n391) );
  NAND2_X1 U560 ( .A1(n452), .A2(n353), .ZN(n392) );
  XNOR2_X1 U561 ( .A(n426), .B(n625), .ZN(n626) );
  XNOR2_X1 U562 ( .A(n435), .B(n709), .ZN(n434) );
  NAND2_X1 U563 ( .A1(n673), .A2(n415), .ZN(n547) );
  NAND2_X1 U564 ( .A1(n440), .A2(n595), .ZN(n439) );
  NAND2_X1 U565 ( .A1(n434), .A2(n710), .ZN(n433) );
  NAND2_X1 U566 ( .A1(n570), .A2(n571), .ZN(n397) );
  XNOR2_X1 U567 ( .A(n486), .B(n399), .ZN(n398) );
  XNOR2_X1 U568 ( .A(n487), .B(n534), .ZN(n405) );
  NAND2_X1 U569 ( .A1(n414), .A2(n412), .ZN(n400) );
  XNOR2_X1 U570 ( .A(n611), .B(KEYINPUT98), .ZN(n411) );
  NOR2_X1 U571 ( .A1(n690), .A2(n442), .ZN(n441) );
  NOR2_X1 U572 ( .A1(n441), .A2(n439), .ZN(n438) );
  XNOR2_X2 U573 ( .A(n445), .B(G469), .ZN(n557) );
  NAND2_X1 U574 ( .A1(n438), .A2(n437), .ZN(n448) );
  XNOR2_X2 U575 ( .A(n405), .B(n485), .ZN(n736) );
  XNOR2_X2 U576 ( .A(n617), .B(KEYINPUT82), .ZN(n737) );
  NAND2_X1 U577 ( .A1(n408), .A2(n407), .ZN(n431) );
  INV_X1 U578 ( .A(n554), .ZN(n408) );
  XNOR2_X1 U579 ( .A(n431), .B(KEYINPUT74), .ZN(n556) );
  XNOR2_X2 U580 ( .A(n491), .B(KEYINPUT87), .ZN(n616) );
  NAND2_X1 U581 ( .A1(n416), .A2(n350), .ZN(n617) );
  XNOR2_X1 U582 ( .A(n573), .B(KEYINPUT48), .ZN(n416) );
  NOR2_X1 U583 ( .A1(n543), .A2(n674), .ZN(n526) );
  XNOR2_X1 U584 ( .A(n525), .B(G472), .ZN(n543) );
  XNOR2_X2 U585 ( .A(n418), .B(n417), .ZN(n721) );
  NOR2_X2 U586 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U587 ( .A(n423), .B(n422), .ZN(G51) );
  NAND2_X1 U588 ( .A1(n700), .A2(n710), .ZN(n423) );
  NAND2_X1 U589 ( .A1(n661), .A2(n425), .ZN(n424) );
  NAND2_X1 U590 ( .A1(n642), .A2(n678), .ZN(n554) );
  NOR2_X2 U591 ( .A1(n553), .A2(n587), .ZN(n642) );
  XNOR2_X1 U592 ( .A(n433), .B(n432), .ZN(G60) );
  NAND2_X1 U593 ( .A1(n690), .A2(KEYINPUT34), .ZN(n437) );
  XNOR2_X2 U594 ( .A(n448), .B(KEYINPUT35), .ZN(n745) );
  INV_X1 U595 ( .A(n620), .ZN(n452) );
  XOR2_X1 U596 ( .A(n501), .B(n500), .Z(n460) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n528), .B(n523), .ZN(n524) );
  XNOR2_X1 U599 ( .A(n736), .B(n524), .ZN(n624) );
  INV_X1 U600 ( .A(n594), .ZN(n595) );
  INV_X1 U601 ( .A(KEYINPUT65), .ZN(n597) );
  XNOR2_X1 U602 ( .A(n480), .B(G475), .ZN(n481) );
  XNOR2_X1 U603 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U604 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U605 ( .A(n630), .B(n629), .ZN(G57) );
  XNOR2_X1 U606 ( .A(KEYINPUT105), .B(G478), .ZN(n471) );
  XOR2_X1 U607 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n461) );
  NAND2_X1 U608 ( .A1(n498), .A2(G217), .ZN(n469) );
  XNOR2_X1 U609 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U610 ( .A(n467), .B(n466), .ZN(n468) );
  NOR2_X1 U611 ( .A1(G902), .A2(n622), .ZN(n470) );
  XNOR2_X1 U612 ( .A(n471), .B(n470), .ZN(n566) );
  XNOR2_X1 U613 ( .A(n473), .B(n472), .ZN(n479) );
  NAND2_X1 U614 ( .A1(G214), .A2(n520), .ZN(n474) );
  XNOR2_X1 U615 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U616 ( .A(n477), .B(n502), .ZN(n478) );
  XOR2_X1 U617 ( .A(n479), .B(n478), .Z(n708) );
  NOR2_X1 U618 ( .A1(G902), .A2(n708), .ZN(n482) );
  AND2_X1 U619 ( .A1(n566), .A2(n546), .ZN(n646) );
  XOR2_X1 U620 ( .A(G140), .B(KEYINPUT94), .Z(n489) );
  NAND2_X1 U621 ( .A1(G227), .A2(n738), .ZN(n488) );
  XNOR2_X1 U622 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U623 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n495) );
  XNOR2_X2 U624 ( .A(G902), .B(KEYINPUT15), .ZN(n491) );
  INV_X1 U625 ( .A(n616), .ZN(n492) );
  NAND2_X1 U626 ( .A1(n492), .A2(G234), .ZN(n493) );
  XNOR2_X1 U627 ( .A(n493), .B(KEYINPUT20), .ZN(n503) );
  NAND2_X1 U628 ( .A1(n503), .A2(G217), .ZN(n494) );
  NAND2_X1 U629 ( .A1(n498), .A2(G221), .ZN(n499) );
  XOR2_X1 U630 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n505) );
  NAND2_X1 U631 ( .A1(n503), .A2(G221), .ZN(n504) );
  XNOR2_X1 U632 ( .A(KEYINPUT75), .B(n507), .ZN(n508) );
  NAND2_X1 U633 ( .A1(G952), .A2(n508), .ZN(n688) );
  NOR2_X1 U634 ( .A1(G953), .A2(n688), .ZN(n585) );
  NAND2_X1 U635 ( .A1(n509), .A2(G953), .ZN(n583) );
  NOR2_X1 U636 ( .A1(G900), .A2(n583), .ZN(n510) );
  NOR2_X1 U637 ( .A1(n585), .A2(n510), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G214), .A2(n538), .ZN(n511) );
  XNOR2_X1 U639 ( .A(KEYINPUT91), .B(n511), .ZN(n674) );
  NAND2_X1 U640 ( .A1(KEYINPUT70), .A2(n512), .ZN(n515) );
  NAND2_X1 U641 ( .A1(n513), .A2(G119), .ZN(n514) );
  XNOR2_X1 U642 ( .A(G116), .B(G113), .ZN(n518) );
  NAND2_X1 U643 ( .A1(n520), .A2(G210), .ZN(n521) );
  XNOR2_X1 U644 ( .A(n522), .B(n521), .ZN(n523) );
  NOR2_X1 U645 ( .A1(n624), .A2(G902), .ZN(n525) );
  NAND2_X1 U646 ( .A1(G224), .A2(n738), .ZN(n531) );
  XNOR2_X1 U647 ( .A(n534), .B(G125), .ZN(n535) );
  XOR2_X1 U648 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n540) );
  NAND2_X1 U649 ( .A1(G210), .A2(n538), .ZN(n539) );
  INV_X1 U650 ( .A(n581), .ZN(n564) );
  AND2_X1 U651 ( .A1(n646), .A2(n541), .ZN(n653) );
  NAND2_X1 U652 ( .A1(n541), .A2(n644), .ZN(n542) );
  XOR2_X1 U653 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n548) );
  INV_X1 U654 ( .A(n543), .ZN(n612) );
  XNOR2_X1 U655 ( .A(KEYINPUT28), .B(n544), .ZN(n545) );
  NAND2_X1 U656 ( .A1(n545), .A2(n557), .ZN(n553) );
  INV_X1 U657 ( .A(n546), .ZN(n567) );
  XNOR2_X1 U658 ( .A(n549), .B(KEYINPUT46), .ZN(n572) );
  NOR2_X2 U659 ( .A1(n581), .A2(n674), .ZN(n558) );
  XOR2_X1 U660 ( .A(KEYINPUT77), .B(KEYINPUT19), .Z(n551) );
  XNOR2_X1 U661 ( .A(KEYINPUT66), .B(n551), .ZN(n552) );
  NAND2_X1 U662 ( .A1(n554), .A2(KEYINPUT47), .ZN(n555) );
  AND2_X1 U663 ( .A1(n556), .A2(n555), .ZN(n571) );
  BUF_X1 U664 ( .A(n589), .Z(n664) );
  INV_X1 U665 ( .A(n664), .ZN(n563) );
  XNOR2_X1 U666 ( .A(n410), .B(KEYINPUT6), .ZN(n600) );
  AND2_X1 U667 ( .A1(n644), .A2(n600), .ZN(n579) );
  NAND2_X1 U668 ( .A1(n579), .A2(n558), .ZN(n559) );
  XOR2_X1 U669 ( .A(KEYINPUT36), .B(n561), .Z(n562) );
  NOR2_X1 U670 ( .A1(n563), .A2(n562), .ZN(n650) );
  NAND2_X1 U671 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U672 ( .A1(n567), .A2(n566), .ZN(n594) );
  NOR2_X1 U673 ( .A1(n568), .A2(n594), .ZN(n569) );
  XNOR2_X1 U674 ( .A(n569), .B(KEYINPUT108), .ZN(n750) );
  NOR2_X1 U675 ( .A1(n660), .A2(n664), .ZN(n601) );
  INV_X1 U676 ( .A(n661), .ZN(n574) );
  NOR2_X1 U677 ( .A1(n674), .A2(n574), .ZN(n575) );
  NAND2_X1 U678 ( .A1(n601), .A2(n575), .ZN(n576) );
  NOR2_X1 U679 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U680 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U681 ( .A(KEYINPUT43), .B(n580), .ZN(n582) );
  NAND2_X1 U682 ( .A1(n582), .A2(n581), .ZN(n654) );
  NOR2_X1 U683 ( .A1(G898), .A2(n583), .ZN(n584) );
  NOR2_X1 U684 ( .A1(n585), .A2(n584), .ZN(n586) );
  AND2_X1 U685 ( .A1(n661), .A2(n676), .ZN(n596) );
  INV_X1 U686 ( .A(n601), .ZN(n602) );
  NOR2_X1 U687 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n604), .A2(n410), .ZN(n639) );
  NAND2_X1 U689 ( .A1(n660), .A2(n605), .ZN(n631) );
  XOR2_X1 U690 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n608) );
  AND2_X1 U691 ( .A1(n606), .A2(n612), .ZN(n670) );
  NAND2_X1 U692 ( .A1(n670), .A2(n443), .ZN(n607) );
  NOR2_X1 U693 ( .A1(n617), .A2(n721), .ZN(n618) );
  NAND2_X1 U694 ( .A1(KEYINPUT2), .A2(n618), .ZN(n657) );
  INV_X1 U695 ( .A(n622), .ZN(n621) );
  NOR2_X1 U696 ( .A1(G952), .A2(n738), .ZN(n623) );
  XOR2_X1 U697 ( .A(n624), .B(KEYINPUT62), .Z(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n710), .ZN(n630) );
  XOR2_X1 U699 ( .A(KEYINPUT110), .B(KEYINPUT84), .Z(n628) );
  INV_X1 U700 ( .A(KEYINPUT63), .ZN(n627) );
  XNOR2_X1 U701 ( .A(G101), .B(n631), .ZN(G3) );
  NAND2_X1 U702 ( .A1(n636), .A2(n644), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(G104), .ZN(G6) );
  XOR2_X1 U704 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n634) );
  XNOR2_X1 U705 ( .A(G107), .B(KEYINPUT111), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(n635) );
  XOR2_X1 U707 ( .A(KEYINPUT26), .B(n635), .Z(n638) );
  NAND2_X1 U708 ( .A1(n636), .A2(n646), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(G9) );
  XNOR2_X1 U710 ( .A(G110), .B(n639), .ZN(G12) );
  XOR2_X1 U711 ( .A(G128), .B(KEYINPUT29), .Z(n641) );
  NAND2_X1 U712 ( .A1(n642), .A2(n646), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(G30) );
  NAND2_X1 U714 ( .A1(n642), .A2(n644), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(G146), .ZN(G48) );
  NAND2_X1 U716 ( .A1(n647), .A2(n644), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(G113), .ZN(G15) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n648), .B(KEYINPUT114), .ZN(n649) );
  XNOR2_X1 U720 ( .A(G116), .B(n649), .ZN(G18) );
  XOR2_X1 U721 ( .A(KEYINPUT37), .B(KEYINPUT115), .Z(n652) );
  XNOR2_X1 U722 ( .A(G125), .B(n650), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(G27) );
  XOR2_X1 U724 ( .A(G134), .B(n653), .Z(G36) );
  XNOR2_X1 U725 ( .A(G140), .B(n654), .ZN(G42) );
  OR2_X1 U726 ( .A1(KEYINPUT2), .A2(n655), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U728 ( .A(KEYINPUT81), .B(n658), .ZN(n659) );
  NOR2_X1 U729 ( .A1(G953), .A2(n659), .ZN(n694) );
  NOR2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT49), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n410), .A2(n663), .ZN(n668) );
  NOR2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n666), .B(KEYINPUT50), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U737 ( .A(KEYINPUT51), .B(n671), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n403), .A2(n672), .ZN(n685) );
  INV_X1 U739 ( .A(n404), .ZN(n683) );
  NAND2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n677) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U746 ( .A(KEYINPUT52), .B(n686), .Z(n687) );
  NOR2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n404), .A2(n689), .ZN(n691) );
  NOR2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U751 ( .A(KEYINPUT53), .B(n695), .Z(G75) );
  XNOR2_X1 U752 ( .A(n696), .B(KEYINPUT54), .ZN(n697) );
  XNOR2_X1 U753 ( .A(n697), .B(KEYINPUT55), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n699), .B(n698), .ZN(n700) );
  INV_X1 U755 ( .A(n710), .ZN(n715) );
  XOR2_X1 U756 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n703) );
  XNOR2_X1 U757 ( .A(n701), .B(KEYINPUT116), .ZN(n702) );
  XNOR2_X1 U758 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U759 ( .A1(n712), .A2(G469), .ZN(n704) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U761 ( .A1(n715), .A2(n706), .ZN(G54) );
  XOR2_X1 U762 ( .A(KEYINPUT59), .B(KEYINPUT85), .Z(n707) );
  XOR2_X1 U763 ( .A(n711), .B(KEYINPUT119), .Z(n714) );
  NAND2_X1 U764 ( .A1(n712), .A2(G217), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n714), .B(n713), .ZN(n716) );
  NOR2_X1 U766 ( .A1(n716), .A2(n715), .ZN(G66) );
  NAND2_X1 U767 ( .A1(G224), .A2(G953), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n717), .B(KEYINPUT120), .ZN(n718) );
  XNOR2_X1 U769 ( .A(KEYINPUT61), .B(n718), .ZN(n719) );
  NAND2_X1 U770 ( .A1(n719), .A2(G898), .ZN(n720) );
  XNOR2_X1 U771 ( .A(KEYINPUT121), .B(n720), .ZN(n724) );
  NOR2_X1 U772 ( .A1(G953), .A2(n721), .ZN(n722) );
  XNOR2_X1 U773 ( .A(n722), .B(KEYINPUT122), .ZN(n723) );
  NOR2_X1 U774 ( .A1(n724), .A2(n723), .ZN(n732) );
  XOR2_X1 U775 ( .A(n726), .B(n725), .Z(n727) );
  XNOR2_X1 U776 ( .A(KEYINPUT123), .B(n727), .ZN(n729) );
  NOR2_X1 U777 ( .A1(G898), .A2(n738), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U779 ( .A(KEYINPUT124), .B(n730), .Z(n731) );
  XNOR2_X1 U780 ( .A(n732), .B(n731), .ZN(G69) );
  XNOR2_X1 U781 ( .A(n733), .B(KEYINPUT126), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(KEYINPUT125), .ZN(n735) );
  XNOR2_X1 U783 ( .A(n736), .B(n735), .ZN(n740) );
  XNOR2_X1 U784 ( .A(n740), .B(n737), .ZN(n739) );
  NAND2_X1 U785 ( .A1(n739), .A2(n738), .ZN(n744) );
  XNOR2_X1 U786 ( .A(G227), .B(n740), .ZN(n741) );
  NAND2_X1 U787 ( .A1(n741), .A2(G900), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(G953), .ZN(n743) );
  NAND2_X1 U789 ( .A1(n744), .A2(n743), .ZN(G72) );
  XNOR2_X1 U790 ( .A(n745), .B(G122), .ZN(n746) );
  XNOR2_X1 U791 ( .A(n746), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U792 ( .A(n747), .B(G119), .ZN(G21) );
  XNOR2_X1 U793 ( .A(G137), .B(n748), .ZN(G39) );
  XNOR2_X1 U794 ( .A(n749), .B(G131), .ZN(G33) );
  XNOR2_X1 U795 ( .A(G143), .B(KEYINPUT113), .ZN(n751) );
  XNOR2_X1 U796 ( .A(n751), .B(n750), .ZN(G45) );
endmodule

