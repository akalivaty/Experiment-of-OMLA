//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G77), .ZN(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n206), .A2(new_n207), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n213), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n202), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT66), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n223), .B(new_n224), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AND2_X1   g0031(.A1(new_n229), .A2(new_n230), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n215), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n218), .B(new_n222), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XOR2_X1   g0035(.A(G226), .B(G232), .Z(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n207), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n201), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  AOI21_X1  g0051(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G222), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n253), .B1(new_n254), .B2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT68), .A2(G223), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT68), .A2(G223), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n252), .B1(G77), .B2(new_n253), .C1(new_n255), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n252), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  OAI211_X1 g0065(.A(G1), .B(G13), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n262), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n263), .B1(G226), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n260), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G200), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(G190), .B2(new_n270), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G150), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT8), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n213), .A2(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  XOR2_X1   g0083(.A(new_n283), .B(KEYINPUT69), .Z(new_n284));
  NAND2_X1  g0084(.A1(new_n209), .A2(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n220), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G50), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n288), .B1(new_n212), .B2(G20), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(G50), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n274), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n288), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n284), .B2(new_n285), .ZN(new_n298));
  INV_X1    g0098(.A(new_n295), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n298), .A2(KEYINPUT9), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n273), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT71), .B1(new_n270), .B2(new_n271), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n273), .C1(new_n296), .C2(new_n300), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n270), .A2(new_n308), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n309), .B1(G169), .B2(new_n270), .C1(new_n298), .C2(new_n299), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n294), .A2(G77), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n312), .A2(new_n282), .B1(new_n213), .B2(new_n227), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n280), .B2(new_n275), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n311), .B1(G77), .B2(new_n292), .C1(new_n314), .C2(new_n297), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT70), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G238), .A2(G1698), .ZN(new_n317));
  INV_X1    g0117(.A(G232), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n253), .B(new_n317), .C1(new_n318), .C2(G1698), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n319), .B(new_n252), .C1(G107), .C2(new_n253), .ZN(new_n320));
  INV_X1    g0120(.A(new_n262), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(new_n266), .A3(G274), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n320), .B(new_n322), .C1(new_n228), .C2(new_n267), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G200), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n323), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n323), .A2(G179), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n323), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n327), .B1(new_n316), .B2(new_n330), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n207), .A2(G20), .A3(G33), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT73), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n202), .A2(G20), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n282), .B2(new_n227), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n288), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT11), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n292), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n291), .A2(KEYINPUT12), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n339), .A2(KEYINPUT12), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n294), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT12), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n341), .B1(new_n343), .B2(G68), .ZN(new_n344));
  OAI211_X1 g0144(.A(KEYINPUT11), .B(new_n288), .C1(new_n333), .C2(new_n335), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n338), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n318), .A2(G1698), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n253), .B(new_n347), .C1(G226), .C2(G1698), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n266), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n322), .B1(new_n267), .B2(new_n226), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT13), .B1(new_n350), .B2(new_n352), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n346), .B1(new_n357), .B2(new_n271), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n356), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n359), .A2(KEYINPUT72), .A3(new_n325), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT72), .B1(new_n359), .B2(new_n325), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(G169), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(KEYINPUT14), .B1(new_n357), .B2(G179), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n329), .B1(new_n355), .B2(new_n356), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n365), .A2(KEYINPUT74), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT74), .B1(new_n365), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n346), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n307), .A2(new_n310), .A3(new_n331), .A4(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n292), .A2(new_n280), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n280), .B2(new_n294), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G58), .A2(G68), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n203), .A2(new_n205), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n275), .A2(G159), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n253), .B2(G20), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n264), .A2(KEYINPUT75), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G33), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT3), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n380), .A2(G20), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n381), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n379), .B1(new_n392), .B2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n288), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n384), .A2(new_n386), .A3(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n388), .A2(G33), .ZN(new_n397));
  AOI21_X1  g0197(.A(G20), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n202), .B1(new_n398), .B2(new_n380), .ZN(new_n399));
  INV_X1    g0199(.A(new_n397), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT75), .B(G33), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(KEYINPUT3), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT7), .B1(new_n402), .B2(G20), .ZN(new_n403));
  AOI211_X1 g0203(.A(new_n395), .B(new_n379), .C1(new_n399), .C2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n374), .B1(new_n394), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT76), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n379), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n396), .A2(new_n397), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(new_n380), .A3(new_n213), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G68), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n398), .A2(new_n380), .ZN(new_n412));
  OAI211_X1 g0212(.A(KEYINPUT16), .B(new_n408), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT3), .B1(new_n384), .B2(new_n386), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n390), .B1(new_n414), .B2(new_n383), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n202), .B1(new_n415), .B2(new_n381), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n395), .B1(new_n416), .B2(new_n379), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n413), .A2(new_n288), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(KEYINPUT76), .A3(new_n374), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n322), .B1(new_n267), .B2(new_n318), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  MUX2_X1   g0221(.A(G223), .B(G226), .S(G1698), .Z(new_n422));
  AOI22_X1  g0222(.A1(new_n402), .A2(new_n422), .B1(G33), .B2(G87), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n423), .B2(new_n266), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n424), .A2(new_n308), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(G169), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n407), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT18), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n402), .A2(new_n422), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n266), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(G200), .B1(new_n432), .B2(new_n420), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n421), .B(G190), .C1(new_n266), .C2(new_n423), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(new_n418), .A3(new_n374), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n435), .A2(new_n418), .A3(new_n438), .A4(new_n374), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n407), .A2(new_n441), .A3(new_n419), .A4(new_n427), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n429), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n372), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT5), .ZN(new_n446));
  AOI211_X1 g0246(.A(G1), .B(new_n445), .C1(new_n446), .C2(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(G41), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n447), .A2(G274), .A3(new_n266), .A4(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n445), .A2(G1), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(KEYINPUT5), .B2(new_n265), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n266), .B(G264), .C1(new_n452), .C2(new_n448), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  MUX2_X1   g0254(.A(G250), .B(G257), .S(G1698), .Z(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(new_n396), .A3(new_n397), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n387), .A2(G294), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n266), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n458), .A2(new_n459), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT85), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n460), .B2(new_n461), .ZN(new_n465));
  OAI21_X1  g0265(.A(G169), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n453), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n458), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n450), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n466), .B1(new_n308), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n397), .A2(new_n382), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n472));
  INV_X1    g0272(.A(G87), .ZN(new_n473));
  NOR4_X1   g0273(.A1(new_n471), .A2(new_n472), .A3(G20), .A4(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n396), .A2(new_n213), .A3(G87), .A4(new_n397), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT22), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT80), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(KEYINPUT80), .A3(KEYINPUT22), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT82), .ZN(new_n481));
  INV_X1    g0281(.A(G107), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G20), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT23), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n387), .A2(G116), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(G20), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT83), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n485), .B(KEYINPUT83), .C1(G20), .C2(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n480), .A2(new_n481), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n481), .B1(new_n480), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT24), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n479), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT80), .B1(new_n475), .B2(KEYINPUT22), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n495), .A2(new_n474), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n489), .A2(new_n490), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT82), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT24), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n480), .A2(new_n481), .A3(new_n491), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n297), .B1(new_n494), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT25), .B1(new_n339), .B2(new_n482), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n339), .A2(KEYINPUT25), .A3(new_n482), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n212), .A2(G33), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n297), .A2(new_n292), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n505), .A2(new_n506), .B1(new_n509), .B2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n470), .B1(new_n503), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT24), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n288), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n465), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n325), .A3(new_n463), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n469), .A2(new_n271), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n510), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G116), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n287), .A2(new_n220), .B1(G20), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  INV_X1    g0324(.A(G97), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n213), .C1(G33), .C2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT79), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT79), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n523), .A2(new_n529), .A3(new_n526), .A4(KEYINPUT20), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n523), .A2(new_n526), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n528), .B(new_n530), .C1(KEYINPUT20), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n339), .A2(new_n522), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n509), .A2(G116), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n266), .B(G270), .C1(new_n452), .C2(new_n448), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n450), .A2(new_n536), .ZN(new_n537));
  MUX2_X1   g0337(.A(G257), .B(G264), .S(G1698), .Z(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(new_n396), .A3(new_n397), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n471), .A2(G303), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n266), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n535), .A2(new_n542), .A3(KEYINPUT21), .A4(G169), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n533), .B1(new_n508), .B2(new_n522), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT20), .B1(new_n523), .B2(new_n526), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(KEYINPUT79), .B2(new_n527), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n547), .B2(new_n530), .ZN(new_n548));
  OAI21_X1  g0348(.A(G169), .B1(new_n537), .B2(new_n541), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n537), .A2(new_n541), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n535), .A2(G179), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n543), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n312), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n292), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n402), .A2(new_n213), .A3(G68), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n349), .B2(new_n213), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n473), .A2(new_n525), .A3(new_n482), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n558), .A2(new_n559), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n555), .B1(new_n562), .B2(new_n288), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n312), .B2(new_n508), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n451), .A2(G250), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n451), .A2(new_n261), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n266), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G238), .A2(G1698), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n228), .B2(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n396), .A3(new_n397), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n570), .A2(new_n486), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n308), .B(new_n567), .C1(new_n571), .C2(new_n266), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n266), .B1(new_n570), .B2(new_n486), .ZN(new_n573));
  INV_X1    g0373(.A(new_n567), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n329), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n572), .A2(KEYINPUT78), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT78), .B1(new_n572), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n564), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n508), .A2(new_n473), .ZN(new_n579));
  AOI211_X1 g0379(.A(new_n555), .B(new_n579), .C1(new_n562), .C2(new_n288), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n573), .A2(new_n574), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G190), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n582), .C1(new_n271), .C2(new_n581), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n551), .A2(G190), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n584), .B(new_n548), .C1(new_n271), .C2(new_n551), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n553), .A2(new_n578), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G257), .B(new_n266), .C1(new_n452), .C2(new_n448), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n450), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n228), .A2(G1698), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n396), .A2(new_n397), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT77), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT4), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n402), .A2(KEYINPUT77), .A3(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n589), .A2(KEYINPUT4), .B1(G250), .B2(G1698), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n524), .B1(new_n595), .B2(new_n471), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n588), .B1(new_n598), .B2(new_n252), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n482), .A2(KEYINPUT6), .A3(G97), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n525), .A2(new_n482), .ZN(new_n602));
  NOR2_X1   g0402(.A1(G97), .A2(G107), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n601), .B1(new_n604), .B2(KEYINPUT6), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n605), .A2(G20), .B1(G77), .B2(new_n275), .ZN(new_n606));
  INV_X1    g0406(.A(new_n392), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n482), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n288), .ZN(new_n609));
  INV_X1    g0409(.A(new_n588), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n596), .B1(new_n592), .B2(new_n593), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(new_n266), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G200), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n292), .A2(G97), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n509), .B2(G97), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n600), .A2(new_n609), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n609), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n329), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n610), .B(new_n308), .C1(new_n611), .C2(new_n266), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n586), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n444), .A2(new_n521), .A3(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n310), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n369), .A2(new_n370), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n316), .A2(new_n330), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n362), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n440), .ZN(new_n628));
  INV_X1    g0428(.A(new_n405), .ZN(new_n629));
  INV_X1    g0429(.A(new_n427), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT18), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n624), .B1(new_n633), .B2(new_n307), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n574), .A2(KEYINPUT86), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT86), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n567), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n635), .B(new_n637), .C1(new_n266), .C2(new_n571), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n329), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(new_n564), .A3(new_n572), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n617), .A2(new_n618), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(new_n619), .A3(new_n578), .A4(new_n583), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n620), .A2(KEYINPUT88), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n617), .A2(new_n618), .A3(new_n646), .A4(new_n619), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n638), .A2(G200), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n580), .A3(new_n582), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n640), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n512), .A2(new_n553), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n620), .A3(new_n616), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n494), .A2(new_n502), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n511), .B1(new_n658), .B2(new_n288), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n659), .B2(new_n519), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n656), .A2(new_n660), .A3(KEYINPUT87), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT87), .B1(new_n656), .B2(new_n660), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n655), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n444), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n634), .B1(new_n664), .B2(new_n665), .ZN(G369));
  NAND2_X1  g0466(.A1(new_n291), .A2(new_n213), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT89), .Z(new_n671));
  INV_X1    g0471(.A(KEYINPUT90), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(G343), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(G343), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n521), .B1(new_n659), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n512), .B2(new_n676), .ZN(new_n678));
  INV_X1    g0478(.A(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n535), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n553), .A3(new_n585), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n553), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n553), .A2(new_n679), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n521), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n515), .A2(new_n510), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n470), .A3(new_n676), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n216), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n559), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n219), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n656), .A2(new_n660), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n649), .B1(new_n648), .B2(new_n652), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n640), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n679), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT29), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT87), .ZN(new_n707));
  INV_X1    g0507(.A(new_n553), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n688), .B2(new_n470), .ZN(new_n709));
  INV_X1    g0509(.A(new_n657), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n520), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n707), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n656), .A2(new_n660), .A3(KEYINPUT87), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n679), .B1(new_n714), .B2(new_n655), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n706), .B1(new_n715), .B2(new_n705), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n512), .A2(new_n520), .A3(new_n622), .A4(new_n676), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT91), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n542), .A2(new_n308), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n468), .A2(new_n581), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n599), .A2(new_n719), .A3(KEYINPUT30), .A4(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n551), .A2(new_n468), .A3(new_n581), .A4(G179), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n612), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n551), .A2(G179), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n612), .A2(new_n725), .A3(new_n469), .A4(new_n638), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n721), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n679), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n718), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI211_X1 g0530(.A(KEYINPUT91), .B(KEYINPUT31), .C1(new_n727), .C2(new_n679), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n728), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT31), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n717), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n716), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n699), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n290), .A2(G20), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G45), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n694), .A2(G1), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n684), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n682), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n213), .A2(new_n325), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n308), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n213), .A2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n271), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n750), .A2(new_n201), .B1(new_n753), .B2(new_n482), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(new_n751), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G159), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n253), .B1(new_n227), .B2(new_n755), .C1(new_n760), .C2(KEYINPUT32), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n748), .A2(new_n752), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n754), .B(new_n761), .C1(G87), .C2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n325), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n207), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n765), .A2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n213), .B1(new_n756), .B2(G190), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n770), .A2(new_n202), .B1(new_n771), .B2(new_n525), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n768), .B(new_n772), .C1(KEYINPUT32), .C2(new_n760), .ZN(new_n773));
  INV_X1    g0573(.A(G322), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n471), .B1(new_n750), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT33), .B(G317), .Z(new_n776));
  INV_X1    g0576(.A(G294), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n770), .A2(new_n776), .B1(new_n777), .B2(new_n771), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n775), .B(new_n778), .C1(G326), .C2(new_n766), .ZN(new_n779));
  INV_X1    g0579(.A(G303), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n762), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n753), .B1(new_n755), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n757), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n781), .B(new_n784), .C1(G329), .C2(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n764), .A2(new_n773), .B1(new_n779), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n220), .B1(G20), .B2(new_n329), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n745), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n788), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n247), .A2(G45), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n216), .A2(new_n409), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT92), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(G45), .C2(new_n697), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n692), .A2(new_n471), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n800), .A2(G355), .B1(new_n522), .B2(new_n692), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n795), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n793), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n682), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n747), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  NAND2_X1  g0607(.A1(new_n316), .A2(new_n679), .ZN(new_n808));
  OAI21_X1  g0608(.A(KEYINPUT94), .B1(new_n626), .B2(new_n676), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT94), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n316), .A2(new_n679), .A3(new_n330), .A4(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n331), .A2(new_n808), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n715), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n745), .B1(new_n814), .B2(new_n739), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n739), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n788), .A2(new_n791), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n753), .A2(new_n473), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G311), .B2(new_n785), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n820), .B1(new_n522), .B2(new_n755), .C1(new_n777), .C2(new_n750), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n471), .B1(new_n771), .B2(new_n525), .C1(new_n482), .C2(new_n762), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n770), .A2(new_n782), .B1(new_n767), .B2(new_n780), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n750), .ZN(new_n825));
  INV_X1    g0625(.A(new_n755), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G143), .A2(new_n825), .B1(new_n826), .B2(G159), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n827), .B1(new_n767), .B2(new_n828), .C1(new_n829), .C2(new_n770), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT34), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n753), .A2(new_n202), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G132), .B2(new_n785), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n207), .B2(new_n762), .ZN(new_n834));
  INV_X1    g0634(.A(new_n771), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n409), .B(new_n834), .C1(G58), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n824), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n745), .B1(G77), .B2(new_n818), .C1(new_n837), .C2(new_n789), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT93), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n792), .B2(new_n813), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n816), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  OR2_X1    g0642(.A1(new_n605), .A2(KEYINPUT35), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n605), .A2(KEYINPUT35), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(G116), .A3(new_n221), .A4(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT36), .Z(new_n846));
  NAND3_X1  g0646(.A1(new_n219), .A2(G77), .A3(new_n375), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n207), .A2(G68), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n212), .B(G13), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n679), .A2(new_n370), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n371), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n371), .A2(new_n851), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n812), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT31), .B1(new_n728), .B2(KEYINPUT99), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(KEYINPUT99), .B2(new_n728), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n717), .A2(new_n856), .A3(new_n734), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n854), .A2(new_n857), .A3(KEYINPUT40), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n436), .B1(new_n629), .B2(new_n630), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n418), .A2(KEYINPUT76), .A3(new_n374), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT76), .B1(new_n418), .B2(new_n374), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT97), .B1(new_n863), .B2(new_n671), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n407), .A2(KEYINPUT97), .A3(new_n419), .A4(new_n671), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n860), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(KEYINPUT98), .A3(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT98), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n407), .A2(new_n419), .A3(new_n671), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT97), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n859), .B1(new_n872), .B2(new_n865), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n436), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n428), .B(new_n877), .C1(new_n864), .C2(new_n866), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n868), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n632), .A2(new_n440), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n872), .A3(new_n865), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n297), .B1(new_n883), .B2(new_n395), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(KEYINPUT95), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n379), .B1(new_n399), .B2(new_n403), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT95), .B(new_n288), .C1(new_n886), .C2(KEYINPUT16), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n413), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n374), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n671), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n427), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n891), .A3(new_n436), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n878), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT96), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n428), .A2(KEYINPUT18), .B1(new_n437), .B2(new_n439), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n895), .B(new_n890), .C1(new_n896), .C2(new_n442), .ZN(new_n897));
  INV_X1    g0697(.A(new_n890), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT96), .B1(new_n443), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n894), .B(KEYINPUT38), .C1(new_n897), .C2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n858), .B1(new_n882), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n854), .A2(new_n857), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n894), .B1(new_n897), .B2(new_n899), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n903), .B1(new_n906), .B2(new_n900), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n902), .B(G330), .C1(KEYINPUT40), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n444), .A2(new_n857), .A3(G330), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT100), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n903), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n443), .A2(new_n898), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n895), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n443), .A2(KEYINPUT96), .A3(new_n898), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n917), .B2(new_n894), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n913), .B1(new_n918), .B2(new_n901), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n921), .A2(new_n444), .A3(new_n857), .A4(new_n902), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n912), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n910), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(KEYINPUT100), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n625), .A2(new_n679), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n882), .A2(new_n901), .A3(KEYINPUT39), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n906), .B2(new_n900), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n926), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n663), .A2(new_n676), .A3(new_n813), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n626), .A2(new_n679), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n906), .A2(new_n900), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n852), .A2(new_n853), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n632), .A2(new_n671), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n930), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n634), .B1(new_n716), .B2(new_n665), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n925), .A2(new_n942), .B1(new_n212), .B2(new_n742), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n925), .A2(new_n942), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n850), .B1(new_n943), .B2(new_n944), .ZN(G367));
  NAND2_X1  g0745(.A1(new_n679), .A2(new_n617), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(new_n616), .A3(new_n620), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n620), .B2(new_n676), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n521), .A2(new_n686), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n620), .B1(new_n512), .B2(new_n947), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n949), .A2(KEYINPUT42), .B1(new_n676), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(KEYINPUT42), .B2(new_n949), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n676), .A2(new_n580), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n640), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT101), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT101), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n652), .A2(new_n953), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n952), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n685), .ZN(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT102), .B1(new_n963), .B2(new_n948), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n963), .A2(KEYINPUT102), .A3(new_n948), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n962), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n693), .B(KEYINPUT41), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n685), .A2(KEYINPUT104), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n690), .A2(new_n948), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT103), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n690), .A2(new_n948), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n971), .A2(new_n972), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n969), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n969), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n973), .A2(new_n980), .A3(new_n977), .A4(new_n975), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n683), .A2(KEYINPUT105), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n687), .B(new_n982), .C1(new_n678), .C2(new_n686), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n683), .A2(KEYINPUT105), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n985), .A2(new_n740), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n968), .B1(new_n987), .B2(new_n740), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n743), .A2(G1), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n965), .B(new_n967), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n798), .A2(new_n243), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n795), .B1(new_n692), .B2(new_n554), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n744), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT106), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n750), .A2(new_n829), .B1(new_n753), .B2(new_n227), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n762), .A2(new_n201), .B1(new_n757), .B2(new_n828), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n771), .A2(new_n202), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n471), .B1(new_n826), .B2(G50), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G143), .A2(new_n766), .B1(new_n769), .B2(G159), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n753), .A2(new_n525), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n750), .A2(new_n780), .B1(new_n755), .B2(new_n782), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(G317), .C2(new_n785), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n763), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT46), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n762), .B2(new_n522), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1006), .B(new_n1008), .C1(new_n777), .C2(new_n770), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT107), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n409), .B1(new_n767), .B2(new_n783), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G107), .B2(new_n835), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1005), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1009), .A2(KEYINPUT107), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1002), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT47), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n788), .B1(new_n1016), .B2(KEYINPUT47), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n994), .B1(new_n1017), .B2(new_n1018), .C1(new_n958), .C2(new_n804), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n990), .A2(new_n1019), .ZN(G387));
  NOR2_X1   g0820(.A1(new_n986), .A2(new_n694), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n740), .B2(new_n985), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n678), .A2(new_n804), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n762), .A2(new_n777), .B1(new_n771), .B2(new_n782), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G317), .A2(new_n825), .B1(new_n826), .B2(G303), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n767), .B2(new_n774), .C1(new_n783), .C2(new_n770), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n753), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G116), .A2(new_n1033), .B1(new_n785), .B2(G326), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1031), .A2(new_n409), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n835), .A2(new_n554), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n770), .B2(new_n281), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n409), .B(new_n1037), .C1(G159), .C2(new_n766), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n762), .A2(new_n227), .B1(new_n757), .B2(new_n829), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT109), .Z(new_n1040));
  NOR2_X1   g0840(.A1(new_n755), .A2(new_n202), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1003), .B(new_n1041), .C1(G50), .C2(new_n825), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n789), .B1(new_n1035), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n695), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n800), .A2(new_n1045), .B1(new_n482), .B2(new_n692), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n240), .A2(G45), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n280), .A2(new_n207), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n695), .B(new_n445), .C1(new_n202), .C2(new_n227), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n798), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1046), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT108), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1055), .A2(new_n794), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n744), .B(new_n1044), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT110), .Z(new_n1058));
  AOI22_X1  g0858(.A1(new_n985), .A2(new_n989), .B1(new_n1023), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1022), .A2(new_n1059), .ZN(G393));
  OAI21_X1  g0860(.A(new_n963), .B1(new_n976), .B2(new_n978), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n973), .A2(new_n685), .A3(new_n977), .A4(new_n975), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n989), .A3(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n825), .A2(G311), .B1(G317), .B2(new_n766), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT52), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n762), .A2(new_n782), .B1(new_n757), .B2(new_n774), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G294), .B2(new_n826), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n771), .A2(new_n522), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n471), .B1(new_n753), .B2(new_n482), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(G303), .C2(new_n769), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1065), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n767), .A2(new_n829), .B1(new_n750), .B2(new_n758), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n819), .B1(G143), .B2(new_n785), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n763), .A2(G68), .B1(new_n826), .B2(new_n280), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n771), .A2(new_n227), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1076), .B(new_n409), .C1(G50), .C2(new_n769), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n789), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n798), .A2(new_n250), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n795), .B1(G97), .B2(new_n692), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n744), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n948), .B2(new_n804), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n987), .A2(new_n693), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n986), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1063), .B(new_n1083), .C1(new_n1084), .C2(new_n1085), .ZN(G390));
  OAI21_X1  g0886(.A(new_n745), .B1(new_n280), .B2(new_n818), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n253), .B(new_n1076), .C1(G87), .C2(new_n763), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n832), .B1(G97), .B2(new_n826), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G116), .A2(new_n825), .B1(new_n785), .B2(G294), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G107), .A2(new_n769), .B1(new_n766), .B2(G283), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(G125), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n253), .B1(new_n757), .B2(new_n1093), .C1(new_n207), .C2(new_n753), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT114), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n762), .A2(new_n829), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1097));
  XNOR2_X1  g0897(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G132), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n750), .A2(new_n1099), .B1(new_n755), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G159), .B2(new_n835), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G128), .A2(new_n766), .B1(new_n769), .B2(G137), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1098), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1092), .B1(new_n1095), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1087), .B1(new_n1105), .B2(new_n788), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n879), .A2(new_n881), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n928), .B(new_n900), .C1(new_n1107), .C2(KEYINPUT38), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n935), .A2(KEYINPUT39), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1106), .B1(new_n1110), .B2(new_n792), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n926), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n882), .B2(new_n901), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n936), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n700), .A2(new_n703), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n676), .A3(new_n813), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(new_n1116), .B2(new_n933), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n812), .A2(new_n737), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n735), .A2(new_n936), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n926), .B1(new_n934), .B2(new_n936), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1118), .B(new_n1120), .C1(new_n1121), .C2(new_n1110), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n932), .B1(new_n715), .B2(new_n813), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1112), .B1(new_n1124), .B2(new_n1114), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n927), .A2(new_n929), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n857), .A2(new_n936), .A3(new_n1119), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n989), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1111), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1116), .A2(new_n1120), .A3(new_n933), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n936), .B1(new_n857), .B2(new_n1119), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n735), .A2(new_n1119), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1114), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT112), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT112), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1135), .A2(new_n1138), .A3(new_n1114), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1128), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1134), .B1(new_n1140), .B2(new_n934), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n909), .A2(KEYINPUT111), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT111), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n444), .A2(new_n857), .A3(new_n1143), .A4(G330), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n634), .B(new_n1145), .C1(new_n716), .C2(new_n665), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1129), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1122), .B(new_n1147), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n693), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1131), .B1(new_n1151), .B2(KEYINPUT113), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(KEYINPUT113), .B2(new_n1151), .ZN(G378));
  INV_X1    g0953(.A(new_n1146), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT120), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT120), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n1157), .A3(new_n1154), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n307), .A2(new_n310), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n671), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n289), .B2(new_n295), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OR3_X1    g0966(.A1(new_n1162), .A2(new_n1163), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n908), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n921), .A2(G330), .A3(new_n902), .A4(new_n1169), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(new_n939), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1174), .A2(KEYINPUT57), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n694), .B1(new_n1159), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT118), .B1(new_n1173), .B2(new_n939), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n930), .A2(new_n937), .A3(new_n938), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT118), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1178), .A2(new_n1179), .A3(new_n1172), .A4(new_n1171), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT117), .B1(new_n1173), .B2(new_n939), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1173), .A2(new_n939), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT117), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT57), .B1(new_n1188), .B2(new_n1159), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1176), .B1(new_n1189), .B2(KEYINPUT121), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT121), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1191), .B(KEYINPUT57), .C1(new_n1188), .C2(new_n1159), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1186), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n989), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT119), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n767), .A2(new_n1093), .B1(new_n771), .B2(new_n829), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1100), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G128), .A2(new_n825), .B1(new_n763), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n828), .B2(new_n755), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1198), .B(new_n1201), .C1(G132), .C2(new_n769), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1033), .A2(G159), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n999), .B1(new_n770), .B2(new_n525), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n825), .A2(G107), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT116), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n402), .A2(G41), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G77), .A2(new_n763), .B1(new_n785), .B2(G283), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n753), .A2(new_n201), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n554), .B2(new_n826), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1209), .B(new_n1216), .C1(G116), .C2(new_n766), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1212), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1208), .A2(new_n1218), .A3(new_n1219), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n788), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n744), .B1(new_n207), .B2(new_n817), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n1169), .C2(new_n792), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1196), .A2(new_n1197), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1130), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1225), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT119), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1193), .A2(new_n1230), .ZN(G375));
  INV_X1    g1031(.A(new_n1141), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1114), .A2(new_n791), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n471), .B1(new_n753), .B2(new_n227), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT122), .Z(new_n1235));
  OAI221_X1 g1035(.A(new_n1036), .B1(new_n767), .B2(new_n777), .C1(new_n522), .C2(new_n770), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n750), .A2(new_n782), .B1(new_n755), .B2(new_n482), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n762), .A2(new_n525), .B1(new_n757), .B2(new_n780), .ZN(new_n1238));
  OR4_X1    g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n767), .A2(new_n1099), .B1(new_n771), .B2(new_n207), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n769), .B2(new_n1199), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n762), .A2(new_n758), .B1(new_n755), .B2(new_n829), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G128), .B2(new_n785), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1214), .B1(G137), .B2(new_n825), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1243), .A3(new_n402), .A4(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n789), .B1(new_n1239), .B2(new_n1245), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n744), .B(new_n1246), .C1(new_n202), .C2(new_n817), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1232), .A2(new_n989), .B1(new_n1233), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n968), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1148), .A2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1232), .A2(new_n1154), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1248), .B1(new_n1250), .B2(new_n1251), .ZN(G381));
  INV_X1    g1052(.A(G375), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1131), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1151), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1022), .A2(new_n806), .A3(new_n841), .A4(new_n1059), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(G387), .A2(new_n1257), .A3(G390), .A4(G381), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1253), .A2(new_n1256), .A3(new_n1258), .ZN(G407));
  NAND3_X1  g1059(.A1(new_n673), .A2(new_n674), .A3(G213), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1253), .A2(new_n1256), .A3(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(G407), .A2(new_n1262), .A3(G213), .ZN(G409));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1230), .B(G378), .C1(new_n1190), .C2(new_n1192), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1188), .A2(new_n1159), .A3(new_n1249), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1174), .A2(KEYINPUT123), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n989), .B1(new_n1174), .B2(KEYINPUT123), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1266), .B(new_n1225), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1256), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1260), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1251), .A2(KEYINPUT60), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n693), .A3(new_n1148), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1251), .A2(KEYINPUT60), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1248), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(new_n841), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n841), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1264), .B1(new_n1272), .B2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1277), .B(new_n1278), .C1(KEYINPUT124), .C2(new_n1260), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1261), .A2(G2897), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1281), .B(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1261), .B1(new_n1265), .B2(new_n1270), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1279), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(KEYINPUT63), .A3(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n990), .A2(new_n1019), .A3(G390), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT125), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(G393), .B(G396), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(G390), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G387), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1290), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1280), .A2(new_n1286), .A3(new_n1289), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1287), .A2(new_n1302), .A3(new_n1288), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1287), .B2(new_n1284), .ZN(new_n1305));
  XOR2_X1   g1105(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1303), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT127), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1299), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1309), .B1(new_n1310), .B2(new_n1297), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1298), .A2(KEYINPUT127), .A3(new_n1299), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1301), .B1(new_n1308), .B2(new_n1313), .ZN(G405));
  OAI211_X1 g1114(.A(new_n1265), .B(new_n1279), .C1(new_n1253), .C2(new_n1255), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1310), .A2(new_n1297), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1255), .B1(new_n1193), .B2(new_n1230), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1265), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1288), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1315), .A2(new_n1316), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1316), .B1(new_n1315), .B2(new_n1319), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(G402));
endmodule


