

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577;

  NOR2_X1 U319 ( .A1(n572), .A2(n575), .ZN(n447) );
  XOR2_X1 U320 ( .A(G29GAT), .B(G43GAT), .Z(n296) );
  NOR2_X1 U321 ( .A1(n535), .A2(n459), .ZN(n460) );
  NOR2_X1 U322 ( .A1(n534), .A2(n514), .ZN(n517) );
  XNOR2_X1 U323 ( .A(n458), .B(KEYINPUT48), .ZN(n535) );
  INV_X1 U324 ( .A(n561), .ZN(n493) );
  NOR2_X1 U325 ( .A1(n518), .A2(n463), .ZN(n365) );
  XOR2_X2 U326 ( .A(n307), .B(n306), .Z(n555) );
  AND2_X1 U327 ( .A1(n567), .A2(n448), .ZN(n449) );
  XNOR2_X1 U328 ( .A(KEYINPUT95), .B(n366), .ZN(n559) );
  AND2_X1 U329 ( .A1(n462), .A2(n461), .ZN(n560) );
  XNOR2_X1 U330 ( .A(n346), .B(n345), .ZN(n518) );
  XOR2_X1 U331 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n287) );
  XOR2_X1 U332 ( .A(n420), .B(n419), .Z(n288) );
  XOR2_X1 U333 ( .A(n443), .B(KEYINPUT101), .Z(n289) );
  XNOR2_X1 U334 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n451) );
  XNOR2_X1 U335 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U336 ( .A(n410), .B(KEYINPUT33), .ZN(n411) );
  XNOR2_X1 U337 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U338 ( .A(n421), .B(n288), .ZN(n422) );
  XNOR2_X1 U339 ( .A(n423), .B(n422), .ZN(n427) );
  INV_X1 U340 ( .A(G183GAT), .ZN(n466) );
  XNOR2_X1 U341 ( .A(n466), .B(KEYINPUT122), .ZN(n467) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n444) );
  XNOR2_X1 U343 ( .A(n468), .B(n467), .ZN(G1350GAT) );
  XNOR2_X1 U344 ( .A(n445), .B(n444), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT73), .B(G92GAT), .Z(n291) );
  XNOR2_X1 U346 ( .A(G134GAT), .B(G106GAT), .ZN(n290) );
  XNOR2_X1 U347 ( .A(n291), .B(n290), .ZN(n307) );
  XOR2_X1 U348 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n293) );
  NAND2_X1 U349 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U350 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U351 ( .A(n294), .B(KEYINPUT64), .Z(n299) );
  XNOR2_X1 U352 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n296), .B(n295), .ZN(n430) );
  XNOR2_X1 U354 ( .A(G36GAT), .B(G190GAT), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n297), .B(G218GAT), .ZN(n367) );
  XNOR2_X1 U356 ( .A(n430), .B(n367), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U358 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n301) );
  XNOR2_X1 U359 ( .A(KEYINPUT74), .B(KEYINPUT11), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U361 ( .A(n303), .B(n302), .Z(n305) );
  XOR2_X1 U362 ( .A(G50GAT), .B(G162GAT), .Z(n360) );
  XOR2_X1 U363 ( .A(G99GAT), .B(G85GAT), .Z(n418) );
  XNOR2_X1 U364 ( .A(n360), .B(n418), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U366 ( .A(KEYINPUT36), .B(n555), .ZN(n575) );
  XOR2_X1 U367 ( .A(KEYINPUT76), .B(KEYINPUT15), .Z(n309) );
  NAND2_X1 U368 ( .A1(G231GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U370 ( .A(n310), .B(KEYINPUT12), .Z(n318) );
  XOR2_X1 U371 ( .A(G155GAT), .B(G211GAT), .Z(n312) );
  XNOR2_X1 U372 ( .A(G22GAT), .B(G127GAT), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U374 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n314) );
  XNOR2_X1 U375 ( .A(G78GAT), .B(G64GAT), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U379 ( .A(G8GAT), .B(G183GAT), .Z(n377) );
  XOR2_X1 U380 ( .A(n319), .B(n377), .Z(n322) );
  XOR2_X1 U381 ( .A(G15GAT), .B(G1GAT), .Z(n437) );
  XNOR2_X1 U382 ( .A(G71GAT), .B(G57GAT), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n320), .B(KEYINPUT13), .ZN(n424) );
  XNOR2_X1 U384 ( .A(n437), .B(n424), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n572) );
  XOR2_X1 U386 ( .A(KEYINPUT84), .B(G71GAT), .Z(n324) );
  XNOR2_X1 U387 ( .A(KEYINPUT82), .B(KEYINPUT20), .ZN(n323) );
  XNOR2_X1 U388 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U389 ( .A(G183GAT), .B(KEYINPUT83), .Z(n326) );
  XNOR2_X1 U390 ( .A(KEYINPUT65), .B(KEYINPUT86), .ZN(n325) );
  XNOR2_X1 U391 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U392 ( .A(n328), .B(n327), .Z(n334) );
  XOR2_X1 U393 ( .A(G99GAT), .B(KEYINPUT85), .Z(n331) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n287), .B(n329), .ZN(n373) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(n373), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U398 ( .A(G190GAT), .B(n332), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U400 ( .A(KEYINPUT81), .B(G176GAT), .Z(n336) );
  NAND2_X1 U401 ( .A1(G227GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U402 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U403 ( .A(n338), .B(n337), .Z(n346) );
  XOR2_X1 U404 ( .A(G120GAT), .B(G127GAT), .Z(n340) );
  XNOR2_X1 U405 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n339) );
  XNOR2_X1 U406 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U407 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n342) );
  XNOR2_X1 U408 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U410 ( .A(n344), .B(n343), .Z(n396) );
  XNOR2_X1 U411 ( .A(G15GAT), .B(n396), .ZN(n345) );
  XOR2_X1 U412 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n348) );
  XNOR2_X1 U413 ( .A(G218GAT), .B(G204GAT), .ZN(n347) );
  XNOR2_X1 U414 ( .A(n348), .B(n347), .ZN(n364) );
  XOR2_X1 U415 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n350) );
  NAND2_X1 U416 ( .A1(G228GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U418 ( .A(n351), .B(KEYINPUT24), .Z(n356) );
  XNOR2_X1 U419 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n352), .B(G211GAT), .ZN(n372) );
  XOR2_X1 U421 ( .A(G155GAT), .B(KEYINPUT2), .Z(n354) );
  XNOR2_X1 U422 ( .A(KEYINPUT88), .B(KEYINPUT3), .ZN(n353) );
  XNOR2_X1 U423 ( .A(n354), .B(n353), .ZN(n392) );
  XNOR2_X1 U424 ( .A(n372), .B(n392), .ZN(n355) );
  XNOR2_X1 U425 ( .A(n356), .B(n355), .ZN(n359) );
  XOR2_X1 U426 ( .A(G78GAT), .B(G148GAT), .Z(n358) );
  XNOR2_X1 U427 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n412) );
  XOR2_X1 U429 ( .A(n359), .B(n412), .Z(n362) );
  XOR2_X1 U430 ( .A(G141GAT), .B(G22GAT), .Z(n438) );
  XNOR2_X1 U431 ( .A(n438), .B(n360), .ZN(n361) );
  XNOR2_X1 U432 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U433 ( .A(n364), .B(n363), .ZN(n463) );
  XOR2_X1 U434 ( .A(KEYINPUT26), .B(n365), .Z(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(KEYINPUT93), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n368), .B(KEYINPUT92), .ZN(n371) );
  XOR2_X1 U437 ( .A(G64GAT), .B(G92GAT), .Z(n370) );
  XNOR2_X1 U438 ( .A(G176GAT), .B(G204GAT), .ZN(n369) );
  XNOR2_X1 U439 ( .A(n370), .B(n369), .ZN(n425) );
  XOR2_X1 U440 ( .A(n371), .B(n425), .Z(n375) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U443 ( .A(n377), .B(n376), .Z(n379) );
  NAND2_X1 U444 ( .A1(G226GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n509) );
  XNOR2_X1 U446 ( .A(n509), .B(KEYINPUT27), .ZN(n402) );
  NAND2_X1 U447 ( .A1(n559), .A2(n402), .ZN(n383) );
  NAND2_X1 U448 ( .A1(n518), .A2(n509), .ZN(n380) );
  NAND2_X1 U449 ( .A1(n463), .A2(n380), .ZN(n381) );
  XOR2_X1 U450 ( .A(KEYINPUT25), .B(n381), .Z(n382) );
  NAND2_X1 U451 ( .A1(n383), .A2(n382), .ZN(n401) );
  XOR2_X1 U452 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n385) );
  XNOR2_X1 U453 ( .A(KEYINPUT4), .B(G57GAT), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n385), .B(n384), .ZN(n400) );
  XOR2_X1 U455 ( .A(G85GAT), .B(G162GAT), .Z(n387) );
  XNOR2_X1 U456 ( .A(G141GAT), .B(G29GAT), .ZN(n386) );
  XNOR2_X1 U457 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U458 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n389) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(G148GAT), .ZN(n388) );
  XNOR2_X1 U460 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U461 ( .A(n391), .B(n390), .Z(n398) );
  XOR2_X1 U462 ( .A(n392), .B(KEYINPUT6), .Z(n394) );
  NAND2_X1 U463 ( .A1(G225GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U465 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U467 ( .A(n400), .B(n399), .Z(n507) );
  INV_X1 U468 ( .A(n507), .ZN(n462) );
  NAND2_X1 U469 ( .A1(n401), .A2(n462), .ZN(n407) );
  NAND2_X1 U470 ( .A1(n507), .A2(n402), .ZN(n534) );
  XNOR2_X1 U471 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n403), .B(n463), .ZN(n514) );
  XNOR2_X1 U473 ( .A(n517), .B(KEYINPUT94), .ZN(n405) );
  INV_X1 U474 ( .A(n518), .ZN(n404) );
  NAND2_X1 U475 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X1 U476 ( .A1(n407), .A2(n406), .ZN(n471) );
  NAND2_X1 U477 ( .A1(n572), .A2(n471), .ZN(n408) );
  NOR2_X1 U478 ( .A1(n575), .A2(n408), .ZN(n409) );
  XNOR2_X1 U479 ( .A(KEYINPUT37), .B(n409), .ZN(n505) );
  AND2_X1 U480 ( .A1(G230GAT), .A2(G233GAT), .ZN(n410) );
  INV_X1 U481 ( .A(KEYINPUT70), .ZN(n413) );
  NAND2_X1 U482 ( .A1(n414), .A2(n413), .ZN(n417) );
  INV_X1 U483 ( .A(n414), .ZN(n415) );
  NAND2_X1 U484 ( .A1(n415), .A2(KEYINPUT70), .ZN(n416) );
  NAND2_X1 U485 ( .A1(n417), .A2(n416), .ZN(n423) );
  XNOR2_X1 U486 ( .A(G120GAT), .B(n418), .ZN(n421) );
  XOR2_X1 U487 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n420) );
  XNOR2_X1 U488 ( .A(KEYINPUT31), .B(KEYINPUT69), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n567) );
  XOR2_X1 U491 ( .A(G113GAT), .B(G36GAT), .Z(n429) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(G50GAT), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n442) );
  XOR2_X1 U494 ( .A(n430), .B(KEYINPUT29), .Z(n432) );
  NAND2_X1 U495 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U496 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U497 ( .A(G8GAT), .B(KEYINPUT30), .Z(n434) );
  XNOR2_X1 U498 ( .A(G197GAT), .B(KEYINPUT68), .ZN(n433) );
  XNOR2_X1 U499 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U500 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U503 ( .A(n442), .B(n441), .Z(n561) );
  NAND2_X1 U504 ( .A1(n567), .A2(n493), .ZN(n473) );
  NOR2_X1 U505 ( .A1(n505), .A2(n473), .ZN(n443) );
  XNOR2_X1 U506 ( .A(KEYINPUT38), .B(n289), .ZN(n491) );
  NAND2_X1 U507 ( .A1(n491), .A2(n518), .ZN(n445) );
  XNOR2_X1 U508 ( .A(KEYINPUT45), .B(KEYINPUT110), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U510 ( .A(KEYINPUT111), .B(n449), .ZN(n450) );
  NOR2_X1 U511 ( .A1(n493), .A2(n450), .ZN(n457) );
  NAND2_X1 U512 ( .A1(n555), .A2(n572), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n567), .B(KEYINPUT41), .ZN(n539) );
  NAND2_X1 U514 ( .A1(n539), .A2(n493), .ZN(n452) );
  NOR2_X1 U515 ( .A1(n454), .A2(n453), .ZN(n455) );
  XOR2_X1 U516 ( .A(KEYINPUT47), .B(n455), .Z(n456) );
  NOR2_X1 U517 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n509), .B(KEYINPUT121), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n460), .B(KEYINPUT54), .ZN(n461) );
  NAND2_X1 U520 ( .A1(n560), .A2(n463), .ZN(n464) );
  XNOR2_X1 U521 ( .A(KEYINPUT55), .B(n464), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n465), .A2(n518), .ZN(n554) );
  NOR2_X1 U523 ( .A1(n572), .A2(n554), .ZN(n468) );
  INV_X1 U524 ( .A(n572), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n555), .A2(n469), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(n470), .Z(n472) );
  NAND2_X1 U527 ( .A1(n472), .A2(n471), .ZN(n494) );
  NOR2_X1 U528 ( .A1(n473), .A2(n494), .ZN(n481) );
  NAND2_X1 U529 ( .A1(n481), .A2(n507), .ZN(n477) );
  XOR2_X1 U530 ( .A(KEYINPUT97), .B(KEYINPUT34), .Z(n475) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n477), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n481), .A2(n509), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U537 ( .A1(n481), .A2(n518), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n483) );
  NAND2_X1 U540 ( .A1(n481), .A2(n514), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n484), .ZN(G1327GAT) );
  NAND2_X1 U543 ( .A1(n491), .A2(n507), .ZN(n488) );
  XOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n486) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT100), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  XOR2_X1 U548 ( .A(G36GAT), .B(KEYINPUT103), .Z(n490) );
  NAND2_X1 U549 ( .A1(n509), .A2(n491), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1329GAT) );
  NAND2_X1 U551 ( .A1(n491), .A2(n514), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n496) );
  XNOR2_X1 U554 ( .A(KEYINPUT105), .B(n539), .ZN(n550) );
  OR2_X1 U555 ( .A1(n493), .A2(n550), .ZN(n506) );
  NOR2_X1 U556 ( .A1(n506), .A2(n494), .ZN(n501) );
  NAND2_X1 U557 ( .A1(n501), .A2(n507), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U559 ( .A(G57GAT), .B(n497), .Z(G1332GAT) );
  NAND2_X1 U560 ( .A1(n501), .A2(n509), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U562 ( .A1(n501), .A2(n518), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT106), .ZN(n500) );
  XNOR2_X1 U564 ( .A(G71GAT), .B(n500), .ZN(G1334GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U566 ( .A1(n501), .A2(n514), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U568 ( .A(G78GAT), .B(n504), .Z(G1335GAT) );
  NOR2_X1 U569 ( .A1(n505), .A2(n506), .ZN(n513) );
  NAND2_X1 U570 ( .A1(n513), .A2(n507), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n508), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U572 ( .A1(n513), .A2(n509), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n510), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U574 ( .A1(n513), .A2(n518), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(KEYINPUT108), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G99GAT), .B(n512), .ZN(G1338GAT) );
  NAND2_X1 U577 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n515), .B(KEYINPUT44), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G106GAT), .B(n516), .ZN(G1339GAT) );
  XOR2_X1 U580 ( .A(G113GAT), .B(KEYINPUT113), .Z(n522) );
  NAND2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U582 ( .A1(n535), .A2(n519), .ZN(n520) );
  XOR2_X1 U583 ( .A(KEYINPUT112), .B(n520), .Z(n530) );
  OR2_X1 U584 ( .A1(n530), .A2(n561), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(G1340GAT) );
  XNOR2_X1 U586 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n524) );
  NOR2_X1 U587 ( .A1(n550), .A2(n530), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1341GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n526) );
  XNOR2_X1 U590 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n572), .A2(n530), .ZN(n527) );
  XOR2_X1 U593 ( .A(n528), .B(n527), .Z(n529) );
  XNOR2_X1 U594 ( .A(KEYINPUT114), .B(n529), .ZN(G1342GAT) );
  XNOR2_X1 U595 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n532) );
  NOR2_X1 U596 ( .A1(n555), .A2(n530), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U598 ( .A(G134GAT), .B(n533), .Z(G1343GAT) );
  NOR2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U600 ( .A1(n536), .A2(n559), .ZN(n546) );
  NOR2_X1 U601 ( .A1(n561), .A2(n546), .ZN(n537) );
  XOR2_X1 U602 ( .A(KEYINPUT118), .B(n537), .Z(n538) );
  XNOR2_X1 U603 ( .A(G141GAT), .B(n538), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n542) );
  INV_X1 U605 ( .A(n546), .ZN(n540) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U609 ( .A1(n572), .A2(n546), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1346GAT) );
  NOR2_X1 U612 ( .A1(n555), .A2(n546), .ZN(n547) );
  XOR2_X1 U613 ( .A(KEYINPUT120), .B(n547), .Z(n548) );
  XNOR2_X1 U614 ( .A(G162GAT), .B(n548), .ZN(G1347GAT) );
  NOR2_X1 U615 ( .A1(n561), .A2(n554), .ZN(n549) );
  XOR2_X1 U616 ( .A(G169GAT), .B(n549), .Z(G1348GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n554), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(n553), .ZN(G1349GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(n558), .ZN(G1351GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n574) );
  NOR2_X1 U626 ( .A1(n561), .A2(n574), .ZN(n566) );
  XOR2_X1 U627 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n563) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(KEYINPUT59), .B(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1352GAT) );
  NOR2_X1 U632 ( .A1(n574), .A2(n567), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n569) );
  XNOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n574), .ZN(n573) );
  XOR2_X1 U638 ( .A(G211GAT), .B(n573), .Z(G1354GAT) );
  NOR2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT62), .B(n576), .Z(n577) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(n577), .ZN(G1355GAT) );
endmodule

