

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748;

  AND2_X2 U378 ( .A1(n403), .A2(n404), .ZN(n402) );
  XNOR2_X2 U379 ( .A(n514), .B(n513), .ZN(n533) );
  XNOR2_X2 U380 ( .A(n507), .B(n418), .ZN(n484) );
  XNOR2_X2 U381 ( .A(n419), .B(G146), .ZN(n507) );
  INV_X2 U382 ( .A(n566), .ZN(n539) );
  INV_X1 U383 ( .A(n601), .ZN(n677) );
  INV_X1 U384 ( .A(G119), .ZN(n397) );
  NOR2_X1 U385 ( .A1(n702), .A2(n713), .ZN(n366) );
  AND2_X1 U386 ( .A1(n376), .A2(n375), .ZN(n374) );
  NOR2_X1 U387 ( .A1(n625), .A2(n713), .ZN(n365) );
  NOR2_X2 U388 ( .A1(n746), .A2(n634), .ZN(n593) );
  NOR2_X1 U389 ( .A1(n640), .A2(n630), .ZN(n605) );
  OR2_X1 U390 ( .A1(n543), .A2(n559), .ZN(n544) );
  OR2_X1 U391 ( .A1(n604), .A2(n369), .ZN(n368) );
  XNOR2_X2 U392 ( .A(KEYINPUT38), .B(n539), .ZN(n666) );
  AND2_X1 U393 ( .A1(n523), .A2(n367), .ZN(n540) );
  XNOR2_X1 U394 ( .A(n370), .B(KEYINPUT19), .ZN(n572) );
  BUF_X1 U395 ( .A(n533), .Z(n566) );
  XNOR2_X1 U396 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U397 ( .A(n531), .B(KEYINPUT1), .ZN(n670) );
  XNOR2_X1 U398 ( .A(n455), .B(G472), .ZN(n601) );
  XNOR2_X1 U399 ( .A(n444), .B(n360), .ZN(n506) );
  XNOR2_X1 U400 ( .A(n398), .B(n397), .ZN(n396) );
  XNOR2_X1 U401 ( .A(n433), .B(G107), .ZN(n714) );
  INV_X2 U402 ( .A(G953), .ZN(n379) );
  NAND2_X1 U403 ( .A1(n719), .A2(n401), .ZN(n400) );
  NOR2_X2 U404 ( .A1(n743), .A2(n747), .ZN(n556) );
  NOR2_X1 U405 ( .A1(n531), .A2(n671), .ZN(n602) );
  NOR2_X2 U406 ( .A1(n719), .A2(KEYINPUT2), .ZN(n652) );
  XOR2_X1 U407 ( .A(n434), .B(n729), .Z(n444) );
  XNOR2_X1 U408 ( .A(KEYINPUT69), .B(G101), .ZN(n434) );
  XNOR2_X1 U409 ( .A(KEYINPUT10), .B(KEYINPUT72), .ZN(n418) );
  XNOR2_X1 U410 ( .A(G902), .B(KEYINPUT15), .ZN(n610) );
  XNOR2_X1 U411 ( .A(n505), .B(n502), .ZN(n385) );
  NOR2_X1 U412 ( .A1(n570), .A2(n422), .ZN(n571) );
  AND2_X1 U413 ( .A1(G898), .A2(G953), .ZN(n422) );
  NOR2_X1 U414 ( .A1(G953), .A2(G237), .ZN(n485) );
  INV_X1 U415 ( .A(n660), .ZN(n389) );
  XNOR2_X1 U416 ( .A(n745), .B(KEYINPUT70), .ZN(n592) );
  XNOR2_X1 U417 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n501) );
  XNOR2_X1 U418 ( .A(n504), .B(n421), .ZN(n505) );
  XNOR2_X1 U419 ( .A(G122), .B(G113), .ZN(n488) );
  XOR2_X1 U420 ( .A(G104), .B(G143), .Z(n487) );
  INV_X1 U421 ( .A(KEYINPUT87), .ZN(n392) );
  XNOR2_X1 U422 ( .A(n505), .B(n503), .ZN(n383) );
  INV_X1 U423 ( .A(G125), .ZN(n419) );
  INV_X1 U424 ( .A(n714), .ZN(n360) );
  AND2_X1 U425 ( .A1(n719), .A2(n738), .ZN(n650) );
  NAND2_X1 U426 ( .A1(n417), .A2(n416), .ZN(n529) );
  AND2_X1 U427 ( .A1(n673), .A2(n354), .ZN(n416) );
  XNOR2_X1 U428 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U429 ( .A(n495), .B(n494), .ZN(n547) );
  INV_X1 U430 ( .A(G122), .ZN(n498) );
  XNOR2_X1 U431 ( .A(n588), .B(n587), .ZN(n663) );
  INV_X1 U432 ( .A(n582), .ZN(n409) );
  XNOR2_X1 U433 ( .A(n364), .B(G478), .ZN(n546) );
  NOR2_X1 U434 ( .A1(n711), .A2(G902), .ZN(n364) );
  INV_X1 U435 ( .A(n597), .ZN(n407) );
  NAND2_X1 U436 ( .A1(n693), .A2(KEYINPUT121), .ZN(n375) );
  NAND2_X1 U437 ( .A1(n373), .A2(n357), .ZN(n371) );
  INV_X1 U438 ( .A(KEYINPUT121), .ZN(n372) );
  XOR2_X1 U439 ( .A(G128), .B(G143), .Z(n504) );
  XOR2_X1 U440 ( .A(G140), .B(G131), .Z(n482) );
  OR2_X1 U441 ( .A1(G902), .A2(G237), .ZN(n510) );
  NOR2_X1 U442 ( .A1(n355), .A2(n558), .ZN(n413) );
  INV_X1 U443 ( .A(KEYINPUT48), .ZN(n411) );
  XNOR2_X1 U444 ( .A(KEYINPUT95), .B(n436), .ZN(n728) );
  XNOR2_X1 U445 ( .A(n504), .B(G134), .ZN(n471) );
  XNOR2_X1 U446 ( .A(n471), .B(G146), .ZN(n443) );
  NOR2_X1 U447 ( .A1(n671), .A2(n670), .ZN(n598) );
  XNOR2_X1 U448 ( .A(G110), .B(G104), .ZN(n433) );
  XOR2_X1 U449 ( .A(KEYINPUT80), .B(KEYINPUT24), .Z(n429) );
  XNOR2_X1 U450 ( .A(G110), .B(G119), .ZN(n428) );
  XNOR2_X1 U451 ( .A(G140), .B(G128), .ZN(n423) );
  XNOR2_X1 U452 ( .A(G107), .B(G122), .ZN(n472) );
  XNOR2_X1 U453 ( .A(KEYINPUT105), .B(KEYINPUT7), .ZN(n475) );
  XNOR2_X1 U454 ( .A(n727), .B(n492), .ZN(n616) );
  XNOR2_X1 U455 ( .A(n491), .B(n490), .ZN(n492) );
  INV_X1 U456 ( .A(n610), .ZN(n404) );
  XNOR2_X1 U457 ( .A(KEYINPUT45), .B(KEYINPUT65), .ZN(n608) );
  XNOR2_X1 U458 ( .A(n508), .B(n509), .ZN(n695) );
  XNOR2_X1 U459 ( .A(n506), .B(n507), .ZN(n508) );
  NAND2_X1 U460 ( .A1(n383), .A2(n716), .ZN(n382) );
  AND2_X1 U461 ( .A1(n602), .A2(n354), .ZN(n367) );
  NOR2_X1 U462 ( .A1(n521), .A2(n601), .ZN(n522) );
  NAND2_X1 U463 ( .A1(n533), .A2(n665), .ZN(n370) );
  INV_X1 U464 ( .A(KEYINPUT28), .ZN(n414) );
  NOR2_X1 U465 ( .A1(G952), .A2(n379), .ZN(n713) );
  NOR2_X1 U466 ( .A1(n663), .A2(n604), .ZN(n362) );
  XNOR2_X1 U467 ( .A(n578), .B(KEYINPUT66), .ZN(n579) );
  INV_X1 U468 ( .A(KEYINPUT32), .ZN(n578) );
  XNOR2_X1 U469 ( .A(n363), .B(KEYINPUT67), .ZN(n583) );
  NOR2_X1 U470 ( .A1(n581), .A2(n408), .ZN(n363) );
  NAND2_X1 U471 ( .A1(n409), .A2(n601), .ZN(n408) );
  NAND2_X1 U472 ( .A1(n405), .A2(n358), .ZN(n387) );
  NOR2_X1 U473 ( .A1(n582), .A2(n407), .ZN(n406) );
  INV_X1 U474 ( .A(KEYINPUT53), .ZN(n377) );
  AND2_X1 U475 ( .A1(n569), .A2(n465), .ZN(n354) );
  AND2_X1 U476 ( .A1(n538), .A2(n537), .ZN(n355) );
  AND2_X1 U477 ( .A1(n744), .A2(n567), .ZN(n356) );
  AND2_X1 U478 ( .A1(n381), .A2(n372), .ZN(n357) );
  AND2_X1 U479 ( .A1(n406), .A2(n674), .ZN(n358) );
  XNOR2_X1 U480 ( .A(n548), .B(KEYINPUT107), .ZN(n662) );
  XNOR2_X1 U481 ( .A(n393), .B(n392), .ZN(n607) );
  NAND2_X1 U482 ( .A1(n359), .A2(n382), .ZN(n509) );
  NAND2_X1 U483 ( .A1(n384), .A2(n385), .ZN(n359) );
  NOR2_X1 U484 ( .A1(G902), .A2(n622), .ZN(n455) );
  XNOR2_X1 U485 ( .A(n362), .B(KEYINPUT34), .ZN(n590) );
  NAND2_X1 U486 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U487 ( .A1(n695), .A2(n610), .ZN(n514) );
  XNOR2_X1 U488 ( .A(n443), .B(n444), .ZN(n454) );
  NOR2_X2 U489 ( .A1(n361), .A2(n607), .ZN(n609) );
  NAND2_X1 U490 ( .A1(n595), .A2(n596), .ZN(n361) );
  XNOR2_X2 U491 ( .A(n591), .B(KEYINPUT35), .ZN(n745) );
  XOR2_X2 U492 ( .A(G137), .B(KEYINPUT73), .Z(n435) );
  AND2_X2 U493 ( .A1(n410), .A2(n356), .ZN(n738) );
  XNOR2_X1 U494 ( .A(n365), .B(n626), .ZN(G57) );
  XNOR2_X1 U495 ( .A(n366), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X2 U496 ( .A(n368), .B(KEYINPUT22), .ZN(n581) );
  NAND2_X1 U497 ( .A1(n662), .A2(n673), .ZN(n369) );
  XNOR2_X2 U498 ( .A(n573), .B(KEYINPUT0), .ZN(n604) );
  INV_X1 U499 ( .A(n572), .ZN(n568) );
  NAND2_X1 U500 ( .A1(n374), .A2(n371), .ZN(n380) );
  INV_X1 U501 ( .A(n694), .ZN(n373) );
  NAND2_X1 U502 ( .A1(n694), .A2(KEYINPUT121), .ZN(n376) );
  XNOR2_X1 U503 ( .A(n378), .B(n377), .ZN(G75) );
  NAND2_X1 U504 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U505 ( .A(n693), .ZN(n381) );
  INV_X1 U506 ( .A(n716), .ZN(n384) );
  INV_X1 U507 ( .A(n387), .ZN(n627) );
  XNOR2_X1 U508 ( .A(n386), .B(n395), .ZN(n394) );
  NAND2_X1 U509 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U510 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U511 ( .A(n605), .B(n391), .ZN(n390) );
  INV_X1 U512 ( .A(KEYINPUT100), .ZN(n391) );
  XNOR2_X2 U513 ( .A(n545), .B(n544), .ZN(n743) );
  XNOR2_X1 U514 ( .A(n412), .B(n411), .ZN(n410) );
  XNOR2_X2 U515 ( .A(KEYINPUT4), .B(KEYINPUT71), .ZN(n729) );
  NOR2_X2 U516 ( .A1(n619), .A2(n713), .ZN(n621) );
  NAND2_X1 U517 ( .A1(n557), .A2(n413), .ZN(n412) );
  NAND2_X1 U518 ( .A1(n394), .A2(n606), .ZN(n393) );
  INV_X1 U519 ( .A(KEYINPUT108), .ZN(n395) );
  XNOR2_X2 U520 ( .A(n500), .B(n499), .ZN(n716) );
  XNOR2_X2 U521 ( .A(n396), .B(n451), .ZN(n500) );
  XNOR2_X2 U522 ( .A(KEYINPUT75), .B(KEYINPUT3), .ZN(n398) );
  NOR2_X4 U523 ( .A1(n399), .A2(n652), .ZN(n709) );
  NAND2_X2 U524 ( .A1(n402), .A2(n400), .ZN(n399) );
  AND2_X1 U525 ( .A1(n738), .A2(KEYINPUT2), .ZN(n401) );
  OR2_X1 U526 ( .A1(n738), .A2(KEYINPUT2), .ZN(n403) );
  XNOR2_X2 U527 ( .A(n609), .B(n608), .ZN(n719) );
  INV_X1 U528 ( .A(n581), .ZN(n405) );
  XNOR2_X1 U529 ( .A(n415), .B(n414), .ZN(n530) );
  NOR2_X1 U530 ( .A1(n529), .A2(n601), .ZN(n415) );
  INV_X1 U531 ( .A(n575), .ZN(n417) );
  XNOR2_X1 U532 ( .A(n484), .B(n424), .ZN(n425) );
  BUF_X1 U533 ( .A(n575), .Z(n674) );
  XNOR2_X1 U534 ( .A(G116), .B(G113), .ZN(n451) );
  XNOR2_X1 U535 ( .A(n470), .B(n469), .ZN(n575) );
  XNOR2_X1 U536 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X2 U537 ( .A(n550), .B(KEYINPUT41), .ZN(n685) );
  XNOR2_X2 U538 ( .A(n442), .B(n441), .ZN(n531) );
  XOR2_X1 U539 ( .A(n429), .B(n428), .Z(n420) );
  AND2_X1 U540 ( .A1(G224), .A2(n379), .ZN(n421) );
  INV_X1 U541 ( .A(n649), .ZN(n567) );
  XNOR2_X1 U542 ( .A(KEYINPUT23), .B(KEYINPUT76), .ZN(n424) );
  XNOR2_X1 U543 ( .A(n452), .B(n500), .ZN(n453) );
  XNOR2_X1 U544 ( .A(n493), .B(G475), .ZN(n494) );
  XNOR2_X1 U545 ( .A(n454), .B(n453), .ZN(n622) );
  XNOR2_X1 U546 ( .A(n498), .B(KEYINPUT16), .ZN(n499) );
  BUF_X1 U547 ( .A(n695), .Z(n699) );
  INV_X1 U548 ( .A(KEYINPUT39), .ZN(n541) );
  XNOR2_X1 U549 ( .A(n622), .B(KEYINPUT62), .ZN(n623) );
  XNOR2_X1 U550 ( .A(n542), .B(n541), .ZN(n559) );
  XNOR2_X1 U551 ( .A(n624), .B(n623), .ZN(n625) );
  INV_X1 U552 ( .A(KEYINPUT123), .ZN(n614) );
  XNOR2_X1 U553 ( .A(n580), .B(n579), .ZN(n746) );
  XNOR2_X1 U554 ( .A(n423), .B(n435), .ZN(n426) );
  XOR2_X1 U555 ( .A(n426), .B(n425), .Z(n432) );
  NAND2_X1 U556 ( .A1(G234), .A2(n379), .ZN(n427) );
  XOR2_X1 U557 ( .A(KEYINPUT8), .B(n427), .Z(n477) );
  NAND2_X1 U558 ( .A1(G221), .A2(n477), .ZN(n430) );
  XNOR2_X1 U559 ( .A(n430), .B(n420), .ZN(n431) );
  XNOR2_X1 U560 ( .A(n432), .B(n431), .ZN(n612) );
  XNOR2_X1 U561 ( .A(KEYINPUT74), .B(G469), .ZN(n442) );
  XNOR2_X1 U562 ( .A(n506), .B(n443), .ZN(n440) );
  INV_X1 U563 ( .A(n435), .ZN(n436) );
  XOR2_X1 U564 ( .A(n728), .B(n482), .Z(n438) );
  NAND2_X1 U565 ( .A1(G227), .A2(n379), .ZN(n437) );
  XNOR2_X1 U566 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U567 ( .A(n439), .B(n440), .ZN(n703) );
  NOR2_X1 U568 ( .A1(G902), .A2(n703), .ZN(n441) );
  XOR2_X1 U569 ( .A(KEYINPUT91), .B(n409), .Z(n574) );
  INV_X1 U570 ( .A(n574), .ZN(n518) );
  XOR2_X1 U571 ( .A(KEYINPUT36), .B(KEYINPUT88), .Z(n516) );
  XOR2_X1 U572 ( .A(KEYINPUT98), .B(KEYINPUT78), .Z(n446) );
  XNOR2_X1 U573 ( .A(G137), .B(G131), .ZN(n445) );
  XNOR2_X1 U574 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U575 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n448) );
  NAND2_X1 U576 ( .A1(n485), .A2(G210), .ZN(n447) );
  XNOR2_X1 U577 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U578 ( .A(n450), .B(n449), .Z(n452) );
  XNOR2_X1 U579 ( .A(KEYINPUT6), .B(KEYINPUT106), .ZN(n456) );
  XOR2_X1 U580 ( .A(n677), .B(n456), .Z(n585) );
  INV_X1 U581 ( .A(n585), .ZN(n597) );
  NAND2_X1 U582 ( .A1(G214), .A2(n510), .ZN(n457) );
  XNOR2_X1 U583 ( .A(KEYINPUT94), .B(n457), .ZN(n665) );
  XOR2_X1 U584 ( .A(KEYINPUT21), .B(KEYINPUT96), .Z(n460) );
  NAND2_X1 U585 ( .A1(G234), .A2(n610), .ZN(n458) );
  XNOR2_X1 U586 ( .A(KEYINPUT20), .B(n458), .ZN(n466) );
  NAND2_X1 U587 ( .A1(n466), .A2(G221), .ZN(n459) );
  XNOR2_X1 U588 ( .A(n460), .B(n459), .ZN(n673) );
  NAND2_X1 U589 ( .A1(G237), .A2(G234), .ZN(n461) );
  XNOR2_X1 U590 ( .A(n461), .B(KEYINPUT14), .ZN(n690) );
  OR2_X1 U591 ( .A1(n379), .A2(G902), .ZN(n462) );
  NAND2_X1 U592 ( .A1(n690), .A2(n462), .ZN(n464) );
  NOR2_X1 U593 ( .A1(G953), .A2(G952), .ZN(n463) );
  NOR2_X1 U594 ( .A1(n464), .A2(n463), .ZN(n569) );
  NAND2_X1 U595 ( .A1(G953), .A2(G900), .ZN(n465) );
  NOR2_X1 U596 ( .A1(G902), .A2(n612), .ZN(n470) );
  XOR2_X1 U597 ( .A(KEYINPUT25), .B(KEYINPUT79), .Z(n468) );
  NAND2_X1 U598 ( .A1(n466), .A2(G217), .ZN(n467) );
  XNOR2_X1 U599 ( .A(n468), .B(n467), .ZN(n469) );
  INV_X1 U600 ( .A(n471), .ZN(n733) );
  XOR2_X1 U601 ( .A(KEYINPUT103), .B(G116), .Z(n473) );
  XNOR2_X1 U602 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U603 ( .A(n733), .B(n474), .ZN(n481) );
  XNOR2_X1 U604 ( .A(n475), .B(KEYINPUT104), .ZN(n476) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n476), .Z(n479) );
  NAND2_X1 U606 ( .A1(G217), .A2(n477), .ZN(n478) );
  XNOR2_X1 U607 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U608 ( .A(n481), .B(n480), .ZN(n711) );
  INV_X1 U609 ( .A(n482), .ZN(n483) );
  XNOR2_X1 U610 ( .A(n484), .B(n483), .ZN(n727) );
  NAND2_X1 U611 ( .A1(n485), .A2(G214), .ZN(n486) );
  XNOR2_X1 U612 ( .A(n487), .B(n486), .ZN(n491) );
  XOR2_X1 U613 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n489) );
  XNOR2_X1 U614 ( .A(n489), .B(n488), .ZN(n490) );
  NOR2_X1 U615 ( .A1(G902), .A2(n616), .ZN(n495) );
  XNOR2_X1 U616 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n493) );
  XOR2_X1 U617 ( .A(n547), .B(KEYINPUT102), .Z(n519) );
  NAND2_X1 U618 ( .A1(n546), .A2(n519), .ZN(n543) );
  NOR2_X1 U619 ( .A1(n529), .A2(n543), .ZN(n496) );
  NAND2_X1 U620 ( .A1(n665), .A2(n496), .ZN(n497) );
  NOR2_X1 U621 ( .A1(n597), .A2(n497), .ZN(n562) );
  XOR2_X1 U622 ( .A(n501), .B(KEYINPUT18), .Z(n503) );
  INV_X1 U623 ( .A(n503), .ZN(n502) );
  XOR2_X1 U624 ( .A(KEYINPUT93), .B(KEYINPUT81), .Z(n512) );
  NAND2_X1 U625 ( .A1(G210), .A2(n510), .ZN(n511) );
  NAND2_X1 U626 ( .A1(n562), .A2(n566), .ZN(n515) );
  XNOR2_X1 U627 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U628 ( .A1(n518), .A2(n517), .ZN(n646) );
  XNOR2_X1 U629 ( .A(n646), .B(KEYINPUT86), .ZN(n528) );
  NOR2_X1 U630 ( .A1(n546), .A2(n519), .ZN(n644) );
  INV_X1 U631 ( .A(n543), .ZN(n641) );
  NOR2_X1 U632 ( .A1(n644), .A2(n641), .ZN(n660) );
  NAND2_X1 U633 ( .A1(KEYINPUT47), .A2(n660), .ZN(n520) );
  XNOR2_X1 U634 ( .A(KEYINPUT83), .B(n520), .ZN(n525) );
  INV_X1 U635 ( .A(n665), .ZN(n521) );
  XNOR2_X1 U636 ( .A(KEYINPUT30), .B(n522), .ZN(n523) );
  NAND2_X1 U637 ( .A1(n673), .A2(n575), .ZN(n671) );
  NOR2_X1 U638 ( .A1(n546), .A2(n547), .ZN(n589) );
  NAND2_X1 U639 ( .A1(n540), .A2(n589), .ZN(n524) );
  NOR2_X1 U640 ( .A1(n539), .A2(n524), .ZN(n637) );
  NOR2_X1 U641 ( .A1(n525), .A2(n637), .ZN(n526) );
  XNOR2_X1 U642 ( .A(n526), .B(KEYINPUT82), .ZN(n527) );
  NAND2_X1 U643 ( .A1(n528), .A2(n527), .ZN(n558) );
  INV_X1 U644 ( .A(n644), .ZN(n560) );
  NAND2_X1 U645 ( .A1(n560), .A2(n543), .ZN(n534) );
  NOR2_X1 U646 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U647 ( .A(KEYINPUT111), .B(n532), .ZN(n551) );
  NOR2_X1 U648 ( .A1(n551), .A2(n568), .ZN(n638) );
  NAND2_X1 U649 ( .A1(n534), .A2(n638), .ZN(n536) );
  INV_X1 U650 ( .A(KEYINPUT47), .ZN(n535) );
  NAND2_X1 U651 ( .A1(n536), .A2(n535), .ZN(n538) );
  NAND2_X1 U652 ( .A1(n638), .A2(KEYINPUT47), .ZN(n537) );
  XOR2_X1 U653 ( .A(KEYINPUT40), .B(KEYINPUT112), .Z(n545) );
  NAND2_X1 U654 ( .A1(n540), .A2(n666), .ZN(n542) );
  NAND2_X1 U655 ( .A1(n666), .A2(n665), .ZN(n659) );
  INV_X1 U656 ( .A(n659), .ZN(n549) );
  NAND2_X1 U657 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U658 ( .A1(n549), .A2(n662), .ZN(n550) );
  INV_X1 U659 ( .A(n551), .ZN(n552) );
  NAND2_X1 U660 ( .A1(n685), .A2(n552), .ZN(n553) );
  XOR2_X1 U661 ( .A(KEYINPUT42), .B(n553), .Z(n747) );
  XOR2_X1 U662 ( .A(KEYINPUT46), .B(KEYINPUT85), .Z(n554) );
  XNOR2_X1 U663 ( .A(KEYINPUT64), .B(n554), .ZN(n555) );
  XNOR2_X1 U664 ( .A(n556), .B(n555), .ZN(n557) );
  NOR2_X1 U665 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U666 ( .A(n561), .B(KEYINPUT113), .ZN(n744) );
  XOR2_X1 U667 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n564) );
  NAND2_X1 U668 ( .A1(n562), .A2(n670), .ZN(n563) );
  XNOR2_X1 U669 ( .A(n564), .B(n563), .ZN(n565) );
  NOR2_X1 U670 ( .A1(n566), .A2(n565), .ZN(n649) );
  INV_X1 U671 ( .A(n569), .ZN(n570) );
  NAND2_X1 U672 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U673 ( .A1(n581), .A2(n574), .ZN(n577) );
  NOR2_X1 U674 ( .A1(n674), .A2(n407), .ZN(n576) );
  NAND2_X1 U675 ( .A1(n577), .A2(n576), .ZN(n580) );
  INV_X1 U676 ( .A(n670), .ZN(n582) );
  NOR2_X1 U677 ( .A1(n674), .A2(n583), .ZN(n634) );
  NAND2_X1 U678 ( .A1(KEYINPUT70), .A2(n593), .ZN(n584) );
  NAND2_X1 U679 ( .A1(n584), .A2(KEYINPUT44), .ZN(n596) );
  NAND2_X1 U680 ( .A1(n585), .A2(n598), .ZN(n588) );
  XOR2_X1 U681 ( .A(KEYINPUT33), .B(KEYINPUT77), .Z(n586) );
  XNOR2_X1 U682 ( .A(KEYINPUT109), .B(n586), .ZN(n587) );
  NOR2_X1 U683 ( .A1(KEYINPUT44), .A2(n592), .ZN(n594) );
  NAND2_X1 U684 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U685 ( .A1(n677), .A2(n598), .ZN(n681) );
  NOR2_X1 U686 ( .A1(n604), .A2(n681), .ZN(n600) );
  XNOR2_X1 U687 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n599) );
  XNOR2_X1 U688 ( .A(n600), .B(n599), .ZN(n640) );
  NAND2_X1 U689 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U690 ( .A1(n604), .A2(n603), .ZN(n630) );
  NAND2_X1 U691 ( .A1(n745), .A2(KEYINPUT44), .ZN(n606) );
  NAND2_X1 U692 ( .A1(G217), .A2(n709), .ZN(n611) );
  XNOR2_X1 U693 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X2 U694 ( .A1(n613), .A2(n713), .ZN(n615) );
  XNOR2_X1 U695 ( .A(n615), .B(n614), .ZN(G66) );
  XOR2_X1 U696 ( .A(n616), .B(KEYINPUT59), .Z(n618) );
  NAND2_X1 U697 ( .A1(n709), .A2(G475), .ZN(n617) );
  XNOR2_X1 U698 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U699 ( .A(KEYINPUT60), .B(KEYINPUT68), .ZN(n620) );
  XNOR2_X1 U700 ( .A(n621), .B(n620), .ZN(G60) );
  NAND2_X1 U701 ( .A1(n709), .A2(G472), .ZN(n624) );
  XOR2_X1 U702 ( .A(KEYINPUT63), .B(KEYINPUT114), .Z(n626) );
  XNOR2_X1 U703 ( .A(n627), .B(G101), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT115), .ZN(G3) );
  NAND2_X1 U705 ( .A1(n630), .A2(n641), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n629), .B(G104), .ZN(G6) );
  XOR2_X1 U707 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n632) );
  NAND2_X1 U708 ( .A1(n630), .A2(n644), .ZN(n631) );
  XNOR2_X1 U709 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U710 ( .A(G107), .B(n633), .ZN(G9) );
  XOR2_X1 U711 ( .A(G110), .B(n634), .Z(G12) );
  XOR2_X1 U712 ( .A(G128), .B(KEYINPUT29), .Z(n636) );
  NAND2_X1 U713 ( .A1(n638), .A2(n644), .ZN(n635) );
  XNOR2_X1 U714 ( .A(n636), .B(n635), .ZN(G30) );
  XOR2_X1 U715 ( .A(G143), .B(n637), .Z(G45) );
  NAND2_X1 U716 ( .A1(n638), .A2(n641), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n639), .B(G146), .ZN(G48) );
  NAND2_X1 U718 ( .A1(n640), .A2(n641), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n642), .B(KEYINPUT116), .ZN(n643) );
  XNOR2_X1 U720 ( .A(G113), .B(n643), .ZN(G15) );
  NAND2_X1 U721 ( .A1(n640), .A2(n644), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n645), .B(G116), .ZN(G18) );
  XNOR2_X1 U723 ( .A(KEYINPUT117), .B(KEYINPUT37), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U725 ( .A(G125), .B(n648), .ZN(G27) );
  XOR2_X1 U726 ( .A(G140), .B(n649), .Z(G42) );
  NAND2_X1 U727 ( .A1(KEYINPUT2), .A2(n650), .ZN(n655) );
  NOR2_X1 U728 ( .A1(n738), .A2(KEYINPUT2), .ZN(n651) );
  XNOR2_X1 U729 ( .A(n651), .B(KEYINPUT84), .ZN(n653) );
  NOR2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n658) );
  INV_X1 U732 ( .A(n663), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n685), .A2(n656), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n694) );
  NOR2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(n664) );
  NOR2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n668) );
  OR2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n669), .B(KEYINPUT120), .ZN(n688) );
  NAND2_X1 U741 ( .A1(n671), .A2(n409), .ZN(n672) );
  XNOR2_X1 U742 ( .A(KEYINPUT50), .B(n672), .ZN(n679) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U744 ( .A(KEYINPUT49), .B(n675), .Z(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n680), .B(KEYINPUT118), .ZN(n682) );
  NAND2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U749 ( .A(n683), .B(KEYINPUT119), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n684), .B(KEYINPUT51), .ZN(n686) );
  NAND2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U753 ( .A(KEYINPUT52), .B(n689), .Z(n692) );
  NAND2_X1 U754 ( .A1(n690), .A2(G952), .ZN(n691) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U756 ( .A1(n709), .A2(G210), .ZN(n701) );
  XOR2_X1 U757 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n697) );
  XNOR2_X1 U758 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n696) );
  XNOR2_X1 U759 ( .A(n697), .B(n696), .ZN(n698) );
  XOR2_X1 U760 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n705) );
  XNOR2_X1 U761 ( .A(n703), .B(KEYINPUT122), .ZN(n704) );
  XNOR2_X1 U762 ( .A(n705), .B(n704), .ZN(n707) );
  NAND2_X1 U763 ( .A1(n709), .A2(G469), .ZN(n706) );
  XNOR2_X1 U764 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U765 ( .A1(n713), .A2(n708), .ZN(G54) );
  NAND2_X1 U766 ( .A1(G478), .A2(n709), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U768 ( .A1(n713), .A2(n712), .ZN(G63) );
  XOR2_X1 U769 ( .A(n714), .B(G101), .Z(n715) );
  XNOR2_X1 U770 ( .A(n716), .B(n715), .ZN(n718) );
  NOR2_X1 U771 ( .A1(G898), .A2(n379), .ZN(n717) );
  NOR2_X1 U772 ( .A1(n718), .A2(n717), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n719), .A2(n379), .ZN(n720) );
  XNOR2_X1 U774 ( .A(n720), .B(KEYINPUT124), .ZN(n724) );
  NAND2_X1 U775 ( .A1(G953), .A2(G224), .ZN(n721) );
  XNOR2_X1 U776 ( .A(KEYINPUT61), .B(n721), .ZN(n722) );
  NAND2_X1 U777 ( .A1(n722), .A2(G898), .ZN(n723) );
  NAND2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(G69) );
  XNOR2_X1 U780 ( .A(n727), .B(KEYINPUT125), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n728), .B(n729), .ZN(n730) );
  XNOR2_X1 U782 ( .A(n731), .B(n730), .ZN(n732) );
  XOR2_X1 U783 ( .A(n733), .B(n732), .Z(n739) );
  INV_X1 U784 ( .A(n739), .ZN(n734) );
  XNOR2_X1 U785 ( .A(G227), .B(n734), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n735), .A2(G900), .ZN(n736) );
  NAND2_X1 U787 ( .A1(G953), .A2(n736), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n737), .B(KEYINPUT126), .ZN(n742) );
  XNOR2_X1 U789 ( .A(n739), .B(n738), .ZN(n740) );
  NAND2_X1 U790 ( .A1(n740), .A2(n379), .ZN(n741) );
  NAND2_X1 U791 ( .A1(n742), .A2(n741), .ZN(G72) );
  XOR2_X1 U792 ( .A(G131), .B(n743), .Z(G33) );
  XNOR2_X1 U793 ( .A(G134), .B(n744), .ZN(G36) );
  XOR2_X1 U794 ( .A(G122), .B(n745), .Z(G24) );
  XOR2_X1 U795 ( .A(n746), .B(G119), .Z(G21) );
  XNOR2_X1 U796 ( .A(G137), .B(KEYINPUT127), .ZN(n748) );
  XNOR2_X1 U797 ( .A(n748), .B(n747), .ZN(G39) );
endmodule

