//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G15gat), .ZN(new_n204));
  INV_X1    g003(.A(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G15gat), .A2(G22gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(new_n209), .A3(new_n207), .ZN(new_n212));
  XOR2_X1   g011(.A(KEYINPUT89), .B(G8gat), .Z(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n215), .A2(G71gat), .A3(G78gat), .ZN(new_n216));
  INV_X1    g015(.A(G71gat), .ZN(new_n217));
  INV_X1    g016(.A(G78gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G57gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G64gat), .ZN(new_n221));
  INV_X1    g020(.A(G64gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G57gat), .ZN(new_n223));
  OAI22_X1  g022(.A1(new_n216), .A2(new_n219), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT9), .B1(new_n221), .B2(new_n223), .ZN(new_n225));
  XNOR2_X1  g024(.A(G71gat), .B(G78gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT93), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(G57gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n220), .A2(G64gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n215), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT93), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n231), .A2(new_n232), .A3(new_n226), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n224), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT21), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n212), .A2(KEYINPUT87), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n206), .A2(new_n237), .A3(new_n209), .A4(new_n207), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n211), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(KEYINPUT88), .A3(G8gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT88), .B1(new_n239), .B2(G8gat), .ZN(new_n242));
  OAI221_X1 g041(.A(new_n214), .B1(new_n234), .B2(new_n235), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G183gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n234), .A2(new_n235), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n246), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n247), .A2(G231gat), .A3(G233gat), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G231gat), .A2(G233gat), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n245), .A2(new_n246), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n245), .A2(new_n246), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G127gat), .B(G155gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G211gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n249), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n249), .B2(new_n253), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n203), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(new_n253), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n255), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n249), .A2(new_n253), .A3(new_n256), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(new_n202), .A3(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(G232gat), .A2(G233gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(KEYINPUT41), .ZN(new_n266));
  XNOR2_X1  g065(.A(G134gat), .B(G162gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G190gat), .B(G218gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G85gat), .ZN(new_n272));
  INV_X1    g071(.A(G92gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G99gat), .ZN(new_n275));
  INV_X1    g074(.A(G106gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT8), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G85gat), .A2(G92gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n278), .A2(KEYINPUT7), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(KEYINPUT7), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n274), .B(new_n277), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G99gat), .B(G106gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n278), .B(KEYINPUT7), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n285), .A2(new_n282), .A3(new_n274), .A4(new_n277), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n288));
  INV_X1    g087(.A(G50gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G43gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G50gat), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT15), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR3_X1   g093(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT84), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT84), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n298), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n289), .A2(G43gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(new_n293), .A3(KEYINPUT15), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G29gat), .ZN(new_n304));
  INV_X1    g103(.A(G36gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR4_X1   g105(.A1(new_n294), .A2(new_n300), .A3(new_n303), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n299), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n305), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(KEYINPUT14), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n295), .A2(KEYINPUT85), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n306), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n302), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n307), .A2(new_n315), .A3(KEYINPUT17), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n303), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n300), .A2(new_n303), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n291), .A2(new_n293), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT15), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n314), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n317), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n287), .B1(new_n316), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT94), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n265), .A2(KEYINPUT41), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n326), .A2(KEYINPUT94), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n307), .A2(new_n315), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(new_n287), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n271), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NOR4_X1   g134(.A1(new_n329), .A2(new_n330), .A3(new_n270), .A4(new_n333), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n269), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n331), .A2(new_n271), .A3(new_n334), .ZN(new_n338));
  INV_X1    g137(.A(new_n330), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n339), .A2(new_n334), .A3(new_n327), .A4(new_n328), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n270), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(new_n341), .A3(new_n268), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n264), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G230gat), .A2(G233gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n234), .A2(new_n287), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n225), .A2(new_n227), .A3(KEYINPUT93), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n232), .B1(new_n231), .B2(new_n226), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n349), .A2(new_n224), .A3(new_n286), .A4(new_n284), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n345), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G120gat), .B(G148gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G176gat), .B(G204gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT96), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n346), .A2(new_n358), .A3(new_n350), .ZN(new_n359));
  INV_X1    g158(.A(new_n287), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n360), .A2(KEYINPUT10), .A3(new_n349), .A4(new_n224), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT95), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n359), .B2(new_n361), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n357), .B1(new_n365), .B2(new_n345), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n359), .A2(new_n361), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT95), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n368), .A2(new_n357), .A3(new_n345), .A4(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n352), .B(new_n356), .C1(new_n366), .C2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n345), .B(KEYINPUT97), .Z(new_n373));
  NAND2_X1  g172(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT98), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n367), .A2(KEYINPUT98), .A3(new_n373), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n352), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n355), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT91), .ZN(new_n381));
  NAND2_X1  g180(.A1(G229gat), .A2(G233gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT13), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n214), .B1(new_n241), .B2(new_n242), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n319), .A2(new_n324), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n239), .A2(G8gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT88), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n240), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n332), .B1(new_n391), .B2(new_n214), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n384), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT90), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n385), .A2(new_n386), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n332), .A3(new_n214), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT90), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n384), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n214), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n390), .B2(new_n240), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n316), .B2(new_n325), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n395), .A3(new_n382), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT18), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT18), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n403), .A2(new_n406), .A3(new_n395), .A4(new_n382), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G169gat), .B(G197gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G113gat), .B(G141gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT12), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n400), .A2(new_n408), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n400), .B2(new_n408), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n381), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n414), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n405), .A2(new_n407), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n398), .B1(new_n397), .B2(new_n384), .ZN(new_n420));
  AOI211_X1 g219(.A(KEYINPUT90), .B(new_n383), .C1(new_n395), .C2(new_n396), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n418), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n400), .A2(new_n408), .A3(new_n414), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(KEYINPUT91), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(KEYINPUT64), .B(G169gat), .Z(new_n427));
  INV_X1    g226(.A(KEYINPUT23), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G176gat), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT25), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n428), .B1(G169gat), .B2(G176gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(G183gat), .A2(G190gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT24), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n434), .A2(KEYINPUT24), .ZN(new_n436));
  INV_X1    g235(.A(G190gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n244), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n435), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n431), .A2(new_n432), .A3(new_n433), .A4(new_n439), .ZN(new_n440));
  OR3_X1    g239(.A1(new_n428), .A2(G169gat), .A3(G176gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n433), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n432), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT25), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT27), .B(G183gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n437), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT65), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT28), .ZN(new_n448));
  OR3_X1    g247(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n432), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(new_n452), .A3(new_n437), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n448), .A2(new_n434), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n440), .A2(new_n444), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G226gat), .ZN(new_n456));
  INV_X1    g255(.A(G233gat), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(KEYINPUT71), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT71), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n440), .A2(new_n444), .A3(new_n460), .A4(new_n454), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n456), .A2(new_n457), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(KEYINPUT29), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n458), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G197gat), .B(G204gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT22), .ZN(new_n467));
  INV_X1    g266(.A(G211gat), .ZN(new_n468));
  INV_X1    g267(.A(G218gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(G211gat), .B(G218gat), .Z(new_n472));
  XOR2_X1   g271(.A(new_n471), .B(new_n472), .Z(new_n473));
  INV_X1    g272(.A(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(KEYINPUT70), .A3(new_n472), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n465), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT72), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n464), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n459), .B2(new_n461), .ZN(new_n483));
  NOR4_X1   g282(.A1(new_n483), .A2(new_n458), .A3(new_n480), .A4(new_n477), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G8gat), .B(G36gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(new_n273), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT73), .B(G64gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n487), .B(new_n488), .Z(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n459), .A2(new_n463), .A3(new_n461), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n455), .A2(new_n464), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n478), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n481), .A2(new_n485), .A3(new_n490), .A4(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT72), .B1(new_n465), .B2(new_n478), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n498), .A2(new_n484), .A3(new_n493), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT30), .A3(new_n490), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n485), .A3(new_n494), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n489), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n497), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G1gat), .B(G29gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(G85gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT0), .B(G57gat), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n505), .B(new_n506), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n509));
  XOR2_X1   g308(.A(G113gat), .B(G120gat), .Z(new_n510));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G127gat), .B(G134gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT66), .B1(new_n513), .B2(KEYINPUT67), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT1), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n510), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G155gat), .A2(G162gat), .ZN(new_n519));
  INV_X1    g318(.A(G155gat), .ZN(new_n520));
  INV_X1    g319(.A(G162gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G141gat), .B(G148gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n519), .B(new_n522), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n523), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n519), .B1(new_n522), .B2(KEYINPUT2), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n518), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT5), .ZN(new_n531));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT4), .ZN(new_n535));
  INV_X1    g334(.A(new_n518), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n529), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n525), .A2(new_n528), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n518), .A2(KEYINPUT4), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT3), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT76), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n529), .A2(KEYINPUT3), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n536), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(new_n542), .A3(new_n544), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n540), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n532), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n548), .B2(new_n532), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n508), .B(new_n534), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT40), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT39), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n530), .A2(new_n532), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(KEYINPUT81), .ZN(new_n559));
  OAI221_X1 g358(.A(new_n559), .B1(KEYINPUT81), .B2(new_n558), .C1(new_n548), .C2(new_n532), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n547), .A2(new_n545), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(new_n537), .A3(new_n539), .ZN(new_n562));
  INV_X1    g361(.A(new_n532), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n557), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(new_n564), .A3(new_n507), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n555), .B1(new_n556), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n503), .B(new_n566), .C1(new_n556), .C2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(G228gat), .A2(G233gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT29), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n477), .B1(new_n569), .B2(new_n542), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n473), .A2(KEYINPUT29), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n538), .B1(new_n571), .B2(new_n541), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT80), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n541), .B1(new_n478), .B2(KEYINPUT29), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(new_n575), .B2(new_n529), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(G228gat), .A3(G233gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(G78gat), .B(G106gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(G22gat), .B(G50gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  AND3_X1   g381(.A1(new_n574), .A2(new_n577), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n574), .B2(new_n577), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT6), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n549), .B1(new_n562), .B2(new_n563), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n533), .B1(new_n587), .B2(new_n551), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n588), .B2(new_n508), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n589), .A2(new_n555), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n491), .A2(new_n478), .A3(new_n492), .ZN(new_n591));
  OAI211_X1 g390(.A(KEYINPUT37), .B(new_n591), .C1(new_n465), .C2(new_n478), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n499), .B2(KEYINPUT37), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n489), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT78), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n588), .A2(new_n596), .A3(KEYINPUT6), .A4(new_n508), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT78), .B1(new_n554), .B2(new_n586), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n590), .A2(new_n595), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT37), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n501), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n499), .A2(KEYINPUT37), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n490), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n495), .B1(new_n603), .B2(new_n594), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n567), .B(new_n585), .C1(new_n599), .C2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n497), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n500), .A2(new_n502), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(KEYINPUT74), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n598), .B(new_n597), .C1(new_n555), .C2(new_n589), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT74), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n500), .A2(new_n502), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n585), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n455), .A2(new_n536), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT68), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n455), .A2(new_n536), .ZN(new_n617));
  NAND2_X1  g416(.A1(G227gat), .A2(G233gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT68), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n455), .A2(new_n619), .A3(new_n536), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT34), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT32), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n624));
  INV_X1    g423(.A(new_n618), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT33), .B1(new_n624), .B2(new_n625), .ZN(new_n627));
  XNOR2_X1  g426(.A(G15gat), .B(G43gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G71gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n275), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n626), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n622), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n627), .A2(new_n631), .ZN(new_n636));
  INV_X1    g435(.A(new_n626), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n622), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n632), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT36), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT69), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n635), .A2(new_n644), .A3(new_n640), .ZN(new_n645));
  OAI211_X1 g444(.A(KEYINPUT69), .B(new_n622), .C1(new_n633), .C2(new_n634), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(KEYINPUT36), .A3(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n605), .A2(new_n614), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n641), .A2(new_n609), .A3(new_n585), .ZN(new_n650));
  INV_X1    g449(.A(new_n503), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT82), .B(KEYINPUT35), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n609), .A2(new_n611), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n645), .A2(new_n646), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n655), .A2(new_n585), .A3(new_n656), .A4(new_n608), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n654), .B1(new_n657), .B2(KEYINPUT35), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n426), .B1(new_n649), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT92), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g460(.A(KEYINPUT92), .B(new_n426), .C1(new_n649), .C2(new_n658), .ZN(new_n662));
  AOI211_X1 g461(.A(new_n344), .B(new_n380), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n609), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g465(.A1(new_n663), .A2(new_n503), .ZN(new_n667));
  NAND2_X1  g466(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n668));
  OR2_X1    g467(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(G8gat), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n667), .A2(KEYINPUT42), .A3(new_n668), .A4(new_n669), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(G1325gat));
  AOI21_X1  g475(.A(G15gat), .B1(new_n663), .B2(new_n641), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n648), .A2(new_n204), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n663), .B2(new_n678), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n613), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  INV_X1    g481(.A(new_n343), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n649), .B2(new_n658), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n264), .A2(new_n380), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n423), .A2(new_n424), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT99), .Z(new_n690));
  OAI211_X1 g489(.A(KEYINPUT44), .B(new_n683), .C1(new_n649), .C2(new_n658), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n609), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT45), .ZN(new_n694));
  INV_X1    g493(.A(new_n687), .ZN(new_n695));
  AOI211_X1 g494(.A(new_n343), .B(new_n695), .C1(new_n661), .C2(new_n662), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(new_n304), .A3(new_n664), .ZN(new_n697));
  MUX2_X1   g496(.A(KEYINPUT45), .B(new_n694), .S(new_n697), .Z(G1328gat));
  NAND3_X1  g497(.A1(new_n696), .A2(new_n305), .A3(new_n503), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n699), .A2(KEYINPUT46), .ZN(new_n700));
  OAI21_X1  g499(.A(G36gat), .B1(new_n692), .B2(new_n651), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(KEYINPUT46), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(G1329gat));
  AOI21_X1  g502(.A(new_n695), .B1(new_n661), .B2(new_n662), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n288), .A2(new_n290), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n704), .A2(new_n641), .A3(new_n705), .A4(new_n683), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n696), .A2(KEYINPUT100), .A3(new_n641), .A4(new_n705), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n648), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n686), .A2(new_n690), .A3(new_n711), .A4(new_n691), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n705), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n710), .A2(KEYINPUT47), .A3(new_n717), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n708), .A2(new_n709), .B1(new_n715), .B2(new_n712), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(KEYINPUT47), .B2(new_n719), .ZN(G1330gat));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n704), .A2(new_n289), .A3(new_n613), .A4(new_n683), .ZN(new_n722));
  OAI21_X1  g521(.A(G50gat), .B1(new_n692), .B2(new_n585), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n722), .B2(new_n723), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n727), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(KEYINPUT48), .A3(new_n725), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1331gat));
  INV_X1    g530(.A(new_n688), .ZN(new_n732));
  INV_X1    g531(.A(new_n380), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n344), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n732), .B(new_n734), .C1(new_n649), .C2(new_n658), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n609), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n220), .ZN(G1332gat));
  NOR2_X1   g536(.A1(new_n735), .A2(new_n651), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  AND2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n738), .B2(new_n739), .ZN(G1333gat));
  INV_X1    g541(.A(new_n641), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n735), .A2(KEYINPUT103), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT103), .B1(new_n735), .B2(new_n743), .ZN(new_n745));
  AOI21_X1  g544(.A(G71gat), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n735), .A2(new_n648), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n217), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT104), .B(KEYINPUT50), .Z(new_n750));
  XOR2_X1   g549(.A(new_n749), .B(new_n750), .Z(G1334gat));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n585), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n218), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n264), .A2(new_n688), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n686), .A2(new_n380), .A3(new_n691), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n609), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n683), .B(new_n754), .C1(new_n649), .C2(new_n658), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n760), .A2(KEYINPUT105), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n757), .A2(new_n758), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(KEYINPUT105), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n664), .A2(new_n272), .A3(new_n380), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT106), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n756), .B1(new_n764), .B2(new_n766), .ZN(G1336gat));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  OAI21_X1  g567(.A(G92gat), .B1(new_n755), .B2(new_n651), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n651), .A2(G92gat), .A3(new_n733), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n768), .B(new_n769), .C1(new_n764), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n760), .A2(new_n762), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n769), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(KEYINPUT107), .A3(KEYINPUT52), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT107), .B1(new_n775), .B2(KEYINPUT52), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n772), .B1(new_n776), .B2(new_n777), .ZN(G1337gat));
  NOR2_X1   g577(.A1(new_n764), .A2(new_n733), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(new_n275), .A3(new_n641), .ZN(new_n780));
  OAI21_X1  g579(.A(G99gat), .B1(new_n755), .B2(new_n648), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1338gat));
  NOR2_X1   g581(.A1(new_n585), .A2(G106gat), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n761), .A2(new_n380), .A3(new_n763), .A4(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT108), .B(G106gat), .Z(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n755), .B2(new_n585), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(KEYINPUT109), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n380), .A3(new_n783), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n786), .C1(new_n755), .C2(new_n585), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n788), .B1(new_n793), .B2(new_n785), .ZN(G1339gat));
  NAND2_X1  g593(.A1(new_n259), .A2(new_n263), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n367), .A2(new_n373), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT54), .B(new_n797), .C1(new_n366), .C2(new_n371), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT54), .B1(new_n376), .B2(new_n377), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n800), .A3(new_n356), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n367), .A2(KEYINPUT98), .A3(new_n373), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT98), .B1(new_n367), .B2(new_n373), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT110), .B1(new_n805), .B2(new_n355), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n798), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n800), .B1(new_n799), .B2(new_n356), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(KEYINPUT110), .A3(new_n355), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n798), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n809), .A2(new_n688), .A3(new_n372), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n397), .A2(new_n384), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n382), .B1(new_n403), .B2(new_n395), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n413), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n424), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n380), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n683), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n813), .A2(new_n372), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT55), .B1(new_n812), .B2(new_n798), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n822), .A2(new_n823), .A3(new_n343), .A4(new_n818), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n795), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n264), .A2(new_n732), .A3(new_n343), .A4(new_n733), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n613), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n656), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n609), .A2(new_n503), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(G113gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n688), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n827), .A2(new_n641), .A3(new_n829), .ZN(new_n833));
  INV_X1    g632(.A(new_n426), .ZN(new_n834));
  OAI21_X1  g633(.A(G113gat), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(G1340gat));
  INV_X1    g635(.A(G120gat), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n830), .A2(new_n837), .A3(new_n380), .ZN(new_n838));
  OAI21_X1  g637(.A(G120gat), .B1(new_n833), .B2(new_n733), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(G1341gat));
  INV_X1    g639(.A(G127gat), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n833), .A2(new_n841), .A3(new_n795), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n830), .A2(new_n264), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n841), .ZN(G1342gat));
  INV_X1    g643(.A(G134gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n845), .A3(new_n683), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT111), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(KEYINPUT111), .ZN(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n833), .B2(new_n343), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(G1343gat));
  AOI21_X1  g651(.A(new_n585), .B1(new_n825), .B2(new_n826), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n853), .A2(KEYINPUT112), .A3(KEYINPUT57), .ZN(new_n854));
  XNOR2_X1  g653(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n807), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n426), .A2(new_n856), .A3(new_n372), .A4(new_n813), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n683), .B1(new_n857), .B2(new_n820), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n795), .B1(new_n858), .B2(new_n824), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n826), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(KEYINPUT57), .A3(new_n613), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT112), .B1(new_n853), .B2(KEYINPUT57), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n854), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n648), .A2(new_n829), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G141gat), .B1(new_n866), .B2(new_n834), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n865), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n869), .A2(G141gat), .A3(new_n834), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n863), .A2(new_n688), .A3(new_n865), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n872), .A2(new_n873), .A3(G141gat), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n872), .B2(G141gat), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n870), .B(KEYINPUT115), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n871), .B1(new_n877), .B2(new_n868), .ZN(G1344gat));
  NAND2_X1  g677(.A1(new_n825), .A2(new_n826), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n613), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n264), .A2(new_n343), .A3(new_n733), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n859), .B1(new_n426), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n585), .A2(KEYINPUT57), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n880), .A2(KEYINPUT57), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n884), .A2(new_n380), .A3(new_n865), .ZN(new_n885));
  INV_X1    g684(.A(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT59), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n866), .B2(new_n733), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n889), .B2(new_n886), .ZN(new_n890));
  INV_X1    g689(.A(new_n869), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n886), .A3(new_n380), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1345gat));
  AOI21_X1  g692(.A(G155gat), .B1(new_n891), .B2(new_n264), .ZN(new_n894));
  INV_X1    g693(.A(new_n866), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n795), .A2(new_n520), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(G1346gat));
  AOI21_X1  g696(.A(G162gat), .B1(new_n891), .B2(new_n683), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n343), .A2(new_n521), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n895), .B2(new_n899), .ZN(G1347gat));
  NAND3_X1  g699(.A1(new_n641), .A2(new_n609), .A3(new_n503), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT116), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n901), .A2(KEYINPUT116), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n827), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n834), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT117), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n664), .A2(new_n651), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n828), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n427), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n688), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n906), .A2(new_n910), .ZN(G1348gat));
  NOR3_X1   g710(.A1(new_n904), .A2(new_n430), .A3(new_n733), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n380), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n430), .ZN(G1349gat));
  NAND3_X1  g713(.A1(new_n908), .A2(new_n445), .A3(new_n264), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n904), .B2(new_n795), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(KEYINPUT118), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n908), .A2(new_n437), .A3(new_n683), .ZN(new_n919));
  OAI21_X1  g718(.A(G190gat), .B1(new_n904), .B2(new_n343), .ZN(new_n920));
  XOR2_X1   g719(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n921));
  AND2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT120), .Z(G1351gat));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n884), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n648), .A2(new_n907), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n884), .A2(new_n926), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G197gat), .B1(new_n931), .B2(new_n834), .ZN(new_n932));
  NOR4_X1   g731(.A1(new_n880), .A2(G197gat), .A3(new_n732), .A4(new_n928), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT121), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT123), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1352gat));
  NOR2_X1   g738(.A1(new_n880), .A2(new_n928), .ZN(new_n940));
  INV_X1    g739(.A(G204gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n941), .A3(new_n380), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g742(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n943), .B(new_n944), .Z(new_n945));
  OAI21_X1  g744(.A(G204gat), .B1(new_n931), .B2(new_n733), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1353gat));
  NOR3_X1   g746(.A1(new_n415), .A2(new_n416), .A3(new_n381), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT91), .B1(new_n423), .B2(new_n424), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n368), .A2(new_n345), .A3(new_n369), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT96), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n796), .B1(new_n951), .B2(new_n370), .ZN(new_n952));
  AOI22_X1  g751(.A1(new_n811), .A2(new_n810), .B1(new_n952), .B2(KEYINPUT54), .ZN(new_n953));
  INV_X1    g752(.A(new_n855), .ZN(new_n954));
  OAI22_X1  g753(.A1(new_n948), .A2(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n820), .B1(new_n955), .B2(new_n822), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n343), .ZN(new_n957));
  INV_X1    g756(.A(new_n824), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n264), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR4_X1   g758(.A1(new_n795), .A2(new_n426), .A3(new_n683), .A4(new_n380), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n883), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT57), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n961), .B(new_n264), .C1(new_n962), .C2(new_n853), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT125), .B1(new_n963), .B2(new_n928), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n884), .A2(new_n965), .A3(new_n264), .A4(new_n929), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n964), .A2(G211gat), .A3(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n964), .A2(new_n966), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n940), .A2(new_n468), .A3(new_n264), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n971), .A2(KEYINPUT126), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1354gat));
  AOI21_X1  g776(.A(G218gat), .B1(new_n940), .B2(new_n683), .ZN(new_n978));
  INV_X1    g777(.A(new_n931), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n683), .A2(G218gat), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT127), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n978), .B1(new_n979), .B2(new_n981), .ZN(G1355gat));
endmodule


