//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n214), .A2(new_n215), .B1(new_n202), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G68), .B2(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n218), .B1(new_n203), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G20), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g0037(.A1(G58), .A2(G68), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G50), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  AOI211_X1 g0041(.A(new_n213), .B(new_n231), .C1(new_n237), .C2(new_n241), .ZN(G361));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G264), .ZN(new_n248));
  INV_X1    g0048(.A(G270), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G358));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n254), .B(new_n257), .Z(G351));
  OAI21_X1  g0058(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n259), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n264), .B2(new_n223), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n262), .A2(KEYINPUT67), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT67), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n268), .B1(new_n271), .B2(new_n236), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G222), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G223), .A2(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n274), .B(new_n279), .C1(G77), .C2(new_n275), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n266), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G200), .ZN(new_n283));
  INV_X1    g0083(.A(G190), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n236), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n206), .A2(G20), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G50), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n235), .A2(G33), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  INV_X1    g0093(.A(G150), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n297), .A2(KEYINPUT68), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(KEYINPUT68), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n207), .B1(new_n238), .B2(new_n222), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n288), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n291), .B1(G50), .B2(new_n285), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n283), .B1(new_n284), .B2(new_n282), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n304), .B2(new_n303), .ZN(new_n306));
  XOR2_X1   g0106(.A(new_n306), .B(KEYINPUT10), .Z(new_n307));
  NOR2_X1   g0107(.A1(new_n282), .A2(G179), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n282), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n303), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G238), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n261), .B1(new_n264), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT71), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(G226), .A2(G1698), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n228), .B2(G1698), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(new_n275), .B1(G33), .B2(G97), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n273), .B2(new_n319), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n320), .A2(KEYINPUT13), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(KEYINPUT13), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT14), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n326), .A3(G169), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n325), .B(new_n327), .C1(new_n328), .C2(new_n323), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n292), .A2(new_n224), .B1(new_n207), .B2(G68), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT73), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n296), .A2(new_n222), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n288), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT11), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT70), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n285), .B(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G68), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(KEYINPUT12), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT12), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n285), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n336), .A2(new_n302), .A3(new_n290), .ZN(new_n342));
  OAI21_X1  g0142(.A(G68), .B1(new_n342), .B2(new_n340), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n334), .A2(new_n339), .A3(new_n341), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n329), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n323), .A2(G200), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT72), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n323), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n344), .B1(new_n349), .B2(G190), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n261), .B1(new_n264), .B2(new_n225), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n353), .A2(KEYINPUT69), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G238), .A2(G1698), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n275), .B(new_n355), .C1(new_n228), .C2(G1698), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n274), .B(new_n356), .C1(G107), .C2(new_n275), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(KEYINPUT69), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n309), .ZN(new_n360));
  INV_X1    g0160(.A(new_n293), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT65), .B(G20), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n361), .A2(new_n295), .B1(new_n362), .B2(G77), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n292), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n288), .A2(new_n365), .B1(new_n342), .B2(G77), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(G77), .B2(new_n336), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n360), .B(new_n367), .C1(G179), .C2(new_n359), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n359), .A2(G200), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n284), .B2(new_n359), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n368), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(G58), .B(G68), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(G20), .B1(G159), .B2(new_n295), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G33), .ZN(new_n377));
  AOI21_X1  g0177(.A(G20), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT75), .B1(new_n378), .B2(KEYINPUT7), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT75), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n275), .C2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n376), .A2(KEYINPUT74), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT74), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n386), .A3(new_n269), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n362), .B1(new_n387), .B2(new_n377), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n374), .B1(new_n390), .B2(G68), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT76), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n379), .A2(new_n382), .B1(new_n388), .B2(KEYINPUT7), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n373), .B1(new_n393), .B2(new_n338), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n269), .B1(new_n384), .B2(new_n386), .ZN(new_n398));
  INV_X1    g0198(.A(new_n375), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT7), .B1(new_n400), .B2(G20), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n376), .A2(KEYINPUT74), .ZN(new_n403));
  OAI21_X1  g0203(.A(G33), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n375), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(new_n381), .A3(new_n235), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(new_n406), .A3(G68), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT16), .A3(new_n373), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n392), .A2(new_n397), .A3(new_n288), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n289), .A2(new_n290), .A3(new_n361), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n285), .B2(new_n361), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT77), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n223), .A2(G1698), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n400), .B(new_n414), .C1(G223), .C2(G1698), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n269), .A2(new_n214), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n273), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n261), .B1(new_n264), .B2(new_n228), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G179), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n309), .B2(new_n420), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n413), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT18), .ZN(new_n424));
  OAI21_X1  g0224(.A(G200), .B1(new_n418), .B2(new_n419), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n420), .A2(G190), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n409), .A2(new_n425), .A3(new_n426), .A4(new_n412), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NOR4_X1   g0229(.A1(new_n312), .A2(new_n352), .A3(new_n371), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n206), .A2(G33), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n289), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G107), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n435));
  OR3_X1    g0235(.A1(new_n285), .A2(G107), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n435), .B1(new_n285), .B2(G107), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(KEYINPUT23), .A2(G107), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G116), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n362), .A2(new_n444), .B1(new_n207), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n235), .B(new_n375), .C1(new_n449), .C2(new_n269), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT22), .B1(new_n450), .B2(new_n214), .ZN(new_n451));
  AND2_X1   g0251(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n453));
  OAI21_X1  g0253(.A(G87), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n375), .A2(new_n377), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n454), .A2(new_n455), .A3(new_n362), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n448), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n459));
  XOR2_X1   g0259(.A(new_n459), .B(KEYINPUT84), .Z(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n443), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n404), .A2(G87), .A3(new_n235), .A4(new_n375), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n456), .B1(new_n463), .B2(KEYINPUT22), .ZN(new_n464));
  NOR4_X1   g0264(.A1(new_n464), .A2(new_n442), .A3(new_n460), .A4(new_n448), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n441), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g0266(.A(new_n434), .B(new_n440), .C1(new_n466), .C2(new_n288), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n216), .A2(new_n276), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n375), .B(new_n468), .C1(new_n449), .C2(new_n269), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT87), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n404), .A2(G250), .A3(new_n276), .A4(new_n375), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT87), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n404), .A2(new_n472), .A3(new_n375), .A4(new_n468), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G294), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n470), .A2(new_n471), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n475), .A2(KEYINPUT88), .A3(new_n274), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT88), .B1(new_n475), .B2(new_n274), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT89), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n206), .A2(G45), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n263), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n219), .ZN(new_n487));
  INV_X1    g0287(.A(new_n484), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n480), .B1(new_n488), .B2(new_n482), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G274), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n478), .A2(new_n479), .A3(new_n284), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n475), .A2(new_n274), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n475), .A2(KEYINPUT88), .A3(new_n274), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n496), .A2(new_n284), .A3(new_n492), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n492), .ZN(new_n500));
  INV_X1    g0300(.A(G200), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n493), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n467), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n451), .A2(new_n457), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n461), .A3(new_n447), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n442), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n458), .A2(new_n443), .A3(new_n461), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n507), .A2(new_n508), .B1(KEYINPUT85), .B2(KEYINPUT24), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n433), .B(new_n439), .C1(new_n509), .C2(new_n302), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n494), .A2(G179), .A3(new_n492), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n496), .A2(new_n492), .A3(new_n497), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(G169), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n504), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G116), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n337), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n336), .A2(G116), .A3(new_n302), .A4(new_n431), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n235), .B(new_n520), .C1(G33), .C2(new_n202), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n287), .A2(new_n236), .B1(G20), .B2(new_n517), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n521), .A2(KEYINPUT20), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT20), .B1(new_n521), .B2(new_n522), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n518), .B(new_n519), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G257), .A2(G1698), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n276), .A2(G264), .ZN(new_n527));
  NOR4_X1   g0327(.A1(new_n398), .A2(new_n399), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G303), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n275), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n274), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n489), .A2(new_n262), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(G270), .B1(G274), .B2(new_n489), .ZN(new_n533));
  AND4_X1   g0333(.A1(G179), .A2(new_n525), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n533), .A3(KEYINPUT81), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT81), .ZN(new_n536));
  INV_X1    g0336(.A(new_n526), .ZN(new_n537));
  INV_X1    g0337(.A(new_n527), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n404), .A2(new_n375), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n530), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n273), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n490), .B1(new_n486), .B2(new_n249), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND4_X1   g0343(.A1(G169), .A2(new_n535), .A3(new_n543), .A4(new_n525), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n534), .B1(new_n544), .B2(KEYINPUT21), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n535), .A2(new_n543), .A3(new_n525), .A4(G169), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT82), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT82), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n545), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n535), .A2(new_n543), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  INV_X1    g0354(.A(new_n525), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n554), .B(new_n555), .C1(new_n501), .C2(new_n553), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n203), .B1(new_n383), .B2(new_n389), .ZN(new_n558));
  XNOR2_X1  g0358(.A(G97), .B(G107), .ZN(new_n559));
  NOR2_X1   g0359(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(KEYINPUT6), .A2(G107), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(KEYINPUT79), .B2(KEYINPUT6), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n362), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n296), .A2(new_n224), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n566), .A2(KEYINPUT78), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(KEYINPUT78), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n288), .B1(new_n558), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n286), .A2(new_n202), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n432), .A2(G97), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n276), .A2(KEYINPUT4), .A3(G244), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n215), .B2(new_n276), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n275), .ZN(new_n576));
  NOR4_X1   g0376(.A1(new_n398), .A2(new_n225), .A3(new_n399), .A4(G1698), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n520), .B(new_n576), .C1(new_n577), .C2(KEYINPUT4), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n274), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n491), .B1(G257), .B2(new_n532), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(G179), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n309), .B1(new_n579), .B2(new_n580), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n573), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n292), .B2(new_n202), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n404), .A2(G68), .A3(new_n235), .A4(new_n375), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n585), .A2(new_n269), .A3(new_n202), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n588), .A2(new_n362), .B1(G87), .B2(new_n204), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n288), .ZN(new_n591));
  INV_X1    g0391(.A(new_n364), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n432), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n337), .A2(new_n364), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n481), .A2(new_n260), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n480), .A2(new_n215), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n263), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G238), .A2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n225), .B2(G1698), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n446), .B1(new_n400), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n598), .B1(new_n601), .B2(new_n273), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n309), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n328), .B(new_n598), .C1(new_n601), .C2(new_n273), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n595), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n590), .A2(new_n288), .B1(new_n337), .B2(new_n364), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n404), .A2(new_n375), .A3(new_n600), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n273), .B1(new_n445), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n598), .ZN(new_n609));
  OAI21_X1  g0409(.A(G200), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(G190), .B(new_n598), .C1(new_n601), .C2(new_n273), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n432), .A2(G87), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n606), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n564), .A2(new_n362), .B1(KEYINPUT78), .B2(new_n566), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n567), .C1(new_n393), .C2(new_n203), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n616), .A2(new_n288), .B1(G97), .B2(new_n432), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n404), .A2(G244), .A3(new_n276), .A4(new_n375), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT4), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n618), .A2(new_n619), .B1(new_n275), .B2(new_n575), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n273), .B1(new_n620), .B2(new_n520), .ZN(new_n621));
  INV_X1    g0421(.A(new_n580), .ZN(new_n622));
  OAI21_X1  g0422(.A(G200), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n579), .A2(G190), .A3(new_n580), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n617), .A2(new_n623), .A3(new_n571), .A4(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n584), .A2(new_n614), .A3(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(KEYINPUT80), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(KEYINPUT80), .ZN(new_n628));
  NOR4_X1   g0428(.A1(new_n516), .A2(new_n557), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n430), .A2(new_n629), .ZN(G372));
  XNOR2_X1  g0430(.A(new_n368), .B(KEYINPUT92), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n351), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n345), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT93), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(KEYINPUT93), .A3(new_n345), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n428), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n424), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n307), .B1(new_n303), .B2(new_n310), .ZN(new_n640));
  INV_X1    g0440(.A(new_n430), .ZN(new_n641));
  INV_X1    g0441(.A(new_n626), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n504), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n434), .B1(new_n466), .B2(new_n288), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n513), .B1(new_n644), .B2(new_n439), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n545), .A2(new_n549), .A3(new_n551), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT90), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n605), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT91), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT91), .ZN(new_n651));
  OAI21_X1  g0451(.A(G169), .B1(new_n621), .B2(new_n622), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n581), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n613), .B(new_n573), .C1(new_n650), .C2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n584), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n613), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n649), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n552), .A2(new_n515), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n626), .B1(new_n467), .B2(new_n503), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n648), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n640), .B1(new_n641), .B2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(new_n516), .ZN(new_n667));
  INV_X1    g0467(.A(G13), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n362), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n206), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n667), .B1(new_n467), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n515), .B2(new_n676), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n676), .A2(new_n555), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n646), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n557), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n660), .A2(new_n504), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n676), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT94), .Z(G399));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n657), .A2(KEYINPUT26), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n613), .B(new_n691), .C1(new_n685), .C2(new_n657), .ZN(new_n692));
  INV_X1    g0492(.A(new_n625), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n605), .B(new_n690), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n689), .B1(new_n694), .B2(new_n676), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n665), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n602), .A2(new_n541), .A3(new_n542), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(new_n494), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n581), .A2(new_n487), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT30), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT96), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT96), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n553), .B1(new_n579), .B2(new_n580), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(new_n328), .A3(new_n602), .A4(new_n500), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT30), .B1(new_n700), .B2(new_n701), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n675), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  XOR2_X1   g0509(.A(KEYINPUT95), .B(KEYINPUT31), .Z(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n629), .B2(new_n676), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n698), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n697), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(KEYINPUT97), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(KEYINPUT97), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n206), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n210), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G1), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n214), .A2(new_n202), .A3(new_n203), .A4(new_n517), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n726), .A2(new_n727), .B1(new_n240), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n722), .A2(new_n729), .ZN(G364));
  XOR2_X1   g0530(.A(new_n682), .B(KEYINPUT98), .Z(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n726), .B1(G45), .B2(new_n669), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n732), .B(new_n734), .C1(G330), .C2(new_n681), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n236), .B1(G20), .B2(new_n309), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n235), .A2(G190), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(G179), .A3(new_n501), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT101), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT101), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n328), .A2(new_n284), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n362), .A2(new_n501), .A3(new_n744), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n743), .A2(new_n224), .B1(new_n227), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT102), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n362), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n202), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n738), .A2(new_n748), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G159), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT32), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n501), .A2(G179), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n738), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n203), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n738), .A2(G179), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n501), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n338), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n757), .A2(new_n455), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n362), .A2(G200), .A3(new_n744), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G50), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n758), .A2(G20), .A3(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G87), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n753), .A2(new_n765), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G294), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n751), .A2(new_n773), .B1(new_n529), .B2(new_n769), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n755), .A2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  XOR2_X1   g0576(.A(KEYINPUT33), .B(G317), .Z(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(new_n776), .B2(new_n759), .C1(new_n763), .C2(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n774), .B(new_n778), .C1(G311), .C2(new_n740), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n767), .A2(G326), .ZN(new_n780));
  INV_X1    g0580(.A(new_n745), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G322), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n779), .A2(new_n455), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n737), .B1(new_n772), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n736), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT100), .Z(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n210), .A2(new_n275), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT99), .Z(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G355), .ZN(new_n793));
  INV_X1    g0593(.A(G45), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n254), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n723), .A2(new_n400), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n240), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n793), .B1(G116), .B2(new_n210), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n784), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n787), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n733), .C1(new_n681), .C2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n735), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  INV_X1    g0603(.A(KEYINPUT105), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n631), .A2(new_n367), .A3(new_n675), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n367), .A2(new_n675), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n371), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n665), .B2(new_n675), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n664), .A2(new_n676), .A3(new_n808), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(KEYINPUT104), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT104), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n664), .A2(new_n813), .A3(new_n676), .A4(new_n808), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n716), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n716), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(new_n734), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n808), .A2(new_n786), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n455), .B1(new_n763), .B2(new_n776), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n752), .B(new_n823), .C1(G107), .C2(new_n770), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n767), .A2(G303), .ZN(new_n825));
  INV_X1    g0625(.A(new_n743), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G116), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n754), .A2(new_n828), .B1(new_n773), .B2(new_n745), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n759), .A2(new_n214), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n824), .A2(new_n825), .A3(new_n827), .A4(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(KEYINPUT103), .B(G143), .Z(new_n833));
  AOI22_X1  g0633(.A1(new_n762), .A2(G150), .B1(new_n781), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  INV_X1    g0635(.A(G159), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n766), .C1(new_n743), .C2(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  INV_X1    g0638(.A(new_n759), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n839), .A2(G68), .B1(G58), .B2(new_n750), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n405), .B1(G50), .B2(new_n770), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n754), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n832), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n736), .A2(new_n785), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n844), .A2(new_n736), .B1(new_n224), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n734), .B1(new_n822), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n804), .B1(new_n820), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n820), .A2(new_n804), .A3(new_n848), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  AOI21_X1  g0653(.A(new_n517), .B1(new_n564), .B2(KEYINPUT35), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n854), .B(new_n237), .C1(KEYINPUT35), .C2(new_n564), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT36), .ZN(new_n856));
  OAI21_X1  g0656(.A(G77), .B1(new_n227), .B2(new_n338), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n240), .A2(new_n857), .B1(G50), .B2(new_n338), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(G1), .A3(new_n668), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n629), .A2(new_n676), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n860), .A2(new_n709), .A3(new_n710), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n709), .A2(KEYINPUT31), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(new_n808), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT16), .B1(new_n407), .B2(new_n373), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT108), .B1(new_n865), .B2(new_n302), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n408), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n865), .A2(KEYINPUT108), .A3(new_n302), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n412), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n673), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n424), .B2(new_n428), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n413), .A2(new_n870), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT109), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT109), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n413), .A2(new_n875), .A3(new_n870), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n423), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(KEYINPUT110), .A3(new_n878), .A4(new_n427), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT110), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n413), .A2(new_n422), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n875), .B1(new_n413), .B2(new_n870), .ZN(new_n882));
  AOI211_X1 g0682(.A(KEYINPUT109), .B(new_n673), .C1(new_n409), .C2(new_n412), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n427), .B(new_n881), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n880), .B1(new_n884), .B2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n869), .A2(new_n422), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n871), .A2(new_n887), .A3(new_n427), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n872), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT38), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n879), .A2(new_n885), .B1(KEYINPUT37), .B2(new_n884), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n883), .B(new_n882), .C1(new_n424), .C2(new_n428), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n352), .A2(new_n344), .A3(new_n675), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n344), .A2(new_n675), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n345), .A2(new_n351), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n864), .A2(KEYINPUT40), .A3(new_n896), .A4(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n879), .A2(new_n885), .B1(KEYINPUT37), .B2(new_n888), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n892), .B1(new_n902), .B2(new_n872), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n891), .A2(new_n903), .ZN(new_n904));
  AND4_X1   g0704(.A1(new_n808), .A2(new_n904), .A3(new_n900), .A4(new_n863), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(KEYINPUT40), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n863), .A2(new_n430), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n906), .B(new_n907), .Z(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(G330), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT106), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n368), .A2(new_n675), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n815), .B2(new_n912), .ZN(new_n913));
  AOI211_X1 g0713(.A(KEYINPUT106), .B(new_n911), .C1(new_n812), .C2(new_n814), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n900), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT107), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(KEYINPUT107), .B(new_n900), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n904), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n424), .A2(new_n870), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n891), .A2(new_n903), .A3(KEYINPUT39), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT39), .B1(new_n891), .B2(new_n895), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n345), .A2(new_n675), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n430), .B1(new_n695), .B2(new_n696), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n640), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n909), .A2(new_n929), .B1(new_n206), .B2(new_n669), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT111), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n909), .A2(new_n929), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n856), .B(new_n859), .C1(new_n931), .C2(new_n932), .ZN(G367));
  NOR2_X1   g0733(.A1(new_n763), .A2(new_n773), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n767), .A2(G311), .B1(G107), .B2(new_n750), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n769), .A2(new_n517), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n935), .B1(KEYINPUT46), .B2(new_n936), .C1(new_n529), .C2(new_n745), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n934), .B(new_n937), .C1(KEYINPUT46), .C2(new_n936), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n839), .A2(G97), .ZN(new_n939));
  INV_X1    g0739(.A(G317), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n939), .B(new_n405), .C1(new_n940), .C2(new_n754), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT112), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n938), .B(new_n942), .C1(new_n776), .C2(new_n743), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n743), .A2(new_n222), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n275), .B1(new_n759), .B2(new_n224), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT113), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n751), .A2(new_n338), .ZN(new_n947));
  INV_X1    g0747(.A(new_n833), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n754), .A2(new_n835), .B1(new_n766), .B2(new_n948), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n947), .B(new_n949), .C1(G150), .C2(new_n781), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n762), .A2(G159), .B1(G58), .B2(new_n770), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n946), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n943), .B1(new_n944), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT47), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n736), .ZN(new_n955));
  INV_X1    g0755(.A(new_n796), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n790), .B1(new_n210), .B2(new_n364), .C1(new_n250), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n606), .A2(new_n612), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n675), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n614), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n605), .B2(new_n959), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(new_n800), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n955), .A2(new_n733), .A3(new_n957), .A4(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n573), .B(new_n675), .C1(new_n650), .C2(new_n653), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n573), .A2(new_n675), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n584), .A2(new_n625), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n552), .A2(new_n675), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n667), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT42), .Z(new_n971));
  AOI21_X1  g0771(.A(new_n657), .B1(new_n968), .B2(new_n645), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n971), .B1(new_n675), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n968), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n684), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n975), .A2(new_n977), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n206), .B1(new_n669), .B2(G45), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n686), .A2(new_n968), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT45), .Z(new_n987));
  NAND3_X1  g0787(.A1(new_n685), .A2(new_n676), .A3(new_n967), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT44), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(new_n684), .ZN(new_n991));
  MUX2_X1   g0791(.A(new_n678), .B(new_n516), .S(new_n969), .Z(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n731), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n683), .B2(new_n992), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n720), .A2(new_n721), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n724), .B(KEYINPUT41), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n985), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n964), .B1(new_n984), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(G387));
  INV_X1    g0800(.A(new_n721), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n994), .B1(new_n1001), .B2(new_n719), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n994), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n720), .A2(new_n721), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1004), .A3(new_n724), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n985), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n994), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n678), .A2(new_n800), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n796), .B1(new_n246), .B2(new_n794), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n792), .A2(new_n727), .ZN(new_n1010));
  AOI211_X1 g0810(.A(G45), .B(new_n727), .C1(G68), .C2(G77), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n293), .A2(G50), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT50), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1009), .A2(new_n1010), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n210), .A2(G107), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n790), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n762), .A2(G311), .B1(G317), .B2(new_n781), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n743), .B2(new_n529), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G322), .B2(new_n767), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT48), .Z(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n776), .B2(new_n751), .C1(new_n773), .C2(new_n769), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT49), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n400), .B1(new_n755), .B2(G326), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n517), .C2(new_n759), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n751), .A2(new_n364), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G159), .B2(new_n767), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n338), .B2(new_n739), .C1(new_n294), .C2(new_n754), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n361), .B2(new_n762), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n781), .A2(G50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n405), .B1(G77), .B2(new_n770), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1028), .A2(new_n939), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n733), .B(new_n1016), .C1(new_n1032), .C2(new_n737), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1008), .B1(new_n1033), .B2(KEYINPUT114), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(KEYINPUT114), .B2(new_n1033), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1005), .A2(new_n1007), .A3(new_n1035), .ZN(G393));
  NAND2_X1  g0836(.A1(new_n991), .A2(new_n1006), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n828), .A2(new_n745), .B1(new_n766), .B2(new_n940), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n203), .B2(new_n759), .C1(new_n529), .C2(new_n763), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G294), .B2(new_n740), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n750), .A2(G116), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n755), .A2(G322), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n275), .B1(new_n770), .B2(G283), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n294), .A2(new_n766), .B1(new_n745), .B2(new_n836), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT51), .Z(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n826), .B2(new_n361), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n751), .A2(new_n224), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n754), .A2(new_n948), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n830), .B(new_n1051), .C1(G50), .C2(new_n762), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n405), .B1(G68), .B2(new_n770), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1048), .A2(new_n1050), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n737), .B1(new_n1045), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n210), .A2(new_n202), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1056), .B(new_n789), .C1(new_n257), .C2(new_n796), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1055), .A2(new_n734), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n968), .B2(new_n800), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1002), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n991), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n724), .B1(new_n1060), .B2(new_n991), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1037), .B(new_n1059), .C1(new_n1062), .C2(new_n1063), .ZN(G390));
  INV_X1    g0864(.A(new_n924), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n923), .B1(new_n915), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n900), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n694), .A2(new_n676), .A3(new_n808), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n912), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n896), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n924), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n716), .A2(new_n808), .A3(new_n900), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n861), .A2(G330), .A3(new_n808), .A4(new_n862), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1073), .A2(KEYINPUT115), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1066), .A2(new_n1071), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(KEYINPUT115), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n923), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n815), .A2(new_n912), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(KEYINPUT106), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n815), .A2(new_n910), .A3(new_n912), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1067), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1079), .B1(new_n1083), .B2(new_n924), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1071), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1078), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1006), .B1(new_n1075), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT118), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n923), .A2(new_n786), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n845), .A2(new_n293), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  XOR2_X1   g0891(.A(KEYINPUT54), .B(G143), .Z(new_n1092));
  AOI22_X1  g0892(.A1(new_n826), .A2(new_n1092), .B1(G137), .B2(new_n762), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(KEYINPUT116), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n770), .A2(G150), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT117), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT53), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1096), .A2(new_n1097), .B1(G132), .B2(new_n781), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n766), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1094), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1093), .A2(KEYINPUT116), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n755), .A2(G125), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1096), .A2(new_n1097), .B1(new_n836), .B2(new_n751), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n455), .B(new_n1104), .C1(G50), .C2(new_n839), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n762), .A2(G107), .B1(G116), .B2(new_n781), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n338), .B2(new_n759), .C1(new_n776), .C2(new_n766), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1049), .B(new_n1108), .C1(G97), .C2(new_n826), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n755), .A2(G294), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1109), .A2(new_n455), .A3(new_n771), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n737), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1112));
  NOR4_X1   g0912(.A1(new_n1089), .A2(new_n734), .A3(new_n1091), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1087), .A2(new_n1088), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n900), .B1(new_n716), .B2(new_n808), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1076), .A2(new_n1116), .B1(new_n913), .B2(new_n914), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1072), .A2(new_n912), .A3(new_n1068), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n863), .A2(new_n430), .A3(G330), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n640), .A2(new_n927), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1075), .B2(new_n1086), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1074), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1072), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1084), .A2(new_n1085), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1123), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n1120), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1077), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1125), .A2(new_n724), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n985), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1134));
  OAI21_X1  g0934(.A(KEYINPUT118), .B1(new_n1134), .B2(new_n1113), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1115), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT119), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1115), .A2(new_n1133), .A3(new_n1135), .A4(KEYINPUT119), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(G378));
  NAND2_X1  g0940(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n901), .B(G330), .C1(KEYINPUT40), .C2(new_n905), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n919), .A2(new_n1142), .A3(new_n925), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n919), .B2(new_n925), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n303), .A2(new_n870), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n312), .B(new_n1146), .Z(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1148));
  XNOR2_X1  g0948(.A(new_n1147), .B(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1149), .B(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1144), .A2(new_n1145), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1149), .B(new_n1150), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1142), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n926), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1154), .B1(new_n1156), .B2(new_n1143), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1141), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1141), .B(KEYINPUT57), .C1(new_n1153), .C2(new_n1157), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n724), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1154), .A2(new_n785), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n269), .A2(new_n270), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT120), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n222), .B(new_n1166), .C1(new_n400), .C2(G41), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n745), .A2(new_n1099), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n767), .A2(G125), .B1(G150), .B2(new_n750), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT121), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n770), .C2(new_n1092), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n842), .B2(new_n763), .C1(new_n835), .C2(new_n739), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT59), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1166), .B1(new_n755), .B2(G124), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n836), .B2(new_n759), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1167), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n759), .A2(new_n227), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n781), .A2(G107), .B1(G77), .B2(new_n770), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n517), .B2(new_n766), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(G97), .C2(new_n762), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n755), .A2(G283), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n947), .A2(G41), .A3(new_n400), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n740), .A2(new_n592), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT58), .Z(new_n1185));
  OAI21_X1  g0985(.A(new_n736), .B1(new_n1176), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n845), .A2(new_n222), .ZN(new_n1187));
  AND4_X1   g0987(.A1(new_n733), .A2(new_n1164), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1189), .B2(new_n1006), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1163), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(G375));
  NAND2_X1  g0993(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n1130), .A3(new_n996), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1177), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n835), .B2(new_n745), .C1(new_n836), .C2(new_n769), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n762), .B2(new_n1092), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n842), .B2(new_n766), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n405), .B(new_n1199), .C1(G150), .C2(new_n740), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n222), .B2(new_n751), .C1(new_n1099), .C2(new_n754), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n455), .B1(new_n759), .B2(new_n224), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT125), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1025), .B(new_n1203), .C1(G303), .C2(new_n755), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n767), .A2(G294), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n826), .A2(G107), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n762), .A2(G116), .B1(G283), .B2(new_n781), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n769), .A2(new_n202), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1201), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n736), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n733), .B(new_n1211), .C1(new_n900), .C2(new_n786), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n338), .B2(new_n845), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n985), .B(KEYINPUT124), .Z(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1120), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1195), .A2(new_n1215), .ZN(G381));
  INV_X1    g1016(.A(new_n1136), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1192), .A2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1005), .A2(new_n802), .A3(new_n1007), .A4(new_n1035), .ZN(new_n1219));
  OR3_X1    g1019(.A1(G387), .A2(G384), .A3(new_n1219), .ZN(new_n1220));
  OR4_X1    g1020(.A1(G390), .A2(new_n1218), .A3(G381), .A4(new_n1220), .ZN(G407));
  OAI211_X1 g1021(.A(G407), .B(G213), .C1(G343), .C2(new_n1218), .ZN(G409));
  NOR2_X1   g1022(.A1(G390), .A2(new_n999), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G390), .A2(new_n999), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(KEYINPUT127), .A3(new_n1219), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(G390), .A2(new_n999), .A3(new_n1219), .A4(new_n1225), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1223), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1226), .A2(new_n999), .A3(G390), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(G343), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT60), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1130), .B(new_n724), .C1(new_n1194), .C2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT60), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1215), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  OR3_X1    g1038(.A1(new_n1237), .A2(new_n1238), .A3(G384), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(G384), .A2(new_n1238), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n852), .A2(KEYINPUT126), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1237), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G378), .A2(new_n1162), .A3(new_n1190), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1214), .B1(new_n1141), .B2(new_n996), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1217), .B1(new_n1248), .B2(new_n1188), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1233), .B(new_n1244), .C1(new_n1245), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1233), .B1(new_n1245), .B2(new_n1249), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1233), .A2(G2897), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1243), .B(new_n1253), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n1250), .A2(new_n1251), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1245), .A2(new_n1249), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1233), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(new_n1251), .A3(new_n1257), .A4(new_n1243), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1231), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1231), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1259), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1250), .B2(KEYINPUT63), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1250), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT63), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1261), .A2(new_n1268), .ZN(G405));
  OAI21_X1  g1069(.A(new_n1217), .B1(new_n1163), .B2(new_n1191), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1262), .B1(new_n1270), .B2(new_n1245), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1262), .A2(new_n1270), .A3(new_n1245), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1244), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1273), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1243), .B1(new_n1275), .B2(new_n1271), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(G402));
endmodule


