

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(G2105), .ZN(n595) );
  NOR2_X1 U551 ( .A1(n603), .A2(n602), .ZN(G164) );
  NOR2_X2 U552 ( .A1(n611), .A2(n610), .ZN(n517) );
  INV_X1 U553 ( .A(KEYINPUT65), .ZN(n516) );
  INV_X1 U554 ( .A(KEYINPUT0), .ZN(n557) );
  NOR2_X1 U555 ( .A1(G2105), .A2(G2104), .ZN(n593) );
  XNOR2_X1 U556 ( .A(n778), .B(n518), .ZN(n521) );
  NAND2_X1 U557 ( .A1(n541), .A2(n538), .ZN(n778) );
  AND2_X1 U558 ( .A1(n535), .A2(n531), .ZN(n530) );
  AND2_X1 U559 ( .A1(n532), .A2(n715), .ZN(n531) );
  XNOR2_X1 U560 ( .A(n726), .B(KEYINPUT31), .ZN(n727) );
  NOR2_X1 U561 ( .A1(G164), .A2(n663), .ZN(n664) );
  BUF_X1 U562 ( .A(n678), .Z(n561) );
  AND2_X1 U563 ( .A1(n623), .A2(G101), .ZN(n607) );
  XNOR2_X1 U564 ( .A(n594), .B(n593), .ZN(n620) );
  XNOR2_X1 U565 ( .A(n557), .B(G543), .ZN(n641) );
  XNOR2_X2 U566 ( .A(n517), .B(n516), .ZN(G160) );
  BUF_X1 U567 ( .A(n620), .Z(n519) );
  INV_X1 U568 ( .A(KEYINPUT101), .ZN(n518) );
  XNOR2_X1 U569 ( .A(n705), .B(n704), .ZN(n537) );
  NAND2_X1 U570 ( .A1(n716), .A2(G8), .ZN(n772) );
  XNOR2_X2 U571 ( .A(n729), .B(KEYINPUT94), .ZN(n742) );
  INV_X1 U572 ( .A(n710), .ZN(n533) );
  XNOR2_X1 U573 ( .A(G305), .B(n766), .ZN(n1050) );
  NAND2_X1 U574 ( .A1(n523), .A2(n552), .ZN(n549) );
  NAND2_X1 U575 ( .A1(n523), .A2(KEYINPUT102), .ZN(n553) );
  NAND2_X1 U576 ( .A1(n811), .A2(n552), .ZN(n551) );
  XNOR2_X1 U577 ( .A(n707), .B(KEYINPUT28), .ZN(n708) );
  INV_X1 U578 ( .A(KEYINPUT90), .ZN(n693) );
  NAND2_X1 U579 ( .A1(n534), .A2(n533), .ZN(n532) );
  INV_X1 U580 ( .A(n708), .ZN(n534) );
  OR2_X1 U581 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U582 ( .A1(n529), .A2(n533), .ZN(n528) );
  XNOR2_X1 U583 ( .A(n757), .B(n756), .ZN(n1048) );
  INV_X1 U584 ( .A(KEYINPUT102), .ZN(n552) );
  INV_X1 U585 ( .A(n765), .ZN(n540) );
  NOR2_X1 U586 ( .A1(n595), .A2(G2104), .ZN(n599) );
  NAND2_X1 U587 ( .A1(n549), .A2(n548), .ZN(n547) );
  NAND2_X1 U588 ( .A1(n811), .A2(KEYINPUT102), .ZN(n548) );
  NOR2_X1 U589 ( .A1(n526), .A2(n546), .ZN(n545) );
  INV_X1 U590 ( .A(n554), .ZN(n546) );
  XNOR2_X1 U591 ( .A(G168), .B(n592), .ZN(G286) );
  NOR2_X2 U592 ( .A1(n641), .A2(n559), .ZN(n520) );
  OR2_X1 U593 ( .A1(n706), .A2(G299), .ZN(n522) );
  OR2_X1 U594 ( .A1(n810), .A2(KEYINPUT103), .ZN(n523) );
  OR2_X1 U595 ( .A1(n772), .A2(KEYINPUT33), .ZN(n524) );
  NAND2_X1 U596 ( .A1(n744), .A2(n743), .ZN(n525) );
  AND2_X1 U597 ( .A1(n553), .A2(n551), .ZN(n526) );
  AND2_X1 U598 ( .A1(n1050), .A2(n542), .ZN(n527) );
  NAND2_X1 U599 ( .A1(n530), .A2(n528), .ZN(n728) );
  INV_X1 U600 ( .A(n537), .ZN(n529) );
  NAND2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n535) );
  AND2_X1 U602 ( .A1(n708), .A2(n710), .ZN(n536) );
  AND2_X1 U603 ( .A1(n777), .A2(n539), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n527), .A2(n540), .ZN(n539) );
  NAND2_X1 U605 ( .A1(n761), .A2(n527), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n765), .A2(n524), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n521), .A2(n554), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n550), .A2(n543), .ZN(n827) );
  NAND2_X1 U609 ( .A1(n544), .A2(n547), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n521), .A2(n545), .ZN(n550) );
  INV_X2 U611 ( .A(n716), .ZN(n666) );
  NAND2_X2 U612 ( .A1(G160), .A2(n664), .ZN(n716) );
  NAND2_X1 U613 ( .A1(n807), .A2(n824), .ZN(n554) );
  AND2_X1 U614 ( .A1(n661), .A2(n660), .ZN(n555) );
  AND2_X1 U615 ( .A1(n716), .A2(n668), .ZN(n556) );
  OR2_X1 U616 ( .A1(n716), .A2(n696), .ZN(n699) );
  XNOR2_X1 U617 ( .A(KEYINPUT30), .B(KEYINPUT93), .ZN(n719) );
  XNOR2_X1 U618 ( .A(n720), .B(n719), .ZN(n722) );
  NOR2_X1 U619 ( .A1(n657), .A2(n656), .ZN(n659) );
  NOR2_X1 U620 ( .A1(n618), .A2(n617), .ZN(G171) );
  INV_X1 U621 ( .A(G651), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G73), .A2(n520), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT2), .B(n558), .Z(n567) );
  NOR2_X1 U624 ( .A1(G543), .A2(n559), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT1), .B(n560), .Z(n678) );
  NAND2_X1 U626 ( .A1(n561), .A2(G61), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT82), .ZN(n564) );
  NOR2_X2 U628 ( .A1(G651), .A2(G543), .ZN(n844) );
  NAND2_X1 U629 ( .A1(G86), .A2(n844), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT83), .B(n565), .Z(n566) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n571) );
  NOR2_X1 U633 ( .A1(n641), .A2(G651), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT64), .ZN(n653) );
  INV_X1 U635 ( .A(n653), .ZN(n569) );
  INV_X1 U636 ( .A(n569), .ZN(n847) );
  NAND2_X1 U637 ( .A1(G48), .A2(n847), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(G305) );
  NAND2_X1 U639 ( .A1(G65), .A2(n561), .ZN(n573) );
  NAND2_X1 U640 ( .A1(G53), .A2(n847), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U642 ( .A(KEYINPUT70), .B(n574), .Z(n578) );
  NAND2_X1 U643 ( .A1(G91), .A2(n844), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G78), .A2(n520), .ZN(n575) );
  AND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(G299) );
  XNOR2_X1 U647 ( .A(KEYINPUT6), .B(KEYINPUT76), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G63), .A2(n561), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G51), .A2(n847), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U651 ( .A(n582), .B(n581), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n520), .A2(G76), .ZN(n583) );
  XNOR2_X1 U653 ( .A(KEYINPUT75), .B(n583), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n844), .A2(G89), .ZN(n584) );
  XOR2_X1 U655 ( .A(KEYINPUT4), .B(n584), .Z(n585) );
  NOR2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U657 ( .A(n587), .B(KEYINPUT5), .ZN(n588) );
  NOR2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U659 ( .A(n590), .B(KEYINPUT7), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT77), .ZN(G168) );
  INV_X1 U661 ( .A(KEYINPUT8), .ZN(n592) );
  XNOR2_X2 U662 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n620), .A2(G138), .ZN(n597) );
  AND2_X4 U664 ( .A1(n595), .A2(G2104), .ZN(n623) );
  NAND2_X1 U665 ( .A1(G102), .A2(n623), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT86), .ZN(n603) );
  AND2_X1 U668 ( .A1(G2105), .A2(G2104), .ZN(n936) );
  NAND2_X1 U669 ( .A1(G114), .A2(n936), .ZN(n601) );
  XNOR2_X2 U670 ( .A(n599), .B(KEYINPUT66), .ZN(n937) );
  NAND2_X1 U671 ( .A1(G126), .A2(n937), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n620), .A2(G137), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n936), .A2(G113), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(KEYINPUT68), .ZN(n611) );
  XNOR2_X1 U677 ( .A(n607), .B(KEYINPUT23), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n937), .A2(G125), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G90), .A2(n844), .ZN(n613) );
  NAND2_X1 U681 ( .A1(G77), .A2(n520), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U683 ( .A(KEYINPUT9), .B(n614), .Z(n618) );
  NAND2_X1 U684 ( .A1(G64), .A2(n561), .ZN(n616) );
  NAND2_X1 U685 ( .A1(G52), .A2(n847), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n616), .A2(n615), .ZN(n617) );
  AND2_X1 U687 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U688 ( .A1(G123), .A2(n937), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n619), .B(KEYINPUT18), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n519), .A2(G135), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n628) );
  NAND2_X1 U692 ( .A1(G111), .A2(n936), .ZN(n625) );
  NAND2_X1 U693 ( .A1(G99), .A2(n623), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U695 ( .A(KEYINPUT78), .B(n626), .ZN(n627) );
  NOR2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n629), .B(KEYINPUT79), .ZN(n986) );
  XNOR2_X1 U698 ( .A(G2096), .B(n986), .ZN(n630) );
  OR2_X1 U699 ( .A1(G2100), .A2(n630), .ZN(G156) );
  INV_X1 U700 ( .A(G132), .ZN(G219) );
  INV_X1 U701 ( .A(G82), .ZN(G220) );
  INV_X1 U702 ( .A(G171), .ZN(G301) );
  NAND2_X1 U703 ( .A1(G88), .A2(n844), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G75), .A2(n520), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n847), .A2(G50), .ZN(n633) );
  XOR2_X1 U707 ( .A(KEYINPUT84), .B(n633), .Z(n634) );
  NOR2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n561), .A2(G62), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n637), .A2(n636), .ZN(G303) );
  NAND2_X1 U711 ( .A1(G651), .A2(G74), .ZN(n639) );
  NAND2_X1 U712 ( .A1(G49), .A2(n847), .ZN(n638) );
  NAND2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U714 ( .A1(n561), .A2(n640), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n641), .A2(G87), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n643), .A2(n642), .ZN(G288) );
  NAND2_X1 U717 ( .A1(G85), .A2(n844), .ZN(n645) );
  NAND2_X1 U718 ( .A1(G72), .A2(n520), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U720 ( .A(KEYINPUT69), .B(n646), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n847), .A2(G47), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G60), .A2(n561), .ZN(n647) );
  AND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(G290) );
  NAND2_X1 U725 ( .A1(G92), .A2(n844), .ZN(n652) );
  NAND2_X1 U726 ( .A1(G66), .A2(n678), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n657) );
  NAND2_X1 U728 ( .A1(G54), .A2(n653), .ZN(n655) );
  NAND2_X1 U729 ( .A1(G79), .A2(n520), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U731 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n658) );
  XNOR2_X2 U732 ( .A(n659), .B(n658), .ZN(n689) );
  NAND2_X1 U733 ( .A1(n689), .A2(G2067), .ZN(n661) );
  NAND2_X1 U734 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n660) );
  INV_X1 U735 ( .A(G40), .ZN(n662) );
  OR2_X1 U736 ( .A1(n662), .A2(G1384), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n555), .A2(n666), .ZN(n671) );
  INV_X1 U738 ( .A(G1341), .ZN(n667) );
  AND2_X1 U739 ( .A1(n667), .A2(KEYINPUT26), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n689), .A2(G1348), .ZN(n669) );
  NAND2_X1 U741 ( .A1(n556), .A2(n669), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n684) );
  NAND2_X1 U743 ( .A1(n844), .A2(G81), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n672), .B(KEYINPUT12), .ZN(n674) );
  NAND2_X1 U745 ( .A1(G68), .A2(n520), .ZN(n673) );
  NAND2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U747 ( .A(KEYINPUT13), .B(n675), .Z(n677) );
  AND2_X1 U748 ( .A1(n847), .A2(G43), .ZN(n676) );
  NOR2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n681) );
  NAND2_X1 U750 ( .A1(G56), .A2(n678), .ZN(n679) );
  XNOR2_X1 U751 ( .A(KEYINPUT14), .B(n679), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n1045) );
  NOR2_X1 U753 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n682) );
  NOR2_X1 U754 ( .A1(n1045), .A2(n682), .ZN(n683) );
  NAND2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n692) );
  INV_X1 U756 ( .A(G2067), .ZN(n685) );
  NAND2_X1 U757 ( .A1(n666), .A2(n685), .ZN(n688) );
  INV_X1 U758 ( .A(G1348), .ZN(n686) );
  NAND2_X1 U759 ( .A1(n716), .A2(n686), .ZN(n687) );
  NAND2_X1 U760 ( .A1(n688), .A2(n687), .ZN(n690) );
  INV_X1 U761 ( .A(n689), .ZN(n853) );
  NAND2_X1 U762 ( .A1(n690), .A2(n853), .ZN(n691) );
  NAND2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n694) );
  XNOR2_X1 U764 ( .A(n694), .B(n693), .ZN(n703) );
  INV_X1 U765 ( .A(KEYINPUT27), .ZN(n695) );
  AND2_X1 U766 ( .A1(n695), .A2(G2072), .ZN(n696) );
  NOR2_X1 U767 ( .A1(KEYINPUT27), .A2(G1956), .ZN(n697) );
  NAND2_X1 U768 ( .A1(n716), .A2(n697), .ZN(n698) );
  NAND2_X1 U769 ( .A1(n699), .A2(n698), .ZN(n702) );
  INV_X1 U770 ( .A(G2072), .ZN(n700) );
  NAND2_X1 U771 ( .A1(n700), .A2(KEYINPUT27), .ZN(n701) );
  NAND2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n703), .A2(n522), .ZN(n705) );
  INV_X1 U774 ( .A(KEYINPUT91), .ZN(n704) );
  NAND2_X1 U775 ( .A1(n706), .A2(G299), .ZN(n707) );
  INV_X1 U776 ( .A(KEYINPUT92), .ZN(n709) );
  XNOR2_X1 U777 ( .A(n709), .B(KEYINPUT29), .ZN(n710) );
  XOR2_X1 U778 ( .A(G2078), .B(KEYINPUT25), .Z(n1026) );
  INV_X1 U779 ( .A(n1026), .ZN(n711) );
  OR2_X1 U780 ( .A1(n716), .A2(n711), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n716), .A2(G1961), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n723) );
  INV_X1 U783 ( .A(n723), .ZN(n714) );
  NAND2_X1 U784 ( .A1(n714), .A2(G171), .ZN(n715) );
  OR2_X1 U785 ( .A1(n772), .A2(G1966), .ZN(n744) );
  INV_X1 U786 ( .A(G2084), .ZN(n717) );
  NAND2_X1 U787 ( .A1(n666), .A2(n717), .ZN(n743) );
  AND2_X1 U788 ( .A1(n743), .A2(G8), .ZN(n718) );
  NAND2_X1 U789 ( .A1(n744), .A2(n718), .ZN(n720) );
  INV_X1 U790 ( .A(G168), .ZN(n721) );
  NAND2_X1 U791 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U792 ( .A1(n723), .A2(G301), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U795 ( .A1(n742), .A2(G286), .ZN(n731) );
  INV_X1 U796 ( .A(KEYINPUT95), .ZN(n730) );
  XNOR2_X1 U797 ( .A(n731), .B(n730), .ZN(n737) );
  NOR2_X1 U798 ( .A1(n716), .A2(G2090), .ZN(n732) );
  XNOR2_X1 U799 ( .A(n732), .B(KEYINPUT96), .ZN(n735) );
  OR2_X1 U800 ( .A1(n772), .A2(G1971), .ZN(n733) );
  NAND2_X1 U801 ( .A1(n733), .A2(G303), .ZN(n734) );
  NAND2_X1 U802 ( .A1(n737), .A2(n736), .ZN(n739) );
  INV_X1 U803 ( .A(KEYINPUT97), .ZN(n738) );
  XNOR2_X1 U804 ( .A(n739), .B(n738), .ZN(n740) );
  NAND2_X1 U805 ( .A1(n740), .A2(G8), .ZN(n741) );
  XNOR2_X1 U806 ( .A(n741), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U807 ( .A1(n525), .A2(G8), .ZN(n746) );
  INV_X1 U808 ( .A(KEYINPUT89), .ZN(n745) );
  NAND2_X1 U809 ( .A1(n746), .A2(n745), .ZN(n750) );
  NAND2_X1 U810 ( .A1(G8), .A2(KEYINPUT89), .ZN(n747) );
  NOR2_X1 U811 ( .A1(n747), .A2(G2084), .ZN(n748) );
  NAND2_X1 U812 ( .A1(n666), .A2(n748), .ZN(n749) );
  NAND2_X1 U813 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U814 ( .A1(n742), .A2(n751), .ZN(n752) );
  NAND2_X1 U815 ( .A1(n753), .A2(n752), .ZN(n767) );
  NOR2_X1 U816 ( .A1(G1971), .A2(G303), .ZN(n754) );
  NOR2_X1 U817 ( .A1(G1976), .A2(G288), .ZN(n762) );
  NOR2_X1 U818 ( .A1(n754), .A2(n762), .ZN(n1061) );
  XNOR2_X1 U819 ( .A(KEYINPUT98), .B(n1061), .ZN(n755) );
  NAND2_X1 U820 ( .A1(n767), .A2(n755), .ZN(n758) );
  NAND2_X1 U821 ( .A1(G288), .A2(G1976), .ZN(n757) );
  INV_X1 U822 ( .A(KEYINPUT99), .ZN(n756) );
  NAND2_X1 U823 ( .A1(n758), .A2(n1048), .ZN(n760) );
  INV_X1 U824 ( .A(KEYINPUT100), .ZN(n759) );
  XNOR2_X1 U825 ( .A(n760), .B(n759), .ZN(n761) );
  INV_X1 U826 ( .A(n762), .ZN(n763) );
  OR2_X1 U827 ( .A1(n772), .A2(n763), .ZN(n764) );
  NAND2_X1 U828 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  INV_X1 U829 ( .A(G1981), .ZN(n766) );
  NOR2_X1 U830 ( .A1(G2090), .A2(G303), .ZN(n768) );
  NAND2_X1 U831 ( .A1(G8), .A2(n768), .ZN(n769) );
  AND2_X1 U832 ( .A1(n769), .A2(n772), .ZN(n770) );
  NAND2_X1 U833 ( .A1(n767), .A2(n770), .ZN(n776) );
  OR2_X1 U834 ( .A1(G305), .A2(G1981), .ZN(n771) );
  XNOR2_X1 U835 ( .A(n771), .B(KEYINPUT24), .ZN(n774) );
  INV_X1 U836 ( .A(n772), .ZN(n773) );
  NAND2_X1 U837 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U838 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U839 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NAND2_X1 U840 ( .A1(n519), .A2(G140), .ZN(n780) );
  NAND2_X1 U841 ( .A1(G104), .A2(n623), .ZN(n779) );
  NAND2_X1 U842 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U843 ( .A(KEYINPUT34), .B(n781), .ZN(n786) );
  NAND2_X1 U844 ( .A1(G116), .A2(n936), .ZN(n783) );
  NAND2_X1 U845 ( .A1(G128), .A2(n937), .ZN(n782) );
  NAND2_X1 U846 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U847 ( .A(KEYINPUT35), .B(n784), .Z(n785) );
  NOR2_X1 U848 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U849 ( .A(KEYINPUT36), .B(n787), .ZN(n912) );
  NOR2_X1 U850 ( .A1(n820), .A2(n912), .ZN(n974) );
  NAND2_X1 U851 ( .A1(n937), .A2(G119), .ZN(n794) );
  NAND2_X1 U852 ( .A1(n519), .A2(G131), .ZN(n789) );
  NAND2_X1 U853 ( .A1(n936), .A2(G107), .ZN(n788) );
  NAND2_X1 U854 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U855 ( .A1(G95), .A2(n623), .ZN(n790) );
  XNOR2_X1 U856 ( .A(KEYINPUT87), .B(n790), .ZN(n791) );
  NOR2_X1 U857 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U858 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U859 ( .A(n795), .B(KEYINPUT88), .ZN(n915) );
  NAND2_X1 U860 ( .A1(G1991), .A2(n915), .ZN(n804) );
  NAND2_X1 U861 ( .A1(n937), .A2(G129), .ZN(n797) );
  NAND2_X1 U862 ( .A1(n519), .A2(G141), .ZN(n796) );
  NAND2_X1 U863 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U864 ( .A1(n623), .A2(G105), .ZN(n798) );
  XOR2_X1 U865 ( .A(KEYINPUT38), .B(n798), .Z(n799) );
  NOR2_X1 U866 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U867 ( .A1(n936), .A2(G117), .ZN(n801) );
  NAND2_X1 U868 ( .A1(n802), .A2(n801), .ZN(n914) );
  NAND2_X1 U869 ( .A1(G1996), .A2(n914), .ZN(n803) );
  NAND2_X1 U870 ( .A1(n804), .A2(n803), .ZN(n973) );
  OR2_X1 U871 ( .A1(n974), .A2(n973), .ZN(n807) );
  OR2_X1 U872 ( .A1(G164), .A2(G1384), .ZN(n805) );
  AND2_X1 U873 ( .A1(n805), .A2(G40), .ZN(n806) );
  AND2_X1 U874 ( .A1(n806), .A2(G160), .ZN(n824) );
  XNOR2_X1 U875 ( .A(G290), .B(G1986), .ZN(n1059) );
  INV_X1 U876 ( .A(n1059), .ZN(n809) );
  INV_X1 U877 ( .A(n824), .ZN(n808) );
  NOR2_X1 U878 ( .A1(n809), .A2(n808), .ZN(n810) );
  INV_X1 U879 ( .A(KEYINPUT103), .ZN(n811) );
  NOR2_X1 U880 ( .A1(G1996), .A2(n914), .ZN(n970) );
  NOR2_X1 U881 ( .A1(n915), .A2(G1991), .ZN(n987) );
  NOR2_X1 U882 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U883 ( .A1(n987), .A2(n812), .ZN(n813) );
  NOR2_X1 U884 ( .A1(n973), .A2(n813), .ZN(n814) );
  XNOR2_X1 U885 ( .A(n814), .B(KEYINPUT104), .ZN(n815) );
  NOR2_X1 U886 ( .A1(n970), .A2(n815), .ZN(n816) );
  XNOR2_X1 U887 ( .A(n816), .B(KEYINPUT39), .ZN(n818) );
  INV_X1 U888 ( .A(n974), .ZN(n817) );
  NAND2_X1 U889 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U890 ( .A(KEYINPUT105), .B(n819), .Z(n823) );
  NAND2_X1 U891 ( .A1(n820), .A2(n912), .ZN(n975) );
  NAND2_X1 U892 ( .A1(n1059), .A2(KEYINPUT103), .ZN(n821) );
  AND2_X1 U893 ( .A1(n975), .A2(n821), .ZN(n822) );
  NAND2_X1 U894 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U895 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U896 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U897 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U898 ( .A1(G7), .A2(G661), .ZN(n829) );
  XNOR2_X1 U899 ( .A(n829), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U900 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n831) );
  INV_X1 U901 ( .A(G223), .ZN(n880) );
  NAND2_X1 U902 ( .A1(G567), .A2(n880), .ZN(n830) );
  XNOR2_X1 U903 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U904 ( .A(KEYINPUT72), .B(n832), .Z(G234) );
  INV_X1 U905 ( .A(G860), .ZN(n837) );
  OR2_X1 U906 ( .A1(n1045), .A2(n837), .ZN(G153) );
  NOR2_X1 U907 ( .A1(n689), .A2(G868), .ZN(n834) );
  INV_X1 U908 ( .A(G868), .ZN(n863) );
  NOR2_X1 U909 ( .A1(n863), .A2(G301), .ZN(n833) );
  NOR2_X1 U910 ( .A1(n834), .A2(n833), .ZN(G284) );
  NOR2_X1 U911 ( .A1(G286), .A2(n863), .ZN(n836) );
  NOR2_X1 U912 ( .A1(G868), .A2(G299), .ZN(n835) );
  NOR2_X1 U913 ( .A1(n836), .A2(n835), .ZN(G297) );
  NAND2_X1 U914 ( .A1(n837), .A2(G559), .ZN(n838) );
  NAND2_X1 U915 ( .A1(n838), .A2(n853), .ZN(n839) );
  XNOR2_X1 U916 ( .A(n839), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U917 ( .A1(G868), .A2(n1045), .ZN(n842) );
  NAND2_X1 U918 ( .A1(n853), .A2(G868), .ZN(n840) );
  NOR2_X1 U919 ( .A1(G559), .A2(n840), .ZN(n841) );
  NOR2_X1 U920 ( .A1(n842), .A2(n841), .ZN(G282) );
  NAND2_X1 U921 ( .A1(G67), .A2(n561), .ZN(n843) );
  XNOR2_X1 U922 ( .A(n843), .B(KEYINPUT80), .ZN(n852) );
  NAND2_X1 U923 ( .A1(G93), .A2(n844), .ZN(n846) );
  NAND2_X1 U924 ( .A1(G80), .A2(n520), .ZN(n845) );
  NAND2_X1 U925 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U926 ( .A1(G55), .A2(n847), .ZN(n848) );
  XNOR2_X1 U927 ( .A(KEYINPUT81), .B(n848), .ZN(n849) );
  NOR2_X1 U928 ( .A1(n850), .A2(n849), .ZN(n851) );
  NAND2_X1 U929 ( .A1(n852), .A2(n851), .ZN(n864) );
  NAND2_X1 U930 ( .A1(n853), .A2(G559), .ZN(n854) );
  XNOR2_X1 U931 ( .A(n854), .B(n1045), .ZN(n861) );
  NOR2_X1 U932 ( .A1(G860), .A2(n861), .ZN(n855) );
  XOR2_X1 U933 ( .A(n864), .B(n855), .Z(G145) );
  INV_X1 U934 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U935 ( .A(G299), .B(G305), .ZN(n860) );
  XNOR2_X1 U936 ( .A(KEYINPUT19), .B(G288), .ZN(n856) );
  XNOR2_X1 U937 ( .A(n856), .B(n864), .ZN(n857) );
  XNOR2_X1 U938 ( .A(G166), .B(n857), .ZN(n858) );
  XNOR2_X1 U939 ( .A(n858), .B(G290), .ZN(n859) );
  XNOR2_X1 U940 ( .A(n860), .B(n859), .ZN(n949) );
  XNOR2_X1 U941 ( .A(n861), .B(n949), .ZN(n862) );
  NAND2_X1 U942 ( .A1(n862), .A2(G868), .ZN(n866) );
  NAND2_X1 U943 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U944 ( .A1(n866), .A2(n865), .ZN(G295) );
  NAND2_X1 U945 ( .A1(G2078), .A2(G2084), .ZN(n867) );
  XOR2_X1 U946 ( .A(KEYINPUT20), .B(n867), .Z(n868) );
  NAND2_X1 U947 ( .A1(G2090), .A2(n868), .ZN(n869) );
  XNOR2_X1 U948 ( .A(KEYINPUT21), .B(n869), .ZN(n870) );
  NAND2_X1 U949 ( .A1(n870), .A2(G2072), .ZN(n871) );
  XOR2_X1 U950 ( .A(KEYINPUT85), .B(n871), .Z(G158) );
  XNOR2_X1 U951 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U952 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U953 ( .A1(G108), .A2(G120), .ZN(n872) );
  NOR2_X1 U954 ( .A1(G237), .A2(n872), .ZN(n873) );
  NAND2_X1 U955 ( .A1(G69), .A2(n873), .ZN(n884) );
  NAND2_X1 U956 ( .A1(n884), .A2(G567), .ZN(n878) );
  NOR2_X1 U957 ( .A1(G220), .A2(G219), .ZN(n874) );
  XOR2_X1 U958 ( .A(KEYINPUT22), .B(n874), .Z(n875) );
  NOR2_X1 U959 ( .A1(G218), .A2(n875), .ZN(n876) );
  NAND2_X1 U960 ( .A1(G96), .A2(n876), .ZN(n885) );
  NAND2_X1 U961 ( .A1(n885), .A2(G2106), .ZN(n877) );
  NAND2_X1 U962 ( .A1(n878), .A2(n877), .ZN(n886) );
  NAND2_X1 U963 ( .A1(G661), .A2(G483), .ZN(n879) );
  NOR2_X1 U964 ( .A1(n886), .A2(n879), .ZN(n883) );
  NAND2_X1 U965 ( .A1(n883), .A2(G36), .ZN(G176) );
  NAND2_X1 U966 ( .A1(G2106), .A2(n880), .ZN(G217) );
  AND2_X1 U967 ( .A1(G15), .A2(G2), .ZN(n881) );
  NAND2_X1 U968 ( .A1(G661), .A2(n881), .ZN(G259) );
  NAND2_X1 U969 ( .A1(G3), .A2(G1), .ZN(n882) );
  NAND2_X1 U970 ( .A1(n883), .A2(n882), .ZN(G188) );
  INV_X1 U972 ( .A(G120), .ZN(G236) );
  INV_X1 U973 ( .A(G108), .ZN(G238) );
  INV_X1 U974 ( .A(G96), .ZN(G221) );
  INV_X1 U975 ( .A(G69), .ZN(G235) );
  NOR2_X1 U976 ( .A1(n885), .A2(n884), .ZN(G325) );
  INV_X1 U977 ( .A(G325), .ZN(G261) );
  INV_X1 U978 ( .A(n886), .ZN(G319) );
  XOR2_X1 U979 ( .A(G2100), .B(G2096), .Z(n888) );
  XNOR2_X1 U980 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U982 ( .A(G2678), .B(G2090), .Z(n890) );
  XNOR2_X1 U983 ( .A(G2067), .B(G2072), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U985 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U986 ( .A(G2078), .B(G2084), .ZN(n893) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(G227) );
  XOR2_X1 U988 ( .A(G1976), .B(G1971), .Z(n896) );
  XNOR2_X1 U989 ( .A(G1986), .B(G1956), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U991 ( .A(G1961), .B(G1966), .Z(n898) );
  XNOR2_X1 U992 ( .A(G1996), .B(G1991), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U995 ( .A(KEYINPUT107), .B(G2474), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n904) );
  XOR2_X1 U997 ( .A(G1981), .B(KEYINPUT41), .Z(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(G229) );
  NAND2_X1 U999 ( .A1(G112), .A2(n936), .ZN(n906) );
  NAND2_X1 U1000 ( .A1(G100), .A2(n623), .ZN(n905) );
  NAND2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(n937), .A2(G124), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n907), .B(KEYINPUT44), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n519), .A2(G136), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(G162) );
  XNOR2_X1 U1007 ( .A(G164), .B(n912), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n913), .B(n986), .ZN(n918) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1010 ( .A(n916), .B(G160), .Z(n917) );
  XOR2_X1 U1011 ( .A(n918), .B(n917), .Z(n923) );
  XOR2_X1 U1012 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n920) );
  XNOR2_X1 U1013 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(KEYINPUT110), .B(n921), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(n923), .B(n922), .ZN(n933) );
  NAND2_X1 U1017 ( .A1(n519), .A2(G142), .ZN(n925) );
  NAND2_X1 U1018 ( .A1(G106), .A2(n623), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(n926), .B(KEYINPUT45), .ZN(n928) );
  NAND2_X1 U1021 ( .A1(G130), .A2(n937), .ZN(n927) );
  NAND2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n931) );
  NAND2_X1 U1023 ( .A1(n936), .A2(G118), .ZN(n929) );
  XOR2_X1 U1024 ( .A(KEYINPUT108), .B(n929), .Z(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1026 ( .A(n933), .B(n932), .Z(n945) );
  NAND2_X1 U1027 ( .A1(n519), .A2(G139), .ZN(n935) );
  NAND2_X1 U1028 ( .A1(G103), .A2(n623), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n943) );
  NAND2_X1 U1030 ( .A1(G115), .A2(n936), .ZN(n939) );
  NAND2_X1 U1031 ( .A1(G127), .A2(n937), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT109), .B(n940), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT47), .B(n941), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n976) );
  XNOR2_X1 U1036 ( .A(n976), .B(G162), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(n945), .B(n944), .ZN(n946) );
  NOR2_X1 U1038 ( .A1(G37), .A2(n946), .ZN(G395) );
  XNOR2_X1 U1039 ( .A(n1045), .B(G286), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(n689), .B(G171), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(n948), .B(n947), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(n950), .B(n949), .ZN(n951) );
  NOR2_X1 U1043 ( .A1(G37), .A2(n951), .ZN(G397) );
  XOR2_X1 U1044 ( .A(G2438), .B(G2454), .Z(n953) );
  XNOR2_X1 U1045 ( .A(G2451), .B(G2430), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(n953), .B(n952), .ZN(n954) );
  XOR2_X1 U1047 ( .A(n954), .B(G2435), .Z(n956) );
  XNOR2_X1 U1048 ( .A(G1348), .B(G1341), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(n956), .B(n955), .ZN(n960) );
  XOR2_X1 U1050 ( .A(G2427), .B(G2446), .Z(n958) );
  XNOR2_X1 U1051 ( .A(G2443), .B(KEYINPUT106), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(n958), .B(n957), .ZN(n959) );
  XOR2_X1 U1053 ( .A(n960), .B(n959), .Z(n961) );
  NAND2_X1 U1054 ( .A1(G14), .A2(n961), .ZN(n968) );
  NAND2_X1 U1055 ( .A1(G319), .A2(n968), .ZN(n965) );
  NOR2_X1 U1056 ( .A1(G227), .A2(G229), .ZN(n962) );
  XOR2_X1 U1057 ( .A(KEYINPUT113), .B(n962), .Z(n963) );
  XNOR2_X1 U1058 ( .A(n963), .B(KEYINPUT49), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(G395), .A2(G397), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(G225) );
  INV_X1 U1062 ( .A(G225), .ZN(G308) );
  INV_X1 U1063 ( .A(n968), .ZN(G401) );
  XOR2_X1 U1064 ( .A(G2090), .B(G162), .Z(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(n971), .B(KEYINPUT51), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n984) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n817), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(G2072), .B(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G164), .B(G2078), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT115), .B(n979), .Z(n980) );
  XNOR2_X1 U1073 ( .A(KEYINPUT50), .B(n980), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n991) );
  XNOR2_X1 U1076 ( .A(G160), .B(G2084), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n988) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1079 ( .A(KEYINPUT114), .B(n989), .Z(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1081 ( .A(KEYINPUT52), .B(n992), .Z(n993) );
  NOR2_X1 U1082 ( .A1(KEYINPUT55), .A2(n993), .ZN(n994) );
  XOR2_X1 U1083 ( .A(KEYINPUT116), .B(n994), .Z(n995) );
  NAND2_X1 U1084 ( .A1(G29), .A2(n995), .ZN(n1074) );
  XOR2_X1 U1085 ( .A(G1961), .B(KEYINPUT124), .Z(n996) );
  XNOR2_X1 U1086 ( .A(G5), .B(n996), .ZN(n1017) );
  XOR2_X1 U1087 ( .A(G1966), .B(G21), .Z(n1005) );
  XOR2_X1 U1088 ( .A(G1971), .B(G22), .Z(n999) );
  XOR2_X1 U1089 ( .A(G24), .B(KEYINPUT126), .Z(n997) );
  XNOR2_X1 U1090 ( .A(n997), .B(G1986), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(KEYINPUT125), .B(G1976), .Z(n1000) );
  XNOR2_X1 U1093 ( .A(G23), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(KEYINPUT58), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1015) );
  XOR2_X1 U1097 ( .A(G1348), .B(G4), .Z(n1006) );
  XNOR2_X1 U1098 ( .A(KEYINPUT59), .B(n1006), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(G20), .B(G1956), .ZN(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(G1341), .B(G19), .ZN(n1010) );
  XNOR2_X1 U1102 ( .A(G1981), .B(G6), .ZN(n1009) );
  NOR2_X1 U1103 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(n1018), .B(KEYINPUT127), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(n1019), .B(KEYINPUT61), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(G16), .B(KEYINPUT123), .ZN(n1020) );
  NAND2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1112 ( .A1(G11), .A2(n1022), .ZN(n1072) );
  XOR2_X1 U1113 ( .A(G29), .B(KEYINPUT118), .Z(n1042) );
  XOR2_X1 U1114 ( .A(G1991), .B(G25), .Z(n1023) );
  NAND2_X1 U1115 ( .A1(n1023), .A2(G28), .ZN(n1032) );
  XNOR2_X1 U1116 ( .A(G1996), .B(G32), .ZN(n1025) );
  XNOR2_X1 U1117 ( .A(G33), .B(G2072), .ZN(n1024) );
  NOR2_X1 U1118 ( .A1(n1025), .A2(n1024), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(G2067), .B(G26), .ZN(n1028) );
  XNOR2_X1 U1120 ( .A(G27), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1121 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1122 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1123 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1124 ( .A(KEYINPUT53), .B(n1033), .Z(n1037) );
  XNOR2_X1 U1125 ( .A(KEYINPUT54), .B(G34), .ZN(n1034) );
  XNOR2_X1 U1126 ( .A(n1034), .B(KEYINPUT117), .ZN(n1035) );
  XNOR2_X1 U1127 ( .A(G2084), .B(n1035), .ZN(n1036) );
  NAND2_X1 U1128 ( .A1(n1037), .A2(n1036), .ZN(n1039) );
  XNOR2_X1 U1129 ( .A(G35), .B(G2090), .ZN(n1038) );
  NOR2_X1 U1130 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1131 ( .A(n1040), .B(KEYINPUT55), .ZN(n1041) );
  NAND2_X1 U1132 ( .A1(n1042), .A2(n1041), .ZN(n1070) );
  XNOR2_X1 U1133 ( .A(KEYINPUT56), .B(G16), .ZN(n1068) );
  XNOR2_X1 U1134 ( .A(G171), .B(G1961), .ZN(n1044) );
  NAND2_X1 U1135 ( .A1(G1971), .A2(G303), .ZN(n1043) );
  NAND2_X1 U1136 ( .A1(n1044), .A2(n1043), .ZN(n1047) );
  XNOR2_X1 U1137 ( .A(G1341), .B(n1045), .ZN(n1046) );
  NOR2_X1 U1138 ( .A1(n1047), .A2(n1046), .ZN(n1049) );
  NAND2_X1 U1139 ( .A1(n1049), .A2(n1048), .ZN(n1056) );
  XNOR2_X1 U1140 ( .A(G1966), .B(G168), .ZN(n1051) );
  NAND2_X1 U1141 ( .A1(n1051), .A2(n1050), .ZN(n1052) );
  XNOR2_X1 U1142 ( .A(n1052), .B(KEYINPUT57), .ZN(n1054) );
  XNOR2_X1 U1143 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n1053) );
  XNOR2_X1 U1144 ( .A(n1054), .B(n1053), .ZN(n1055) );
  NOR2_X1 U1145 ( .A1(n1056), .A2(n1055), .ZN(n1066) );
  XNOR2_X1 U1146 ( .A(G1956), .B(KEYINPUT122), .ZN(n1057) );
  XNOR2_X1 U1147 ( .A(n1057), .B(G299), .ZN(n1058) );
  NOR2_X1 U1148 ( .A1(n1059), .A2(n1058), .ZN(n1060) );
  NAND2_X1 U1149 ( .A1(n1061), .A2(n1060), .ZN(n1064) );
  XOR2_X1 U1150 ( .A(G1348), .B(n689), .Z(n1062) );
  XNOR2_X1 U1151 ( .A(KEYINPUT121), .B(n1062), .ZN(n1063) );
  NOR2_X1 U1152 ( .A1(n1064), .A2(n1063), .ZN(n1065) );
  NAND2_X1 U1153 ( .A1(n1066), .A2(n1065), .ZN(n1067) );
  NAND2_X1 U1154 ( .A1(n1068), .A2(n1067), .ZN(n1069) );
  NAND2_X1 U1155 ( .A1(n1070), .A2(n1069), .ZN(n1071) );
  NOR2_X1 U1156 ( .A1(n1072), .A2(n1071), .ZN(n1073) );
  NAND2_X1 U1157 ( .A1(n1074), .A2(n1073), .ZN(n1075) );
  XOR2_X1 U1158 ( .A(KEYINPUT62), .B(n1075), .Z(G311) );
  INV_X1 U1159 ( .A(G311), .ZN(G150) );
endmodule

