//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n206), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT0), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n217), .A2(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n223), .B1(new_n222), .B2(new_n221), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n214), .A2(new_n224), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n229), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  XNOR2_X1  g0041(.A(KEYINPUT3), .B(G33), .ZN(new_n242));
  INV_X1    g0042(.A(G1698), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n242), .A2(G222), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n242), .A2(G223), .A3(G1698), .ZN(new_n245));
  OAI211_X1 g0045(.A(new_n244), .B(new_n245), .C1(new_n202), .C2(new_n242), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n247), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n246), .A2(KEYINPUT67), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(KEYINPUT67), .B2(new_n246), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n254), .B(G274), .C1(G41), .C2(G45), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n248), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n258), .B2(G226), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G190), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(G200), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n216), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT65), .A2(G20), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT65), .A2(G20), .ZN(new_n267));
  OAI21_X1  g0067(.A(G33), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT8), .A2(G58), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT8), .A2(G58), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n268), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G20), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n277), .A2(new_n279), .B1(new_n201), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n265), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n265), .B1(new_n254), .B2(G20), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(G50), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT9), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n262), .A2(new_n263), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT10), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n264), .A2(new_n216), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n215), .A2(G33), .A3(G77), .ZN(new_n292));
  INV_X1    g0092(.A(G68), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n278), .A2(G50), .B1(G20), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT11), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(KEYINPUT11), .ZN(new_n297));
  OR3_X1    g0097(.A1(new_n283), .A2(KEYINPUT12), .A3(G68), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT12), .B1(new_n283), .B2(G68), .ZN(new_n299));
  AOI22_X1  g0099(.A1(G68), .A2(new_n285), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT3), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G33), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n303), .A2(new_n305), .A3(G232), .A4(G1698), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n303), .A2(new_n305), .A3(G226), .A4(new_n243), .ZN(new_n307));
  INV_X1    g0107(.A(G97), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n306), .B(new_n307), .C1(new_n302), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n250), .A2(new_n251), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n256), .B1(new_n258), .B2(G238), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT13), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(G179), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n314), .B2(new_n316), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT14), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n316), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n315), .B1(new_n311), .B2(new_n312), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n320), .B(G169), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n301), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n322), .A2(new_n323), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n301), .B1(new_n327), .B2(G190), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n327), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n287), .B1(new_n261), .B2(G169), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n260), .A2(G179), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n290), .A2(new_n326), .A3(new_n330), .A4(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT7), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n304), .A2(G33), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n302), .A2(KEYINPUT3), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n336), .B(new_n280), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(KEYINPUT65), .A2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(KEYINPUT65), .A2(G20), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n303), .A2(new_n305), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n339), .B(G68), .C1(new_n342), .C2(new_n336), .ZN(new_n343));
  XNOR2_X1  g0143(.A(G58), .B(G68), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(G20), .B1(new_n303), .B2(new_n305), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n350), .B2(new_n336), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n303), .A2(new_n305), .ZN(new_n352));
  AND3_X1   g0152(.A1(new_n352), .A2(new_n215), .A3(new_n336), .ZN(new_n353));
  OAI211_X1 g0153(.A(KEYINPUT16), .B(new_n345), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n349), .A2(new_n265), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n248), .A2(G232), .A3(new_n257), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n255), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n303), .A2(new_n305), .A3(G226), .A4(G1698), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n303), .A2(new_n305), .A3(G223), .A4(new_n243), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI211_X1 g0162(.A(new_n356), .B(new_n358), .C1(new_n310), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n310), .ZN(new_n364));
  INV_X1    g0164(.A(new_n358), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n329), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n272), .A2(new_n275), .ZN(new_n368));
  INV_X1    g0168(.A(new_n285), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n272), .A2(new_n275), .A3(new_n283), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n355), .A2(new_n367), .A3(KEYINPUT74), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n370), .A2(new_n371), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n354), .A2(new_n265), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n349), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n378), .A2(KEYINPUT74), .A3(KEYINPUT17), .A4(new_n367), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n354), .A2(new_n265), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n347), .B1(new_n343), .B2(new_n345), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n372), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n358), .B1(new_n362), .B2(new_n310), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G179), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n318), .B2(new_n384), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n383), .A2(KEYINPUT18), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT18), .B1(new_n383), .B2(new_n386), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n380), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n340), .A2(G77), .A3(new_n341), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n269), .A2(new_n278), .A3(new_n270), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT15), .B(G87), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n391), .B(new_n392), .C1(new_n268), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n265), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n283), .A2(G77), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n285), .B2(G77), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT70), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(new_n397), .A3(KEYINPUT70), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n303), .A2(new_n305), .A3(G238), .A4(G1698), .ZN(new_n403));
  INV_X1    g0203(.A(G107), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(new_n242), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n242), .A2(G232), .A3(new_n243), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n310), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n256), .B1(new_n258), .B2(G244), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n402), .B1(G200), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n356), .B2(new_n409), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n400), .A2(new_n401), .B1(new_n409), .B2(new_n318), .ZN(new_n412));
  INV_X1    g0212(.A(G179), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n407), .A2(KEYINPUT71), .A3(new_n413), .A4(new_n408), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT71), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n409), .B2(G179), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n412), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT72), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n335), .A2(new_n390), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n303), .A2(new_n305), .A3(G257), .A4(new_n243), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT78), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n242), .A2(KEYINPUT78), .A3(G257), .A4(new_n243), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n242), .A2(G264), .A3(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n352), .A2(G303), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G45), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G1), .ZN(new_n430));
  INV_X1    g0230(.A(G41), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT5), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT5), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G41), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n435), .A2(new_n248), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n428), .A2(new_n310), .B1(G270), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n430), .A2(G274), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(new_n434), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G116), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n264), .A2(new_n216), .B1(G20), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(KEYINPUT75), .A2(G97), .ZN(new_n445));
  NOR2_X1   g0245(.A1(KEYINPUT75), .A2(G97), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n445), .A2(new_n446), .A3(G33), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n266), .B2(new_n267), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n444), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT20), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(KEYINPUT20), .B(new_n444), .C1(new_n447), .C2(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n283), .A2(G116), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n254), .A2(G33), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n283), .A2(new_n457), .A3(new_n216), .A4(new_n264), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(new_n443), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT79), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  AOI211_X1 g0262(.A(new_n462), .B(new_n459), .C1(new_n452), .C2(new_n453), .ZN(new_n463));
  OAI211_X1 g0263(.A(G169), .B(new_n442), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT21), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n453), .ZN(new_n467));
  OR2_X1    g0267(.A1(KEYINPUT75), .A2(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT75), .A2(G97), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n302), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(new_n215), .A3(new_n448), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT20), .B1(new_n471), .B2(new_n444), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n460), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n462), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n454), .A2(KEYINPUT79), .A3(new_n460), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n413), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n442), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n475), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n479), .A2(KEYINPUT21), .A3(G169), .A4(new_n442), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n442), .A2(G200), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n437), .A2(G190), .A3(new_n441), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n481), .A2(new_n474), .A3(new_n475), .A4(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n466), .A2(new_n478), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n303), .A2(new_n305), .A3(G250), .A4(new_n243), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n303), .A2(new_n305), .A3(G257), .A4(G1698), .ZN(new_n486));
  XOR2_X1   g0286(.A(KEYINPUT82), .B(G294), .Z(new_n487));
  OAI211_X1 g0287(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(new_n302), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n440), .B1(new_n488), .B2(new_n310), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n435), .A2(G264), .A3(new_n248), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n318), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n310), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT83), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n435), .A2(KEYINPUT83), .A3(G264), .A4(new_n248), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n493), .A2(new_n441), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n413), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n458), .ZN(new_n500));
  INV_X1    g0300(.A(new_n283), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(KEYINPUT25), .A3(new_n404), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT25), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n283), .B2(G107), .ZN(new_n504));
  AOI22_X1  g0304(.A1(G107), .A2(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(KEYINPUT23), .A2(G107), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n340), .A2(new_n341), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT23), .B1(new_n280), .B2(G107), .ZN(new_n508));
  AND2_X1   g0308(.A1(G33), .A2(G116), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT80), .B1(new_n509), .B2(new_n280), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G116), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT80), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n511), .A2(new_n512), .A3(G20), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n507), .B(new_n508), .C1(new_n510), .C2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n215), .A2(new_n242), .A3(G87), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT22), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT22), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n215), .A2(new_n242), .A3(new_n517), .A4(G87), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n265), .B1(new_n519), .B2(KEYINPUT24), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT24), .ZN(new_n521));
  AOI211_X1 g0321(.A(new_n521), .B(new_n514), .C1(new_n516), .C2(new_n518), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n505), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(KEYINPUT81), .B(new_n505), .C1(new_n520), .C2(new_n522), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n499), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n279), .A2(new_n202), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  AND2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n468), .A2(new_n469), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n404), .A2(KEYINPUT6), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n266), .A2(new_n267), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n528), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n339), .B(G107), .C1(new_n342), .C2(new_n336), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n265), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n283), .A2(G97), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n500), .B2(G97), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(KEYINPUT77), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT77), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n291), .B1(new_n537), .B2(new_n538), .ZN(new_n545));
  INV_X1    g0345(.A(new_n542), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n303), .A2(new_n305), .A3(G244), .A4(new_n243), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT4), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n242), .A2(KEYINPUT4), .A3(G244), .A4(new_n243), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n242), .A2(G250), .A3(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n448), .A4(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n554), .A2(new_n310), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n435), .A2(G257), .A3(new_n248), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT76), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n435), .A2(KEYINPUT76), .A3(G257), .A4(new_n248), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n441), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(G169), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n554), .A2(new_n310), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(G179), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n548), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n248), .ZN(new_n567));
  OAI21_X1  g0367(.A(G250), .B1(new_n429), .B2(G1), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n438), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n303), .A2(new_n305), .A3(G244), .A4(G1698), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n303), .A2(new_n305), .A3(G238), .A4(new_n243), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n511), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n572), .B2(new_n310), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(G169), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n413), .B2(new_n573), .ZN(new_n575));
  INV_X1    g0375(.A(new_n393), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(new_n283), .ZN(new_n577));
  INV_X1    g0377(.A(G87), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n578), .B(new_n404), .C1(new_n445), .C2(new_n446), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n302), .A2(new_n308), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n579), .B(KEYINPUT19), .C1(new_n536), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n215), .A2(new_n242), .A3(G68), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n268), .B2(new_n533), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n577), .B1(new_n585), .B2(new_n265), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n393), .B2(new_n458), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n573), .A2(new_n329), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n356), .B(new_n569), .C1(new_n572), .C2(new_n310), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n458), .A2(new_n578), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n577), .B(new_n591), .C1(new_n585), .C2(new_n265), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n575), .A2(new_n587), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n497), .A2(new_n329), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n489), .A2(new_n356), .A3(new_n490), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n516), .A2(new_n518), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n521), .B1(new_n597), .B2(new_n514), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n519), .A2(KEYINPUT24), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n265), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n600), .A3(new_n505), .ZN(new_n601));
  OAI21_X1  g0401(.A(G200), .B1(new_n555), .B2(new_n560), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n545), .A2(new_n546), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n562), .A2(G190), .A3(new_n563), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n566), .A2(new_n593), .A3(new_n601), .A4(new_n605), .ZN(new_n606));
  NOR4_X1   g0406(.A1(new_n421), .A2(new_n484), .A3(new_n527), .A4(new_n606), .ZN(G372));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n387), .B2(new_n388), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n383), .A2(new_n386), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n383), .A2(KEYINPUT18), .A3(new_n386), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(KEYINPUT84), .A3(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n417), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT14), .B1(new_n327), .B2(new_n318), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n324), .A3(new_n317), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n616), .A2(new_n330), .B1(new_n618), .B2(new_n301), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n615), .B1(new_n619), .B2(new_n380), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n333), .B1(new_n620), .B2(new_n290), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n575), .A2(new_n587), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n590), .A2(new_n592), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT26), .B1(new_n624), .B2(new_n566), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  INV_X1    g0426(.A(new_n603), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n593), .A2(new_n626), .A3(new_n565), .A4(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n622), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n606), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n465), .A2(new_n464), .B1(new_n476), .B2(new_n477), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n480), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n492), .A2(new_n498), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n523), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n631), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n621), .B1(new_n421), .B2(new_n639), .ZN(G369));
  INV_X1    g0440(.A(new_n484), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n215), .A2(G13), .ZN(new_n642));
  OR3_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .A3(G1), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT27), .B1(new_n642), .B2(G1), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n479), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n466), .A2(new_n478), .A3(new_n480), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(new_n648), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT81), .B1(new_n600), .B2(new_n505), .ZN(new_n653));
  INV_X1    g0453(.A(new_n526), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n634), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n647), .B1(new_n653), .B2(new_n654), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(new_n601), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT85), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT85), .A4(new_n601), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n527), .A2(new_n647), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n652), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n650), .A2(new_n647), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n659), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n647), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n636), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n663), .A2(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n220), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G1), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n579), .A2(G116), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n673), .A2(new_n674), .B1(new_n218), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  INV_X1    g0476(.A(G330), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n555), .A2(new_n413), .A3(new_n560), .ZN(new_n678));
  INV_X1    g0478(.A(new_n573), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n497), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n678), .A2(new_n680), .A3(KEYINPUT30), .A4(new_n437), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n495), .A2(new_n496), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n437), .A2(new_n489), .A3(new_n683), .A4(new_n573), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n682), .B1(new_n684), .B2(new_n564), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n562), .A2(new_n563), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n573), .A2(G179), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n442), .A2(new_n686), .A3(new_n497), .A4(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n681), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT31), .B1(new_n689), .B2(new_n647), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n641), .A2(new_n631), .A3(new_n655), .A4(new_n666), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n677), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n655), .A2(new_n480), .A3(new_n632), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT87), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n547), .A2(new_n543), .B1(new_n561), .B2(new_n564), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n566), .A2(KEYINPUT87), .A3(new_n605), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n702), .A3(new_n601), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n626), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n624), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n622), .B(KEYINPUT86), .Z(new_n706));
  NAND2_X1  g0506(.A1(new_n565), .A2(new_n627), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT26), .B1(new_n624), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT29), .B(new_n666), .C1(new_n705), .C2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT88), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n647), .B1(new_n630), .B2(new_n637), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n601), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n700), .B2(new_n701), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n716), .A2(new_n696), .B1(new_n626), .B2(new_n698), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n708), .B(new_n706), .C1(new_n717), .C2(new_n624), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n711), .A3(KEYINPUT29), .A4(new_n666), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n695), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n676), .B1(new_n720), .B2(G1), .ZN(G364));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n651), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n216), .B1(G20), .B2(new_n318), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n670), .A2(new_n352), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT89), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G355), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G116), .B2(new_n220), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n670), .A2(new_n242), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G45), .B2(new_n218), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n240), .B2(G45), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n728), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(G1), .B1(new_n642), .B2(new_n429), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n671), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OR3_X1    g0539(.A1(new_n215), .A2(KEYINPUT92), .A3(G190), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT92), .B1(new_n215), .B2(G190), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n329), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n404), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n356), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n413), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n536), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G97), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n742), .A2(G20), .A3(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n352), .B1(new_n750), .B2(G87), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n215), .A2(new_n413), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n356), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n329), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n748), .B(new_n751), .C1(new_n755), .C2(new_n293), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT91), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n757), .A2(new_n758), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n744), .B(new_n756), .C1(G50), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n740), .A2(new_n741), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT93), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n413), .A2(new_n329), .ZN(new_n767));
  OR3_X1    g0567(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT32), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OR3_X1    g0572(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n771), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n752), .A2(new_n356), .A3(new_n329), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n752), .A2(new_n745), .ZN(new_n775));
  INV_X1    g0575(.A(G58), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n774), .A2(new_n202), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT90), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n764), .A2(new_n772), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n770), .A2(KEYINPUT94), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n770), .A2(KEYINPUT94), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(G329), .ZN(new_n784));
  INV_X1    g0584(.A(new_n743), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n763), .A2(G326), .B1(new_n785), .B2(G283), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n775), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G303), .ZN(new_n789));
  INV_X1    g0589(.A(new_n747), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n352), .B1(new_n789), .B2(new_n749), .C1(new_n790), .C2(new_n487), .ZN(new_n791));
  INV_X1    g0591(.A(new_n774), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n788), .B(new_n791), .C1(G311), .C2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT33), .B(G317), .Z(new_n794));
  OAI211_X1 g0594(.A(new_n786), .B(new_n793), .C1(new_n755), .C2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n779), .B1(new_n784), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n739), .B1(new_n796), .B2(new_n727), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n726), .A2(KEYINPUT95), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT95), .B1(new_n726), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n651), .A2(G330), .ZN(new_n800));
  INV_X1    g0600(.A(new_n738), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n652), .A2(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(new_n802), .ZN(G396));
  OAI21_X1  g0603(.A(KEYINPUT98), .B1(new_n417), .B2(new_n666), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n409), .A2(new_n318), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n402), .A2(new_n416), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT98), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n806), .A2(new_n807), .A3(new_n414), .A4(new_n647), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n402), .A2(new_n647), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n411), .A2(new_n417), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n712), .B(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n695), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n815), .A2(new_n801), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n727), .A2(new_n722), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n801), .B1(new_n202), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n775), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n792), .A2(G159), .B1(new_n820), .B2(G143), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n277), .B2(new_n755), .C1(new_n762), .C2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT34), .Z(new_n824));
  OAI21_X1  g0624(.A(new_n242), .B1(new_n790), .B2(new_n776), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n785), .A2(G68), .ZN(new_n826));
  INV_X1    g0626(.A(G50), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n827), .B2(new_n749), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n825), .B1(new_n828), .B2(KEYINPUT97), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(KEYINPUT97), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n783), .A2(G132), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n783), .A2(G311), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n352), .B1(new_n404), .B2(new_n749), .C1(new_n755), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G294), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n748), .B1(new_n775), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n785), .A2(G87), .B1(new_n837), .B2(KEYINPUT96), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(KEYINPUT96), .B2(new_n837), .C1(new_n789), .C2(new_n762), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n835), .B(new_n839), .C1(G116), .C2(new_n792), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n727), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n819), .B1(new_n723), .B2(new_n812), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n817), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  OAI21_X1  g0645(.A(G77), .B1(new_n776), .B2(new_n293), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n846), .A2(new_n218), .B1(G50), .B2(new_n293), .ZN(new_n847));
  INV_X1    g0647(.A(G13), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(G1), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(G116), .B(new_n217), .C1(new_n535), .C2(KEYINPUT35), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(KEYINPUT35), .B2(new_n535), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT99), .Z(new_n852));
  INV_X1    g0652(.A(KEYINPUT36), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  NOR4_X1   g0655(.A1(new_n484), .A2(new_n606), .A3(new_n527), .A4(new_n647), .ZN(new_n856));
  INV_X1    g0656(.A(new_n692), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n690), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT40), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n345), .B1(new_n351), .B2(new_n353), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n381), .B1(new_n348), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n376), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n645), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n380), .B2(new_n389), .ZN(new_n864));
  INV_X1    g0664(.A(new_n645), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n383), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n355), .A2(new_n367), .A3(new_n372), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n610), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n378), .B2(new_n367), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n861), .A2(new_n376), .B1(new_n386), .B2(new_n865), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n868), .A2(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n869), .B1(new_n866), .B2(KEYINPUT101), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n868), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n874), .A2(new_n867), .A3(new_n610), .A4(new_n866), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n380), .A2(KEYINPUT102), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT102), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n375), .A2(new_n379), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n879), .A2(new_n609), .A3(new_n614), .A4(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n866), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n873), .B1(new_n884), .B2(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n301), .A2(new_n647), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n326), .A2(new_n330), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n618), .A2(new_n301), .A3(new_n647), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n887), .A2(new_n888), .B1(new_n809), .B2(new_n811), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n856), .B2(new_n858), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n859), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n873), .A2(KEYINPUT100), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n864), .B2(new_n872), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n889), .B(new_n859), .C1(new_n856), .C2(new_n858), .ZN(new_n896));
  AOI211_X1 g0696(.A(KEYINPUT100), .B(KEYINPUT38), .C1(new_n864), .C2(new_n872), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n420), .B1(new_n856), .B2(new_n858), .C1(new_n892), .C2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n873), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n881), .A2(new_n609), .A3(new_n614), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n880), .B1(new_n375), .B2(new_n379), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n883), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n878), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT40), .B1(new_n907), .B2(new_n890), .ZN(new_n908));
  INV_X1    g0708(.A(new_n897), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n864), .A2(new_n872), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n906), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(KEYINPUT100), .A3(new_n873), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n891), .A2(new_n859), .A3(new_n909), .A4(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n677), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n420), .A2(new_n695), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n899), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n714), .A2(new_n420), .A3(new_n719), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n918), .A2(new_n621), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT39), .B1(new_n895), .B2(new_n897), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n326), .A2(new_n647), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n903), .B2(new_n904), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(new_n924), .B2(new_n900), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n615), .A2(new_n865), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n895), .A2(new_n897), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n887), .A2(new_n888), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n606), .B1(new_n650), .B2(new_n635), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n666), .B(new_n812), .C1(new_n931), .C2(new_n629), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n417), .A2(new_n647), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n930), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n927), .B1(new_n928), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n926), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT103), .Z(new_n938));
  NAND2_X1  g0738(.A1(new_n920), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n642), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n939), .B1(new_n254), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n920), .A2(new_n938), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n855), .B1(new_n941), .B2(new_n942), .ZN(G367));
  OR3_X1    g0743(.A1(new_n622), .A2(new_n592), .A3(new_n666), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n593), .B1(new_n592), .B2(new_n666), .ZN(new_n945));
  XNOR2_X1  g0745(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n947), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n659), .A2(new_n660), .A3(new_n664), .A4(new_n702), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n702), .B1(new_n603), .B2(new_n666), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n565), .A2(new_n627), .A3(new_n647), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n698), .B1(new_n956), .B2(new_n527), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n952), .B(new_n953), .C1(new_n647), .C2(new_n957), .ZN(new_n958));
  MUX2_X1   g0758(.A(new_n947), .B(new_n950), .S(new_n958), .Z(new_n959));
  NAND2_X1  g0759(.A1(new_n663), .A2(new_n956), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n737), .B(KEYINPUT107), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n665), .A2(new_n667), .A3(new_n956), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  INV_X1    g0767(.A(new_n956), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n668), .A2(KEYINPUT44), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT44), .B1(new_n668), .B2(new_n968), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n966), .A2(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n661), .A2(new_n662), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n665), .B1(new_n972), .B2(new_n664), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n663), .B1(new_n973), .B2(new_n652), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n720), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT105), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT105), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n971), .A2(new_n720), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n720), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n671), .B(KEYINPUT41), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT106), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n963), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n981), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n979), .B2(new_n720), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT106), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n962), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(G311), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n762), .A2(new_n989), .B1(new_n533), .B2(new_n743), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n749), .A2(new_n443), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(KEYINPUT46), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G107), .B2(new_n747), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n242), .B1(new_n991), .B2(KEYINPUT46), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(new_n789), .C2(new_n775), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n755), .A2(new_n487), .B1(new_n834), .B2(new_n774), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n990), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(G317), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n998), .B2(new_n770), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n743), .A2(new_n202), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n242), .B1(new_n776), .B2(new_n749), .C1(new_n755), .C2(new_n771), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G50), .C2(new_n792), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n822), .B2(new_n770), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n820), .A2(G150), .B1(G68), .B2(new_n747), .ZN(new_n1004));
  INV_X1    g0804(.A(G143), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n762), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT109), .Z(new_n1007));
  OAI21_X1  g0807(.A(new_n999), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT47), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n842), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n1009), .B2(new_n1008), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n944), .A2(new_n945), .A3(new_n724), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n233), .A2(new_n733), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n728), .C1(new_n220), .C2(new_n393), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT108), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1016), .A2(new_n1017), .A3(new_n801), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1011), .A2(new_n1012), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n988), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(G387));
  AOI21_X1  g0822(.A(new_n672), .B1(new_n720), .B2(new_n974), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n720), .B2(new_n974), .ZN(new_n1024));
  INV_X1    g0824(.A(G326), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n352), .B1(new_n443), .B2(new_n743), .C1(new_n770), .C2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n792), .A2(G303), .B1(new_n820), .B2(G317), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n989), .B2(new_n755), .C1(new_n762), .C2(new_n787), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n747), .A2(G283), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n487), .C2(new_n749), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1026), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n770), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(G150), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n242), .B1(new_n202), .B2(new_n749), .C1(new_n774), .C2(new_n293), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n368), .B2(new_n754), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n763), .A2(G159), .B1(new_n785), .B2(G97), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n747), .A2(new_n576), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n775), .B2(new_n827), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT113), .Z(new_n1042));
  NAND4_X1  g0842(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n842), .B1(new_n1034), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n972), .A2(new_n725), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n730), .A2(new_n674), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(G107), .B2(new_n220), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n674), .B(KEYINPUT110), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n273), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT50), .B1(new_n273), .B2(G50), .ZN(new_n1050));
  AOI21_X1  g0850(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n733), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT111), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1053), .A2(KEYINPUT111), .B1(new_n229), .B2(G45), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1047), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n728), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n738), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT112), .Z(new_n1059));
  NOR3_X1   g0859(.A1(new_n1044), .A2(new_n1045), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n974), .B2(new_n963), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1024), .A2(new_n1061), .ZN(G393));
  OR2_X1    g0862(.A1(new_n971), .A2(new_n663), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n971), .A2(new_n663), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n720), .A2(new_n974), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n979), .A2(new_n1067), .A3(new_n671), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1063), .A2(new_n963), .A3(new_n1064), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n733), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n728), .B1(new_n220), .B2(new_n533), .C1(new_n237), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT114), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n801), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n352), .B1(new_n749), .B2(new_n834), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n792), .A2(G294), .B1(G116), .B2(new_n747), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n789), .B2(new_n755), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n744), .B(new_n1075), .C1(new_n1078), .C2(KEYINPUT116), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(KEYINPUT116), .B2(new_n1078), .C1(new_n787), .C2(new_n770), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n762), .A2(new_n998), .B1(new_n989), .B2(new_n775), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT52), .Z(new_n1082));
  NOR2_X1   g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n790), .A2(new_n202), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n352), .B(new_n1086), .C1(G68), .C2(new_n750), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n827), .B2(new_n755), .C1(new_n273), .C2(new_n774), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G87), .B2(new_n785), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n762), .A2(new_n277), .B1(new_n771), .B2(new_n775), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1091));
  XNOR2_X1  g0891(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1089), .B(new_n1092), .C1(new_n1005), .C2(new_n770), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1085), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1074), .B1(new_n1095), .B2(new_n727), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n725), .B2(new_n956), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1069), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1068), .A2(new_n1098), .ZN(G390));
  NAND3_X1  g0899(.A1(new_n695), .A2(new_n812), .A3(new_n929), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n924), .A2(new_n900), .B1(new_n326), .B2(new_n647), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n666), .B(new_n812), .C1(new_n705), .C2(new_n709), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n934), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1102), .B1(new_n1104), .B2(new_n929), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n932), .A2(new_n934), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n922), .B1(new_n1106), .B2(new_n929), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n921), .B2(new_n925), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1101), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n905), .A2(new_n906), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT39), .B1(new_n1110), .B2(new_n873), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n923), .B1(new_n912), .B2(new_n909), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1111), .A2(new_n1112), .B1(new_n922), .B2(new_n935), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n930), .B1(new_n1103), .B2(new_n934), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n1100), .C1(new_n1114), .C2(new_n1102), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n918), .A2(new_n621), .A3(new_n915), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n932), .A2(new_n934), .ZN(new_n1118));
  OAI211_X1 g0918(.A(G330), .B(new_n812), .C1(new_n856), .C2(new_n858), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n930), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1118), .B1(new_n1120), .B2(new_n1100), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1104), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1120), .A2(new_n1100), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT118), .B1(new_n1116), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n672), .B1(new_n1116), .B2(new_n1125), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1109), .A2(new_n1115), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1103), .A2(new_n1120), .A3(new_n1100), .A4(new_n934), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1123), .B2(new_n1118), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n919), .A2(new_n915), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT118), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1126), .A2(new_n1127), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n818), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n738), .B1(new_n368), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n826), .B1(new_n782), .B2(new_n836), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1137), .A2(KEYINPUT120), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(KEYINPUT120), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n774), .A2(new_n533), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n242), .B(new_n1086), .C1(G87), .C2(new_n750), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1141), .B1(new_n404), .B2(new_n755), .C1(new_n443), .C2(new_n775), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(G283), .C2(new_n763), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  OR3_X1    g0944(.A1(new_n749), .A2(KEYINPUT53), .A3(new_n277), .ZN(new_n1145));
  OAI21_X1  g0945(.A(KEYINPUT53), .B1(new_n749), .B2(new_n277), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n242), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G132), .B2(new_n820), .ZN(new_n1148));
  INV_X1    g0948(.A(G128), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1148), .B1(new_n827), .B2(new_n743), .C1(new_n762), .C2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT54), .B(G143), .Z(new_n1151));
  NAND2_X1  g0951(.A1(new_n792), .A2(new_n1151), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n771), .B2(new_n790), .C1(new_n755), .C2(new_n822), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1150), .B1(KEYINPUT119), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(G125), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1154), .B1(KEYINPUT119), .B2(new_n1153), .C1(new_n782), .C2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT121), .B1(new_n1144), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(new_n842), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1144), .A2(KEYINPUT121), .A3(new_n1156), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1136), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1160), .B1(new_n723), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT122), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n963), .B2(new_n1116), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1134), .A2(new_n1164), .ZN(G378));
  NAND2_X1  g0965(.A1(new_n937), .A2(new_n914), .ZN(new_n1166));
  OAI21_X1  g0966(.A(G330), .B1(new_n892), .B2(new_n898), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n926), .A3(new_n936), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n290), .B1(new_n332), .B2(new_n331), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n645), .B1(new_n282), .B2(new_n286), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OR3_X1    g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1166), .A2(new_n1168), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT57), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1117), .B1(new_n1116), .B2(new_n1125), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n671), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n919), .B(new_n915), .C1(new_n1128), .C2(new_n1124), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT125), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1179), .A2(new_n1180), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1178), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1167), .B1(new_n926), .B2(new_n936), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n937), .A2(new_n914), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1166), .A2(new_n1168), .A3(new_n1178), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT125), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1184), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1183), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1185), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1190), .A2(KEYINPUT125), .A3(new_n1191), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n963), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1178), .A2(new_n722), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n738), .B1(G50), .B2(new_n1135), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n743), .A2(new_n776), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n431), .B(new_n352), .C1(new_n749), .C2(new_n202), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(new_n783), .C2(G283), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT124), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n820), .A2(G107), .B1(G68), .B2(new_n747), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n393), .B2(new_n774), .C1(new_n308), .C2(new_n755), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G116), .B2(new_n763), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT58), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1205), .A2(KEYINPUT58), .A3(new_n1208), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n775), .A2(new_n1149), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n750), .A2(new_n1151), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n790), .B2(new_n277), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(G137), .C2(new_n792), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n754), .A2(G132), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n1155), .C2(new_n762), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1035), .A2(G124), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n302), .A2(new_n431), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT123), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n785), .B2(G159), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1223), .B(new_n827), .C1(G41), .C2(new_n242), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1211), .A2(new_n1212), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1201), .B1(new_n1227), .B2(new_n727), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1200), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1199), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1195), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(G375));
  AOI21_X1  g1033(.A(new_n801), .B1(new_n293), .B2(new_n818), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n783), .A2(G128), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n754), .A2(new_n1151), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n792), .A2(G150), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n820), .A2(G137), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n242), .B1(new_n749), .B2(new_n771), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G50), .B2(new_n747), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1202), .B(new_n1241), .C1(G132), .C2(new_n763), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n783), .A2(G303), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n242), .B1(new_n750), .B2(G97), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n1040), .C1(new_n775), .C2(new_n834), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G107), .B2(new_n792), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n443), .B2(new_n755), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1000), .B(new_n1247), .C1(G294), .C2(new_n763), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1235), .A2(new_n1242), .B1(new_n1243), .B2(new_n1248), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1234), .B1(new_n723), .B2(new_n929), .C1(new_n1249), .C2(new_n842), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n963), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1250), .B1(new_n1124), .B2(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1125), .A2(new_n985), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G390), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1021), .A2(new_n1257), .A3(new_n1255), .A4(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(G378), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1232), .A2(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1259), .A2(new_n1261), .ZN(G407));
  NOR3_X1   g1062(.A1(new_n1195), .A2(new_n1231), .A3(G378), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n646), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G213), .B(new_n1264), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT126), .ZN(G409));
  OAI21_X1  g1066(.A(G378), .B1(new_n1195), .B2(new_n1231), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT60), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1254), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1117), .A2(KEYINPUT60), .A3(new_n1124), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n671), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT127), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n672), .B1(new_n1268), .B2(new_n1254), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1270), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1252), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n844), .B(new_n1252), .C1(new_n1272), .C2(new_n1275), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G213), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(G343), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1229), .B1(new_n1283), .B2(new_n963), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1134), .A2(new_n1284), .A3(new_n1164), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1182), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n981), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1282), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1267), .A2(new_n1280), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1282), .A2(G2897), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1273), .A2(new_n1274), .A3(new_n1270), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1274), .B1(new_n1273), .B2(new_n1270), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1277), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n844), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1276), .A2(G384), .A3(new_n1277), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1292), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1194), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n672), .B1(new_n1301), .B2(new_n1184), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1286), .B2(KEYINPUT57), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1229), .B1(new_n1198), .B2(new_n963), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1260), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1282), .ZN(new_n1306));
  AOI211_X1 g1106(.A(new_n985), .B(new_n1182), .C1(new_n1197), .C2(new_n1196), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1134), .A2(new_n1284), .A3(new_n1164), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1294), .B(new_n1300), .C1(new_n1305), .C2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1267), .A2(new_n1280), .A3(new_n1288), .A4(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1290), .A2(new_n1291), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1313));
  AND2_X1   g1113(.A1(G393), .A2(G396), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(G393), .A2(G396), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(G390), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1068), .B(new_n1098), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1319), .B1(new_n988), .B2(new_n1020), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n987), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1251), .B1(new_n986), .B2(KEYINPUT106), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n961), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1323), .A2(new_n1019), .A3(new_n1317), .A4(new_n1318), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1320), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1313), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1305), .A2(new_n1327), .A3(new_n1309), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1325), .B1(new_n1328), .B2(KEYINPUT63), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT63), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1289), .A2(new_n1330), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1329), .A2(new_n1291), .A3(new_n1310), .A4(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1326), .A2(new_n1332), .ZN(G405));
  NAND3_X1  g1133(.A1(new_n1261), .A2(new_n1327), .A3(new_n1267), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1280), .B1(new_n1263), .B2(new_n1305), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1325), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1336), .B(new_n1337), .ZN(G402));
endmodule


