//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G107), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n188), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n187), .A2(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G101), .B1(new_n192), .B2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n189), .B1(new_n191), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n193), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n188), .A4(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT0), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n209), .A2(KEYINPUT65), .A3(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT65), .B1(new_n209), .B2(G146), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n206), .B(new_n208), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n209), .A2(G146), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n207), .B2(G143), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n209), .A2(KEYINPUT65), .A3(G146), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(new_n206), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n206), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n209), .A2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n208), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n204), .A2(new_n205), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n227), .B(G101), .C1(new_n192), .C2(new_n196), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n203), .A2(new_n221), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT10), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n216), .A2(new_n217), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n231), .A2(new_n208), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n205), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n218), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT81), .B1(new_n187), .B2(G107), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n188), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n191), .A2(KEYINPUT81), .ZN(new_n239));
  OAI21_X1  g053(.A(G101), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n202), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n230), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n229), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT11), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(G137), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT11), .A3(G134), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G131), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT67), .B(G131), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n252), .A2(new_n246), .A3(new_n248), .A4(new_n249), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n231), .A2(new_n208), .A3(new_n232), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(G143), .B2(new_n207), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n224), .B1(new_n259), .B2(new_n205), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n256), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n257), .B1(new_n256), .B2(new_n260), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT82), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n202), .B2(new_n240), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n202), .A2(new_n240), .A3(new_n264), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n263), .B(KEYINPUT10), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n243), .A2(new_n255), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n270), .A2(G227), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n269), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT10), .B1(new_n266), .B2(new_n265), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n256), .A2(new_n260), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT71), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n256), .A2(new_n257), .A3(new_n260), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n242), .B(new_n229), .C1(new_n276), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n254), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n241), .A2(KEYINPUT82), .ZN(new_n283));
  OAI21_X1  g097(.A(G128), .B1(new_n214), .B2(new_n258), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n218), .A2(new_n232), .B1(new_n284), .B2(new_n224), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n202), .A2(new_n240), .A3(new_n264), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n202), .B(new_n240), .C1(new_n233), .C2(new_n235), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT12), .B1(new_n289), .B2(new_n254), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT12), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n291), .B(new_n255), .C1(new_n287), .C2(new_n288), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n268), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n275), .A2(new_n282), .B1(new_n293), .B2(new_n272), .ZN(new_n294));
  OAI21_X1  g108(.A(G469), .B1(new_n294), .B2(G902), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n281), .A2(new_n254), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n255), .B1(new_n243), .B2(new_n267), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n272), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n268), .B(new_n273), .C1(new_n290), .C2(new_n292), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT83), .B(G469), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G221), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT9), .B(G234), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT15), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT96), .ZN(new_n313));
  INV_X1    g127(.A(G217), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n305), .A2(new_n314), .A3(G953), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G128), .B(G143), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n205), .A2(G143), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT95), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT13), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT95), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n317), .B1(new_n323), .B2(G134), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(G134), .A3(new_n317), .ZN(new_n326));
  INV_X1    g140(.A(G122), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT94), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT94), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G122), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G116), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n327), .A2(G116), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n190), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G116), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n328), .B2(new_n330), .ZN(new_n337));
  OAI21_X1  g151(.A(G107), .B1(new_n337), .B2(new_n333), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n325), .A2(new_n326), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT14), .B1(new_n327), .B2(G116), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n336), .A3(G122), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G107), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n209), .A2(G128), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n345), .A2(new_n318), .A3(G134), .ZN(new_n346));
  AOI21_X1  g160(.A(G134), .B1(new_n345), .B2(new_n318), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n335), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n316), .B1(new_n339), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n190), .B1(new_n332), .B2(new_n334), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n337), .A2(G107), .A3(new_n333), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n323), .A2(G134), .A3(new_n317), .ZN(new_n353));
  OAI22_X1  g167(.A1(new_n351), .A2(new_n352), .B1(new_n353), .B2(new_n324), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n335), .A2(new_n344), .A3(new_n348), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n315), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n313), .B1(new_n357), .B2(new_n307), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n313), .A3(new_n307), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n312), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n358), .A2(new_n311), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT97), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n360), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n311), .B1(new_n364), .B2(new_n358), .ZN(new_n365));
  INV_X1    g179(.A(new_n362), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT97), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n370));
  NOR2_X1   g184(.A1(G237), .A2(G953), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(G143), .A3(G214), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(G143), .B1(new_n371), .B2(G214), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  XNOR2_X1  g190(.A(G125), .B(G140), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n207), .ZN(new_n378));
  INV_X1    g192(.A(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G125), .ZN(new_n380));
  INV_X1    g194(.A(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G146), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n375), .A2(new_n376), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT90), .ZN(new_n386));
  INV_X1    g200(.A(G237), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n270), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n209), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n372), .ZN(new_n390));
  INV_X1    g204(.A(new_n376), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n386), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI211_X1 g206(.A(KEYINPUT90), .B(new_n376), .C1(new_n389), .C2(new_n372), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n385), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n375), .B2(new_n252), .ZN(new_n396));
  INV_X1    g210(.A(new_n252), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n373), .B2(new_n374), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n389), .A2(new_n395), .A3(new_n252), .A4(new_n372), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n381), .A2(KEYINPUT16), .A3(G140), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT77), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n404), .B(G146), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n377), .A2(KEYINPUT19), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n377), .A2(KEYINPUT19), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n207), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n394), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G113), .B(G122), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(new_n187), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT91), .B1(new_n390), .B2(new_n397), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT17), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n398), .A4(new_n399), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n402), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT16), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n406), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n207), .B1(new_n423), .B2(new_n403), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n390), .A2(KEYINPUT17), .A3(new_n397), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n407), .A3(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n414), .B(new_n394), .C1(new_n420), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(G475), .A2(G902), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n429), .B(KEYINPUT92), .Z(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n370), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  AOI211_X1 g246(.A(KEYINPUT20), .B(new_n430), .C1(new_n416), .C2(new_n427), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n394), .B1(new_n420), .B2(new_n426), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n415), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n435), .B2(new_n427), .ZN(new_n436));
  XOR2_X1   g250(.A(KEYINPUT93), .B(G475), .Z(new_n437));
  OAI22_X1  g251(.A1(new_n432), .A2(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(G234), .A2(G237), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(G952), .A3(new_n270), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(G902), .A3(G953), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(G898), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n303), .A2(new_n309), .A3(new_n369), .A4(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n448));
  INV_X1    g262(.A(G113), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n336), .A2(G119), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT5), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT69), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n336), .B2(G119), .ZN(new_n454));
  INV_X1    g268(.A(G119), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT69), .A3(G116), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n336), .A2(G119), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n452), .B1(new_n458), .B2(new_n451), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n449), .A2(KEYINPUT2), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT2), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G113), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n463), .A2(new_n454), .A3(new_n456), .A4(new_n457), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n266), .B2(new_n265), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n460), .A2(new_n462), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n458), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n469), .A2(new_n464), .A3(KEYINPUT70), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT70), .B1(new_n469), .B2(new_n464), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n203), .B(new_n228), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n467), .A2(new_n472), .A3(new_n475), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT6), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n475), .B1(new_n467), .B2(new_n472), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n448), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n480), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n482), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n478), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G224), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(G953), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n219), .B1(new_n218), .B2(new_n206), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n226), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT86), .A3(G125), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(new_n277), .B2(G125), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(G125), .B2(new_n489), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n486), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(G125), .ZN(new_n496));
  INV_X1    g310(.A(new_n493), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n486), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n490), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n484), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G210), .B1(G237), .B2(G902), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(KEYINPUT7), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n490), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n475), .B(KEYINPUT8), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n465), .B1(new_n283), .B2(new_n286), .ZN(new_n508));
  INV_X1    g322(.A(new_n241), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n466), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n478), .A3(new_n511), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(KEYINPUT7), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n498), .B2(new_n490), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n307), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n503), .A2(new_n504), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n520));
  INV_X1    g334(.A(new_n504), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n501), .B1(new_n481), .B2(new_n483), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(new_n522), .B2(new_n517), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G214), .B1(G237), .B2(G902), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT84), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n503), .A2(new_n518), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(KEYINPUT88), .A3(new_n521), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n447), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G110), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT24), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT24), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G110), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT75), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G119), .B(G128), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n533), .B2(new_n535), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n205), .B(G119), .C1(KEYINPUT76), .C2(KEYINPUT23), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT23), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n455), .B2(G128), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT76), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n455), .B2(G128), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n541), .B1(G110), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n424), .A2(new_n407), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n378), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n539), .B1(new_n537), .B2(new_n540), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n532), .B(new_n542), .C1(new_n544), .C2(new_n546), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT78), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n554), .A2(new_n555), .A3(new_n407), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n554), .B2(new_n407), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n550), .B(new_n561), .C1(new_n556), .C2(new_n557), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n314), .B1(G234), .B2(new_n307), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n565), .A2(G902), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n307), .A3(new_n564), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT25), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n563), .A2(KEYINPUT25), .A3(new_n307), .A4(new_n564), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n567), .B1(new_n572), .B2(new_n566), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n226), .B(new_n254), .C1(new_n487), .C2(new_n488), .ZN(new_n575));
  INV_X1    g389(.A(new_n249), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n245), .A2(G137), .ZN(new_n577));
  OAI21_X1  g391(.A(G131), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n253), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(KEYINPUT68), .A3(new_n277), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT68), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n253), .A2(new_n578), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n285), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n575), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n470), .A2(new_n471), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n278), .A2(new_n279), .A3(new_n579), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(KEYINPUT30), .A3(new_n575), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n587), .A3(new_n575), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n371), .A2(G210), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT27), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT26), .B(G101), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n591), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT31), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT31), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n591), .A2(new_n599), .A3(new_n592), .A4(new_n596), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT28), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n592), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n584), .A2(new_n588), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n589), .A2(new_n587), .A3(KEYINPUT28), .A4(new_n575), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT72), .ZN(new_n606));
  INV_X1    g420(.A(new_n596), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n605), .B2(new_n607), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n598), .B(new_n600), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(G472), .A2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT73), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT32), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT73), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n610), .A2(new_n615), .A3(new_n611), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n610), .A2(new_n611), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n605), .A2(new_n596), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n591), .A2(new_n592), .A3(new_n607), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT29), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n587), .B1(new_n589), .B2(new_n575), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT74), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n592), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n592), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT28), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(KEYINPUT29), .A3(new_n596), .A4(new_n602), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n618), .A2(KEYINPUT32), .B1(G472), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n574), .B1(new_n617), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(KEYINPUT79), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT79), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n635), .B(new_n574), .C1(new_n617), .C2(new_n632), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n531), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  NAND2_X1  g452(.A1(new_n610), .A2(new_n307), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n613), .A2(new_n640), .A3(new_n616), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n303), .A2(new_n309), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n641), .A2(new_n642), .A3(new_n574), .ZN(new_n643));
  INV_X1    g457(.A(new_n445), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n310), .A2(G902), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT33), .B1(new_n357), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  AOI211_X1 g462(.A(KEYINPUT99), .B(new_n648), .C1(new_n350), .C2(new_n356), .ZN(new_n649));
  OAI211_X1 g463(.A(KEYINPUT100), .B(new_n645), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n357), .A2(new_n307), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n310), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n354), .A2(new_n355), .A3(new_n315), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n315), .B1(new_n354), .B2(new_n355), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n646), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n648), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n357), .A2(new_n646), .A3(KEYINPUT33), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT100), .B1(new_n659), .B2(new_n645), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n438), .B(new_n644), .C1(new_n653), .C2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n522), .A2(new_n521), .A3(new_n517), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n523), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n528), .A2(KEYINPUT98), .A3(new_n521), .ZN(new_n665));
  AOI211_X1 g479(.A(new_n526), .B(new_n661), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n643), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  NAND2_X1  g483(.A1(new_n428), .A2(new_n431), .ZN(new_n670));
  INV_X1    g484(.A(new_n370), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n428), .A2(new_n370), .A3(new_n431), .ZN(new_n673));
  INV_X1    g487(.A(new_n436), .ZN(new_n674));
  INV_X1    g488(.A(new_n437), .ZN(new_n675));
  AOI22_X1  g489(.A1(new_n672), .A2(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n363), .A2(new_n676), .A3(new_n368), .A4(new_n644), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n526), .B(new_n677), .C1(new_n664), .C2(new_n665), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n643), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G107), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  AND3_X1   g496(.A1(new_n610), .A2(new_n615), .A3(new_n611), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n615), .B1(new_n610), .B2(new_n611), .ZN(new_n684));
  INV_X1    g498(.A(G472), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n610), .B2(new_n307), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n558), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n566), .A2(G902), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n558), .A2(new_n687), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n572), .B2(new_n566), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n683), .A2(new_n684), .A3(new_n686), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n531), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  AOI21_X1  g510(.A(new_n308), .B1(new_n295), .B2(new_n302), .ZN(new_n697));
  INV_X1    g511(.A(new_n692), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n617), .B2(new_n632), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n664), .A2(new_n665), .ZN(new_n702));
  INV_X1    g516(.A(new_n673), .ZN(new_n703));
  OAI22_X1  g517(.A1(new_n703), .A2(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n442), .A2(G900), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n440), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n369), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n701), .A2(new_n702), .A3(new_n527), .A4(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n526), .B1(new_n664), .B2(new_n665), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n701), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n700), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n706), .B(KEYINPUT39), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n697), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n363), .A2(new_n368), .A3(new_n438), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n698), .A2(new_n717), .A3(new_n526), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n524), .A2(new_n529), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT38), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n524), .A2(KEYINPUT38), .A3(new_n529), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n697), .A2(new_n715), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT40), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n628), .A2(new_n596), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(G902), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n591), .A2(new_n592), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n596), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n685), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n618), .B2(KEYINPUT32), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n617), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n719), .A2(new_n724), .A3(new_n726), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G143), .ZN(G45));
  AND3_X1   g549(.A1(new_n303), .A2(new_n309), .A3(new_n698), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT32), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n631), .A2(G472), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n614), .B2(new_n612), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n438), .B(new_n706), .C1(new_n653), .C2(new_n660), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n710), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n207), .ZN(G48));
  INV_X1    g559(.A(KEYINPUT103), .ZN(new_n746));
  INV_X1    g560(.A(new_n299), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n273), .B1(new_n282), .B2(new_n268), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n307), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n746), .B1(new_n749), .B2(G469), .ZN(new_n750));
  INV_X1    g564(.A(G469), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n300), .A2(KEYINPUT103), .A3(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n309), .B(new_n302), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n749), .A2(new_n746), .A3(G469), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT103), .B1(new_n300), .B2(new_n751), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n758), .A3(new_n309), .A4(new_n302), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n633), .A2(new_n666), .A3(new_n754), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G15));
  NAND4_X1  g576(.A1(new_n633), .A2(new_n678), .A3(new_n754), .A4(new_n759), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G116), .ZN(G18));
  NAND3_X1  g578(.A1(new_n698), .A2(new_n369), .A3(new_n446), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n617), .B2(new_n632), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n710), .A3(new_n754), .A4(new_n759), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  AOI211_X1 g582(.A(new_n526), .B(new_n717), .C1(new_n664), .C2(new_n665), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n644), .A3(new_n754), .A4(new_n759), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n598), .A2(new_n600), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n601), .B1(new_n626), .B2(new_n627), .ZN(new_n772));
  INV_X1    g586(.A(new_n602), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n607), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n611), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n640), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n777), .A2(KEYINPUT105), .A3(new_n574), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT105), .ZN(new_n779));
  INV_X1    g593(.A(new_n611), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n771), .B2(new_n774), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n686), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n779), .B1(new_n782), .B2(new_n573), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n770), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n327), .ZN(G24));
  NOR4_X1   g600(.A1(new_n686), .A2(new_n781), .A3(new_n741), .A4(new_n692), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n754), .A2(new_n787), .A3(new_n710), .A4(new_n759), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G125), .ZN(G27));
  NAND2_X1  g603(.A1(new_n617), .A2(new_n632), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n573), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT106), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n720), .A2(new_n527), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n793), .B2(new_n642), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n526), .B1(new_n524), .B2(new_n529), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(KEYINPUT106), .A3(new_n697), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n791), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n741), .A2(KEYINPUT42), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n612), .A2(new_n614), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n574), .B1(new_n632), .B2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n795), .A2(KEYINPUT106), .A3(new_n697), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT106), .B1(new_n795), .B2(new_n697), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n742), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n797), .A2(new_n798), .B1(new_n803), .B2(KEYINPUT42), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G131), .ZN(G33));
  OAI211_X1 g619(.A(new_n633), .B(new_n708), .C1(new_n801), .C2(new_n802), .ZN(new_n806));
  XNOR2_X1  g620(.A(KEYINPUT107), .B(G134), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G36));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT20), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n428), .A2(new_n811), .A3(new_n431), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n672), .A2(new_n812), .B1(new_n674), .B2(new_n675), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n660), .B2(new_n653), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT43), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT43), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n813), .B(new_n816), .C1(new_n660), .C2(new_n653), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n698), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n809), .B1(new_n810), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n810), .A2(new_n818), .A3(new_n809), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT110), .B(new_n809), .C1(new_n810), .C2(new_n818), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT109), .B1(new_n720), .B2(new_n527), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT109), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n825), .B(new_n526), .C1(new_n524), .C2(new_n529), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT45), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n293), .A2(new_n272), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n274), .A2(new_n297), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n294), .A2(KEYINPUT45), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n833), .A3(G469), .ZN(new_n834));
  NAND2_X1  g648(.A1(G469), .A2(G902), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(KEYINPUT46), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT46), .B1(new_n834), .B2(new_n835), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n302), .B(new_n836), .C1(new_n837), .C2(KEYINPUT108), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n837), .A2(KEYINPUT108), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n309), .B(new_n715), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n828), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n247), .ZN(G39));
  OAI21_X1  g656(.A(new_n309), .B1(new_n838), .B2(new_n839), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT47), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n790), .A2(new_n793), .A3(new_n573), .A4(new_n741), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G140), .ZN(G42));
  NOR3_X1   g662(.A1(new_n574), .A2(new_n526), .A3(new_n308), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(KEYINPUT111), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n757), .A2(new_n302), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(KEYINPUT49), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n849), .A2(KEYINPUT111), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n850), .A2(new_n852), .A3(new_n853), .A4(new_n814), .ZN(new_n854));
  INV_X1    g668(.A(new_n733), .ZN(new_n855));
  INV_X1    g669(.A(new_n724), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n851), .A2(KEYINPUT49), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT112), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n365), .A2(new_n366), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n704), .A2(new_n860), .A3(new_n707), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT114), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n740), .A2(new_n793), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n797), .B2(new_n708), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n803), .A2(KEYINPUT42), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n797), .A2(new_n798), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n777), .A2(new_n692), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n742), .B(new_n867), .C1(new_n801), .C2(new_n802), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n361), .A2(new_n362), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT113), .B1(new_n870), .B2(new_n438), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n438), .B1(new_n653), .B2(new_n660), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n813), .A2(new_n873), .A3(new_n860), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n644), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n530), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n643), .A2(new_n877), .B1(new_n531), .B2(new_n693), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n878), .A2(new_n760), .A3(new_n767), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n763), .B1(new_n770), .B2(new_n784), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n881), .A3(new_n637), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n869), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n700), .A2(new_n710), .A3(new_n742), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n642), .A2(new_n698), .A3(new_n707), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n769), .A3(new_n733), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n712), .A2(new_n884), .A3(new_n788), .A4(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n878), .A2(new_n760), .A3(new_n767), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n880), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n740), .A2(new_n793), .A3(new_n862), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n893), .A2(new_n806), .A3(new_n868), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n892), .A2(new_n894), .A3(new_n804), .A4(new_n637), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n702), .A2(new_n527), .A3(new_n708), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT102), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n710), .A2(new_n701), .A3(new_n708), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n740), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n710), .A2(new_n754), .A3(new_n787), .A4(new_n759), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(new_n888), .A3(new_n884), .A4(new_n886), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n887), .A2(KEYINPUT52), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT52), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n895), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n890), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(KEYINPUT53), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n883), .A2(new_n889), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n906), .B1(new_n895), .B2(new_n904), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  OAI22_X1  g731(.A1(new_n909), .A2(new_n910), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n754), .A2(new_n759), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n795), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n815), .A2(new_n441), .A3(new_n817), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT117), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT48), .A4(new_n800), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n919), .A2(new_n710), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n784), .A2(new_n921), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n924), .A2(G952), .A3(new_n270), .A4(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT116), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n574), .A2(new_n440), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n855), .A2(new_n930), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n920), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n929), .B1(new_n920), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n872), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n922), .A2(new_n800), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n937));
  AOI211_X1 g751(.A(new_n928), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT51), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n843), .B(KEYINPUT47), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n309), .B2(new_n851), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n827), .A3(new_n926), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n438), .A2(new_n653), .A3(new_n660), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n932), .A2(new_n933), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n922), .A2(new_n867), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n926), .A2(new_n526), .A3(new_n856), .A4(new_n919), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT50), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n945), .B(new_n946), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n939), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n951), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(KEYINPUT51), .A3(new_n942), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n938), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n918), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(G952), .A2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n859), .B1(new_n956), .B2(new_n957), .ZN(G75));
  AND2_X1   g772(.A1(G210), .A2(G902), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n895), .A2(new_n904), .A3(new_n911), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n890), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT56), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n484), .A2(new_n502), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(new_n522), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT55), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n961), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n270), .A2(G952), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n961), .A2(new_n962), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(KEYINPUT118), .A3(new_n965), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT118), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT56), .B1(new_n915), .B2(new_n959), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(new_n966), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n972), .B2(new_n975), .ZN(G51));
  XNOR2_X1  g790(.A(new_n834), .B(KEYINPUT119), .ZN(new_n977));
  AND4_X1   g791(.A1(KEYINPUT120), .A2(new_n915), .A3(G902), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n307), .B1(new_n913), .B2(new_n914), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT120), .B1(new_n979), .B2(new_n977), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n835), .B(KEYINPUT57), .Z(new_n982));
  AND3_X1   g796(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n916), .B1(new_n913), .B2(new_n914), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n747), .A2(new_n748), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n968), .B1(new_n981), .B2(new_n988), .ZN(G54));
  AND2_X1   g803(.A1(KEYINPUT58), .A2(G475), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n979), .A2(new_n428), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n428), .B1(new_n979), .B2(new_n990), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n991), .A2(new_n992), .A3(new_n968), .ZN(G60));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT59), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n659), .B1(new_n918), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n995), .B1(new_n657), .B2(new_n658), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n983), .B2(new_n984), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n969), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n997), .A2(new_n1000), .ZN(G63));
  INV_X1    g815(.A(KEYINPUT61), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G217), .A2(G902), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT122), .ZN(new_n1004));
  XOR2_X1   g818(.A(KEYINPUT121), .B(KEYINPUT60), .Z(new_n1005));
  XOR2_X1   g819(.A(new_n1004), .B(new_n1005), .Z(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(new_n913), .B2(new_n914), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1008), .A2(new_n690), .A3(new_n688), .ZN(new_n1009));
  INV_X1    g823(.A(new_n565), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n969), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1002), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n915), .A2(new_n1006), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n968), .B1(new_n1013), .B2(new_n565), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1008), .A2(new_n690), .A3(new_n688), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1014), .A2(KEYINPUT61), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1012), .A2(new_n1016), .ZN(G66));
  OAI21_X1  g831(.A(G953), .B1(new_n444), .B2(new_n485), .ZN(new_n1018));
  INV_X1    g832(.A(new_n882), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(G953), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n481), .B(new_n483), .C1(G898), .C2(new_n270), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT123), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1020), .B(new_n1022), .ZN(G69));
  NAND2_X1  g837(.A1(new_n586), .A2(new_n590), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n408), .A2(new_n409), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(G900), .A2(G953), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n800), .A2(new_n769), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n840), .B1(new_n828), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n866), .A2(new_n865), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n899), .A2(new_n744), .A3(new_n900), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1031), .A2(new_n806), .A3(new_n847), .A4(new_n1032), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1026), .B(new_n1027), .C1(new_n1033), .C2(G953), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT127), .ZN(new_n1035));
  AND4_X1   g849(.A1(new_n697), .A2(new_n795), .A3(new_n715), .A4(new_n875), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1036), .B1(new_n634), .B2(new_n636), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1037), .B1(new_n828), .B2(new_n840), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT126), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g854(.A(KEYINPUT126), .B(new_n1037), .C1(new_n828), .C2(new_n840), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT125), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT62), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1032), .A2(new_n1043), .A3(new_n1044), .A4(new_n734), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n712), .A2(new_n734), .A3(new_n884), .A4(new_n788), .ZN(new_n1046));
  OAI21_X1  g860(.A(KEYINPUT125), .B1(new_n1046), .B2(KEYINPUT62), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g862(.A1(new_n845), .A2(new_n846), .B1(new_n1046), .B2(KEYINPUT62), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1042), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(new_n270), .ZN(new_n1051));
  XOR2_X1   g865(.A(new_n1026), .B(KEYINPUT124), .Z(new_n1052));
  INV_X1    g866(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1035), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI211_X1 g868(.A(KEYINPUT127), .B(new_n1052), .C1(new_n1050), .C2(new_n270), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1034), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n270), .B1(G227), .B2(G900), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1057), .ZN(new_n1059));
  OAI211_X1 g873(.A(new_n1059), .B(new_n1034), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1058), .A2(new_n1060), .ZN(G72));
  OR2_X1    g875(.A1(new_n1050), .A2(new_n882), .ZN(new_n1062));
  NAND2_X1  g876(.A1(G472), .A2(G902), .ZN(new_n1063));
  XOR2_X1   g877(.A(new_n1063), .B(KEYINPUT63), .Z(new_n1064));
  AOI21_X1  g878(.A(new_n730), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g879(.A1(new_n1033), .A2(new_n882), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n620), .B1(new_n1066), .B2(new_n1064), .ZN(new_n1067));
  NAND3_X1  g881(.A1(new_n730), .A2(new_n620), .A3(new_n1064), .ZN(new_n1068));
  NOR2_X1   g882(.A1(new_n909), .A2(new_n1068), .ZN(new_n1069));
  NOR4_X1   g883(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .A4(new_n968), .ZN(G57));
endmodule


