//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(new_n202), .A2(G50), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n210), .B(new_n214), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n207), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n208), .A2(G1), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(KEYINPUT69), .A3(G50), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT69), .ZN(new_n253));
  INV_X1    g0053(.A(G50), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n253), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n249), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G50), .B2(new_n245), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT70), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT8), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n208), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n264));
  INV_X1    g0064(.A(G150), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n248), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n258), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G222), .A2(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G223), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n276), .B(new_n279), .C1(G77), .C2(new_n272), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n244), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(new_n278), .A3(G274), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n278), .A2(new_n281), .ZN(new_n284));
  XOR2_X1   g0084(.A(KEYINPUT67), .B(G226), .Z(new_n285));
  OAI211_X1 g0085(.A(new_n280), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(G179), .B2(new_n286), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n271), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(G200), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n270), .A2(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n270), .A2(KEYINPUT9), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI211_X1 g0099(.A(KEYINPUT10), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n291), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n215), .A2(new_n208), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n267), .A2(new_n254), .B1(new_n262), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n248), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  XOR2_X1   g0105(.A(new_n305), .B(KEYINPUT11), .Z(new_n306));
  INV_X1    g0106(.A(KEYINPUT72), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n245), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n244), .A2(KEYINPUT72), .A3(G13), .A4(G20), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(KEYINPUT12), .A3(new_n216), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n245), .A2(G68), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(KEYINPUT12), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n311), .A2(new_n248), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G68), .A3(new_n251), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n228), .A2(G1698), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n272), .B(new_n320), .C1(G226), .C2(G1698), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n278), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n283), .B1(new_n217), .B2(new_n284), .ZN(new_n324));
  OR3_X1    g0124(.A1(new_n323), .A2(KEYINPUT13), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT13), .B1(new_n323), .B2(new_n324), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(G169), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n327), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n327), .B2(G169), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n319), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(G200), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n325), .A2(G190), .A3(new_n326), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n334), .A2(new_n315), .A3(new_n318), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n272), .A2(G238), .A3(G1698), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n272), .A2(G232), .A3(new_n274), .ZN(new_n339));
  INV_X1    g0139(.A(G107), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(new_n272), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n279), .ZN(new_n342));
  INV_X1    g0142(.A(G244), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n342), .B(new_n283), .C1(new_n343), .C2(new_n284), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n293), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G200), .B2(new_n344), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT8), .B(G58), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(new_n267), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n208), .A2(new_n303), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT71), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(new_n262), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n348), .A2(KEYINPUT71), .A3(new_n349), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n248), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n250), .A2(new_n303), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n316), .A2(new_n355), .B1(new_n303), .B2(new_n311), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(KEYINPUT73), .A3(new_n356), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n346), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n344), .A2(G179), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n287), .B2(new_n344), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n360), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n301), .A2(new_n337), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT76), .ZN(new_n368));
  AND2_X1   g0168(.A1(KEYINPUT65), .A2(G68), .ZN(new_n369));
  NOR2_X1   g0169(.A1(KEYINPUT65), .A2(G68), .ZN(new_n370));
  OAI21_X1  g0170(.A(G58), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n208), .B1(new_n371), .B2(new_n202), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n267), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n368), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G33), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT7), .B1(new_n380), .B2(new_n208), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  AOI211_X1 g0182(.A(new_n382), .B(G20), .C1(new_n377), .C2(new_n379), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n215), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n374), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n201), .B1(new_n215), .B2(G58), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT76), .B(new_n385), .C1(new_n386), .C2(new_n208), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n375), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n378), .A2(KEYINPUT75), .A3(G33), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n392), .A2(new_n377), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT7), .B1(new_n394), .B2(G20), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n377), .A3(new_n393), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n382), .A3(new_n208), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(G68), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n398), .A2(KEYINPUT16), .A3(new_n375), .A4(new_n387), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n390), .A2(new_n399), .A3(new_n248), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT77), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n390), .A2(new_n399), .A3(new_n402), .A4(new_n248), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n261), .A2(new_n250), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n249), .B1(new_n246), .B2(new_n261), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n278), .A2(G274), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n281), .ZN(new_n410));
  INV_X1    g0210(.A(new_n284), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(G232), .B2(new_n411), .ZN(new_n412));
  OR2_X1    g0212(.A1(G223), .A2(G1698), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G226), .B2(new_n274), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n396), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT78), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n279), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G169), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n412), .A2(new_n418), .A3(G179), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n407), .A2(new_n408), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G190), .B2(new_n419), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n404), .A2(new_n406), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n406), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n401), .B2(new_n403), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT18), .B1(new_n432), .B2(new_n422), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(KEYINPUT17), .A3(new_n427), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n424), .A2(new_n430), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n367), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n244), .A2(G33), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT79), .ZN(new_n440));
  INV_X1    g0240(.A(new_n248), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n440), .A2(G116), .A3(new_n310), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G116), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n311), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n247), .A2(new_n207), .B1(G20), .B2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  INV_X1    g0246(.A(G97), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n446), .B(new_n208), .C1(G33), .C2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT20), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n445), .A2(KEYINPUT20), .A3(new_n448), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n442), .B(new_n444), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G41), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n244), .B(G45), .C1(new_n452), .C2(KEYINPUT5), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G41), .ZN(new_n455));
  OAI211_X1 g0255(.A(G270), .B(new_n278), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT82), .B1(new_n454), .B2(G41), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT82), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(new_n452), .A3(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(G41), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n457), .A2(new_n459), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n456), .B1(new_n409), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G257), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n274), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(G264), .B2(new_n274), .ZN(new_n468));
  XOR2_X1   g0268(.A(KEYINPUT84), .B(G303), .Z(new_n469));
  OAI22_X1  g0269(.A1(new_n396), .A2(new_n468), .B1(new_n469), .B2(new_n272), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n279), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n451), .A2(new_n472), .A3(G169), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT21), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n464), .B1(new_n279), .B2(new_n470), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G190), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(G200), .ZN(new_n478));
  INV_X1    g0278(.A(new_n451), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n451), .A2(new_n472), .A3(KEYINPUT21), .A4(G169), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n465), .A2(new_n471), .A3(G179), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n451), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n475), .A2(new_n480), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT85), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n483), .A2(new_n481), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(KEYINPUT85), .A3(new_n475), .A4(new_n480), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  OAI21_X1  g0290(.A(G107), .B1(new_n381), .B2(new_n383), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  AND2_X1   g0292(.A1(G97), .A2(G107), .ZN(new_n493));
  NOR2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n340), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n441), .B1(new_n491), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n245), .A2(G97), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n440), .A2(new_n249), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n447), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n490), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(G20), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n266), .A2(G77), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n382), .B1(new_n272), .B2(G20), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n380), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n340), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n248), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n440), .A2(new_n249), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n500), .B1(new_n512), .B2(G97), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT80), .ZN(new_n514));
  AND2_X1   g0314(.A1(KEYINPUT4), .A2(G244), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n377), .A2(new_n379), .A3(new_n515), .A4(new_n274), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT81), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n272), .A2(new_n518), .A3(new_n274), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n343), .A2(G1698), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n392), .A2(new_n393), .A3(new_n521), .A4(new_n377), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n377), .A2(new_n379), .A3(G250), .A4(G1698), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n446), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n520), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n279), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n278), .B1(new_n453), .B2(new_n455), .ZN(new_n530));
  OAI22_X1  g0330(.A1(new_n530), .A2(new_n466), .B1(new_n463), .B2(new_n409), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(G200), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  AOI211_X1 g0333(.A(G190), .B(new_n531), .C1(new_n528), .C2(new_n279), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n504), .B(new_n514), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n511), .A2(new_n513), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n531), .B1(new_n528), .B2(new_n279), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n287), .ZN(new_n538));
  AOI211_X1 g0338(.A(new_n330), .B(new_n531), .C1(new_n528), .C2(new_n279), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT83), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n466), .A2(G1698), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(G250), .B2(G1698), .ZN(new_n545));
  INV_X1    g0345(.A(G294), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n396), .A2(new_n545), .B1(new_n376), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n279), .ZN(new_n548));
  INV_X1    g0348(.A(new_n530), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G264), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n463), .A2(new_n409), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n425), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n547), .A2(new_n279), .B1(new_n549), .B2(G264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n293), .A3(new_n551), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n245), .A2(G107), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n557), .B(KEYINPUT25), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n340), .B2(new_n502), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT22), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n208), .A2(G87), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(new_n380), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G116), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(G20), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n208), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n340), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n392), .A2(new_n393), .A3(new_n208), .A4(new_n377), .ZN(new_n570));
  INV_X1    g0370(.A(G87), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n560), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT24), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n393), .A2(new_n377), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(new_n208), .A3(new_n392), .A4(new_n572), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n562), .A4(new_n568), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n559), .B1(new_n580), .B2(new_n248), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n556), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n552), .A2(new_n287), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n554), .A2(new_n330), .A3(new_n551), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n441), .B1(new_n575), .B2(new_n579), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n559), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n208), .B1(new_n322), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n494), .A2(new_n571), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n588), .A2(new_n589), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(G68), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n570), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n248), .ZN(new_n594));
  INV_X1    g0394(.A(new_n351), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n440), .A2(new_n249), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n311), .A2(new_n351), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G238), .A2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n343), .B2(G1698), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n600), .A2(new_n377), .A3(new_n392), .A4(new_n393), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n278), .B1(new_n601), .B2(new_n563), .ZN(new_n602));
  INV_X1    g0402(.A(G250), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n461), .B2(G1), .ZN(new_n604));
  INV_X1    g0404(.A(G274), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n244), .A2(new_n605), .A3(G45), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n278), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n287), .B1(new_n602), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n343), .A2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(G238), .B2(G1698), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n563), .B1(new_n396), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n608), .B1(new_n612), .B2(new_n279), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n330), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n598), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(G200), .B1(new_n602), .B2(new_n608), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(G190), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n593), .A2(new_n248), .B1(new_n311), .B2(new_n351), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n512), .A2(G87), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n582), .A2(new_n586), .A3(new_n615), .A4(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n499), .A2(new_n490), .A3(new_n503), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT80), .B1(new_n511), .B2(new_n513), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n526), .B1(new_n523), .B2(new_n522), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n278), .B1(new_n625), .B2(new_n520), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n425), .B1(new_n626), .B2(new_n531), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n537), .A2(new_n293), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(G169), .B1(new_n626), .B2(new_n531), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n529), .A2(G179), .A3(new_n532), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n624), .A2(new_n629), .B1(new_n632), .B2(new_n536), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n621), .B1(new_n633), .B2(KEYINPUT83), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n438), .A2(new_n489), .A3(new_n543), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g0435(.A(new_n635), .B(KEYINPUT86), .Z(G372));
  INV_X1    g0436(.A(new_n365), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n336), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(new_n333), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n430), .A2(new_n434), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n433), .B(new_n424), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n299), .A2(new_n300), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n290), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n504), .A2(new_n514), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n632), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n620), .A2(new_n615), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n620), .A2(new_n615), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT26), .B1(new_n540), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n615), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n487), .A2(new_n475), .A3(new_n586), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n535), .A2(new_n540), .A3(new_n648), .A4(new_n582), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(KEYINPUT87), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT87), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n650), .B1(new_n581), .B2(new_n556), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n633), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT88), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n654), .A2(KEYINPUT87), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n633), .A2(new_n657), .A3(new_n656), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .A4(new_n653), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n652), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n643), .B1(new_n437), .B2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(G330), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n244), .A2(new_n208), .A3(G13), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n479), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n486), .B2(new_n488), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n487), .A2(new_n475), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(new_n674), .ZN(new_n677));
  OR3_X1    g0477(.A1(new_n675), .A2(KEYINPUT89), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT89), .B1(new_n675), .B2(new_n677), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n666), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n582), .B(new_n586), .C1(new_n581), .C2(new_n673), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n586), .B2(new_n673), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT90), .Z(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n676), .A2(new_n673), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n586), .A2(new_n672), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n684), .A2(new_n687), .A3(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n212), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n589), .A2(G116), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G1), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n206), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n693), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n633), .A2(new_n657), .A3(new_n653), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT26), .B1(new_n645), .B2(new_n650), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n648), .A2(new_n647), .A3(new_n536), .A4(new_n632), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n615), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n673), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT29), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n659), .A2(new_n663), .ZN(new_n707));
  INV_X1    g0507(.A(new_n652), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n672), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n706), .B1(new_n709), .B2(new_n705), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n476), .A2(G179), .A3(new_n554), .A4(new_n613), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n529), .A2(new_n532), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n476), .A2(G179), .ZN(new_n715));
  INV_X1    g0515(.A(new_n613), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n713), .A2(new_n715), .A3(new_n552), .A4(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n554), .A2(new_n613), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n537), .A3(new_n482), .A4(KEYINPUT30), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n714), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n673), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT91), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT91), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n720), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT92), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n673), .B1(new_n720), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n714), .A2(new_n717), .A3(new_n719), .A4(KEYINPUT92), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT31), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT93), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n720), .A2(new_n728), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n672), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n721), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n720), .A2(new_n725), .A3(new_n722), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n725), .B1(new_n720), .B2(new_n722), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT93), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n735), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n634), .A2(new_n489), .A3(new_n543), .A4(new_n673), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n732), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n710), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n698), .B1(new_n745), .B2(G1), .ZN(G364));
  AOI21_X1  g0546(.A(new_n207), .B1(G20), .B2(new_n287), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n208), .A2(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(G303), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n293), .A2(G179), .A3(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n208), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n749), .A2(new_n293), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n754), .A2(new_n546), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n208), .A2(new_n330), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n759), .A2(G190), .A3(new_n425), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT33), .B(G317), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n752), .B(new_n757), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n749), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G329), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n758), .A2(G190), .A3(new_n425), .ZN(new_n766));
  INV_X1    g0566(.A(G322), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n380), .B1(new_n764), .B2(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n758), .A2(KEYINPUT94), .A3(new_n763), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT94), .B1(new_n758), .B2(new_n763), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n768), .B1(new_n772), .B2(G311), .ZN(new_n773));
  INV_X1    g0573(.A(G326), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT96), .Z(new_n776));
  OAI211_X1 g0576(.A(new_n762), .B(new_n773), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n272), .B1(new_n766), .B2(new_n259), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n775), .A2(new_n254), .B1(new_n750), .B2(new_n571), .ZN(new_n779));
  INV_X1    g0579(.A(new_n754), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n778), .B(new_n779), .C1(G97), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n764), .A2(new_n373), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT95), .B(KEYINPUT32), .Z(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n755), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n782), .A2(new_n784), .B1(new_n785), .B2(G107), .ZN(new_n786));
  INV_X1    g0586(.A(new_n782), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n787), .A2(new_n783), .B1(new_n760), .B2(G68), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n772), .A2(G77), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n781), .A2(new_n786), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n748), .B1(new_n777), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G13), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n244), .B1(new_n793), .B2(G45), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n692), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n272), .A2(new_n212), .ZN(new_n797));
  INV_X1    g0597(.A(G355), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n798), .B1(G116), .B2(new_n212), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n239), .A2(new_n461), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n394), .A2(new_n691), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n461), .B2(new_n206), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n799), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n747), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n796), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n791), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n678), .A2(new_n679), .ZN(new_n812));
  INV_X1    g0612(.A(new_n807), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT97), .Z(new_n815));
  NOR2_X1   g0615(.A1(new_n680), .A2(new_n796), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(G330), .B2(new_n812), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(G396));
  NAND2_X1  g0618(.A1(new_n365), .A2(KEYINPUT98), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT98), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n363), .A2(new_n364), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n361), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n664), .A2(new_n672), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n364), .A2(new_n672), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n819), .A2(new_n361), .A3(new_n827), .A4(new_n821), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n637), .A2(new_n672), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n826), .B1(new_n709), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n796), .B1(new_n831), .B2(new_n743), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n743), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n747), .A2(new_n805), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n796), .B1(G77), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n760), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n837), .A2(new_n756), .B1(new_n340), .B2(new_n750), .ZN(new_n838));
  INV_X1    g0638(.A(new_n775), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(G303), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n772), .A2(G116), .ZN(new_n841));
  INV_X1    g0641(.A(G311), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n380), .B1(new_n764), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n766), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(G294), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n755), .A2(new_n571), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G97), .B2(new_n780), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n840), .A2(new_n841), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  INV_X1    g0649(.A(G143), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n849), .A2(new_n775), .B1(new_n766), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n771), .A2(new_n373), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(G150), .C2(new_n760), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT34), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n754), .A2(new_n259), .B1(new_n755), .B2(new_n592), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n394), .B1(new_n856), .B2(new_n764), .ZN(new_n857));
  INV_X1    g0657(.A(new_n750), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n855), .B(new_n857), .C1(G50), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n853), .A2(KEYINPUT34), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n848), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n836), .B1(new_n862), .B2(new_n747), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n830), .B2(new_n806), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n833), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n793), .A2(new_n244), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n337), .A2(new_n319), .A3(new_n672), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n319), .A2(new_n672), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n333), .A2(new_n336), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n730), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n741), .A2(new_n735), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n873), .A3(new_n830), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n407), .A2(new_n423), .ZN(new_n876));
  INV_X1    g0676(.A(new_n670), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n407), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n876), .A2(new_n878), .A3(new_n428), .A4(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n404), .A2(new_n406), .A3(new_n427), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n395), .A2(G68), .A3(new_n397), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n375), .A2(new_n387), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n389), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n248), .A3(new_n399), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n406), .A2(new_n885), .B1(new_n422), .B2(new_n670), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT99), .B(KEYINPUT37), .C1(new_n881), .C2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT99), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n432), .B2(new_n427), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n880), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n670), .B1(new_n885), .B2(new_n406), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n435), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n895));
  INV_X1    g0695(.A(new_n879), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n428), .B1(new_n432), .B2(new_n422), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n432), .A2(new_n670), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n880), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n435), .A2(new_n898), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n875), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n871), .A2(new_n873), .A3(new_n905), .A4(new_n830), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n892), .A2(new_n894), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT38), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n438), .A3(new_n873), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n910), .ZN(new_n915));
  INV_X1    g0715(.A(new_n906), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n903), .A2(KEYINPUT40), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n438), .A2(new_n873), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n914), .A2(G330), .A3(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT101), .Z(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n895), .B2(new_n902), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n333), .A2(new_n672), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n424), .A2(new_n433), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n670), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n822), .A2(new_n673), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n871), .B1(new_n825), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT38), .B1(new_n892), .B2(new_n894), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n895), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n931), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n929), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n643), .B1(new_n710), .B2(new_n437), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n867), .B1(new_n922), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n922), .B2(new_n941), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n944), .A2(new_n945), .A3(G116), .A4(new_n209), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n206), .A2(G77), .A3(new_n371), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(G50), .B2(new_n592), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n792), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n947), .A3(new_n950), .ZN(G367));
  OAI22_X1  g0751(.A1(new_n754), .A2(new_n340), .B1(new_n755), .B2(new_n447), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n776), .A2(new_n842), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(G294), .C2(new_n760), .ZN(new_n954));
  INV_X1    g0754(.A(G317), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n766), .A2(new_n469), .B1(new_n955), .B2(new_n764), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n750), .A2(new_n443), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n394), .B(new_n956), .C1(KEYINPUT46), .C2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(KEYINPUT46), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT103), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n772), .A2(G283), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n954), .A2(new_n958), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n754), .A2(new_n592), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n755), .A2(new_n303), .B1(new_n750), .B2(new_n259), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(G159), .C2(new_n760), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n272), .B1(new_n764), .B2(new_n849), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G150), .B2(new_n844), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n965), .B(new_n967), .C1(new_n254), .C2(new_n771), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n776), .A2(new_n850), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n747), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n618), .A2(new_n619), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n672), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n648), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n615), .B2(new_n974), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(new_n813), .ZN(new_n977));
  INV_X1    g0777(.A(new_n796), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n235), .A2(new_n802), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n809), .B1(new_n691), .B2(new_n595), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n972), .A2(new_n977), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n633), .B1(new_n624), .B2(new_n673), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n646), .A2(new_n672), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n687), .A2(new_n689), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT45), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n687), .A2(KEYINPUT45), .A3(new_n689), .A4(new_n985), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n985), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n682), .B(KEYINPUT90), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n685), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n991), .B1(new_n993), .B2(new_n688), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(KEYINPUT44), .B(new_n991), .C1(new_n993), .C2(new_n688), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n990), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n684), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n990), .A2(new_n998), .A3(new_n684), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n992), .B(new_n685), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n680), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n745), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n745), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n692), .B(KEYINPUT41), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n795), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n684), .A2(new_n991), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT42), .B1(new_n687), .B2(new_n991), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT42), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n993), .A2(new_n1014), .A3(new_n985), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n540), .B1(new_n991), .B2(new_n586), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n673), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT102), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT102), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1018), .A2(new_n1023), .A3(new_n1019), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1022), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1012), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1024), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1023), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1028), .A2(new_n1029), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n1011), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n982), .B1(new_n1010), .B2(new_n1033), .ZN(G387));
  OAI22_X1  g0834(.A1(new_n797), .A2(new_n694), .B1(G107), .B2(new_n212), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n231), .A2(new_n461), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n694), .ZN(new_n1037));
  AOI211_X1 g0837(.A(G45), .B(new_n1037), .C1(G68), .C2(G77), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n347), .A2(G50), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n802), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1035), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n796), .B1(new_n1042), .B2(new_n809), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n837), .A2(new_n261), .B1(new_n750), .B2(new_n303), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G159), .B2(new_n839), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n754), .A2(new_n351), .B1(new_n755), .B2(new_n447), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n766), .A2(new_n254), .B1(new_n764), .B2(new_n265), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n396), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1045), .B(new_n1048), .C1(new_n592), .C2(new_n771), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT104), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n760), .A2(G311), .B1(new_n844), .B2(G317), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n771), .B2(new_n469), .C1(new_n776), .C2(new_n767), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n780), .A2(G283), .B1(new_n858), .B2(G294), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n396), .B1(new_n764), .B2(new_n774), .C1(new_n443), .C2(new_n755), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1050), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1043), .B1(new_n1063), .B2(new_n747), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT105), .Z(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n992), .B2(new_n807), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1005), .B2(new_n795), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n745), .A2(new_n1005), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n692), .B(KEYINPUT106), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1006), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1067), .B1(new_n1068), .B2(new_n1070), .ZN(G393));
  AND3_X1   g0871(.A1(new_n990), .A2(new_n998), .A3(new_n684), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n684), .B1(new_n990), .B2(new_n998), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n795), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n837), .A2(new_n254), .B1(new_n216), .B2(new_n750), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n754), .A2(new_n303), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1076), .A2(new_n846), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n764), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n396), .B1(new_n1079), .B2(G143), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n347), .C2(new_n771), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n265), .A2(new_n775), .B1(new_n766), .B2(new_n373), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT51), .Z(new_n1083));
  NOR2_X1   g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n842), .A2(new_n766), .B1(new_n775), .B2(new_n955), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT52), .Z(new_n1086));
  AOI21_X1  g0886(.A(new_n272), .B1(new_n785), .B2(G107), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n443), .B2(new_n754), .C1(new_n837), .C2(new_n469), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n771), .A2(new_n546), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n750), .A2(new_n756), .B1(new_n764), .B2(new_n767), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT107), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n747), .B1(new_n1084), .B2(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n808), .B1(new_n447), .B2(new_n212), .C1(new_n802), .C2(new_n242), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n796), .A3(new_n1094), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT108), .Z(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n985), .B2(new_n813), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1075), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT109), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1006), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1074), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1003), .A2(KEYINPUT109), .A3(new_n1006), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1069), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1074), .B2(new_n1100), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1098), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G390));
  AOI22_X1  g0907(.A1(new_n880), .A2(new_n899), .B1(new_n435), .B2(new_n898), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n910), .B1(new_n1108), .B2(KEYINPUT38), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n932), .B1(new_n824), .B2(new_n703), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n927), .B1(new_n1110), .B2(new_n871), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT110), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT110), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1109), .A2(new_n1114), .A3(new_n1111), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n934), .A2(new_n926), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n924), .A2(new_n925), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n742), .A2(G330), .A3(new_n830), .A4(new_n871), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1116), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1115), .A2(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n871), .A2(new_n830), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n873), .A2(G330), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1121), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(new_n794), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1118), .A2(new_n805), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n261), .A2(new_n834), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n775), .A2(new_n756), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1131), .B(new_n1077), .C1(G107), .C2(new_n760), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n772), .A2(G97), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n380), .B1(new_n766), .B2(new_n443), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G294), .B2(new_n1079), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n858), .A2(G87), .B1(new_n785), .B2(G68), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n858), .A2(G150), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT54), .B(G143), .Z(new_n1140));
  NAND2_X1  g0940(.A1(new_n772), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n272), .B1(new_n766), .B2(new_n856), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G125), .B2(new_n1079), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G159), .A2(new_n780), .B1(new_n839), .B2(G128), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n760), .A2(G137), .B1(G50), .B2(new_n785), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1137), .B1(new_n1139), .B2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n978), .B(new_n1130), .C1(new_n1147), .C2(new_n747), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1128), .B1(new_n1129), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT112), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n367), .A2(G330), .A3(new_n436), .A4(new_n873), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n643), .B(new_n1151), .C1(new_n710), .C2(new_n437), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n742), .A2(G330), .A3(new_n830), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n871), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n1126), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n825), .A2(new_n933), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n873), .A2(G330), .A3(new_n830), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1154), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT111), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1110), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT111), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1160), .A2(new_n1164), .A3(new_n1154), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1120), .A4(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1150), .B(new_n1152), .C1(new_n1159), .C2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1125), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1166), .B1(new_n1157), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1152), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT112), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1127), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n1125), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n1121), .C1(new_n1167), .C2(new_n1171), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1069), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1149), .A2(new_n1177), .ZN(G378));
  XOR2_X1   g0978(.A(new_n1152), .B(KEYINPUT119), .Z(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n1172), .B2(new_n1127), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT57), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n270), .A2(new_n877), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT55), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n301), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n301), .A2(new_n1184), .ZN(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OR3_X1    g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n917), .B2(new_n666), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n905), .B1(new_n1109), .B2(new_n875), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1191), .B(G330), .C1(new_n1194), .C2(new_n911), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT120), .B1(new_n1196), .B2(new_n939), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1191), .B1(new_n913), .B2(G330), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1195), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n939), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n928), .A2(new_n937), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1193), .A2(new_n1201), .A3(new_n1195), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1197), .B1(new_n1203), .B2(KEYINPUT120), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1069), .B1(new_n1181), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT118), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1193), .A2(new_n1201), .A3(new_n1195), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1193), .A2(new_n1195), .B1(new_n929), .B2(new_n938), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1200), .A2(KEYINPUT118), .A3(new_n1202), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT57), .B1(new_n1211), .B2(new_n1180), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1205), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n796), .B1(G50), .B2(new_n835), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT115), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n775), .A2(new_n443), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n755), .A2(new_n259), .B1(new_n750), .B2(new_n303), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G97), .C2(new_n760), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n766), .A2(new_n340), .B1(new_n764), .B2(new_n756), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1219), .A2(new_n963), .A3(G41), .A4(new_n394), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n351), .C2(new_n771), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT114), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(G33), .A2(G41), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT113), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G50), .B(new_n1226), .C1(new_n452), .C2(new_n396), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n839), .A2(G125), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n837), .B2(new_n856), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G150), .B2(new_n780), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G128), .A2(new_n844), .B1(new_n858), .B2(new_n1140), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n849), .C2(new_n771), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  INV_X1    g1033(.A(G124), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1226), .B1(new_n1234), .B2(new_n764), .C1(new_n373), .C2(new_n755), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1232), .B2(KEYINPUT59), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1227), .B1(new_n1233), .B2(new_n1236), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1223), .A2(new_n1224), .A3(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1215), .B1(new_n748), .B2(new_n1238), .C1(new_n1191), .C2(new_n806), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT117), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1211), .B2(new_n795), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1213), .A2(new_n1241), .ZN(G375));
  NAND2_X1  g1042(.A1(new_n1169), .A2(new_n795), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1154), .A2(new_n805), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(KEYINPUT121), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(KEYINPUT121), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n796), .B1(G68), .B2(new_n835), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n766), .A2(new_n849), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n396), .B(new_n1248), .C1(G128), .C2(new_n1079), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n754), .A2(new_n254), .B1(new_n750), .B2(new_n373), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G132), .B2(new_n839), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n772), .A2(G150), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n760), .A2(new_n1140), .B1(G58), .B2(new_n785), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n837), .A2(new_n443), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n771), .A2(new_n340), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n380), .B1(new_n755), .B2(new_n303), .C1(new_n756), .C2(new_n766), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n754), .A2(new_n351), .B1(new_n775), .B2(new_n546), .ZN(new_n1258));
  OR4_X1    g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n750), .A2(new_n447), .B1(new_n764), .B2(new_n751), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT122), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1254), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1247), .B1(new_n1262), .B2(new_n747), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT123), .Z(new_n1264));
  NAND3_X1  g1064(.A1(new_n1245), .A2(new_n1246), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1243), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1169), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1152), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(new_n1008), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1266), .B1(new_n1270), .B2(new_n1172), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT124), .ZN(G381));
  OR4_X1    g1072(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1273));
  NOR4_X1   g1073(.A1(new_n1273), .A2(G387), .A3(G378), .A4(G381), .ZN(new_n1274));
  INV_X1    g1074(.A(G375), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(G407));
  AND2_X1   g1076(.A1(new_n1149), .A2(new_n1177), .ZN(new_n1277));
  INV_X1    g1077(.A(G213), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(G343), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G213), .B(G407), .C1(new_n1282), .C2(new_n1283), .ZN(G409));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G378), .B(new_n1241), .C1(new_n1205), .C2(new_n1212), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1207), .A2(new_n1208), .A3(new_n1206), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT118), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1009), .B(new_n1180), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1240), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1204), .B2(new_n794), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1277), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1286), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1279), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1069), .B1(new_n1268), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1172), .A2(KEYINPUT60), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1299), .B2(new_n1268), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n865), .B1(new_n1300), .B2(new_n1266), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1266), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1167), .A2(new_n1171), .A3(new_n1297), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1303), .A2(new_n1269), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G384), .B(new_n1302), .C1(new_n1304), .C2(new_n1298), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1285), .B1(new_n1296), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1279), .A2(G2897), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1301), .A2(new_n1305), .A3(new_n1308), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n982), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1025), .A2(new_n1026), .A3(new_n1012), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1011), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n744), .B1(new_n1074), .B2(new_n1005), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n794), .B1(new_n1318), .B2(new_n1008), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1314), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G390), .A2(new_n1320), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(G393), .B(G396), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G387), .A2(new_n1106), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1321), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1323), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1279), .B1(new_n1286), .B2(new_n1293), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1306), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(KEYINPUT63), .A3(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1307), .A2(new_n1313), .A3(new_n1327), .A4(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1328), .A2(new_n1329), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT61), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1334), .B1(new_n1328), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(KEYINPUT62), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1338), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1339));
  NOR3_X1   g1139(.A1(new_n1333), .A2(new_n1336), .A3(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT127), .ZN(new_n1341));
  NOR3_X1   g1141(.A1(new_n1325), .A2(new_n1326), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1322), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1321), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT127), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1342), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1331), .B1(new_n1340), .B2(new_n1348), .ZN(G405));
  AOI21_X1  g1149(.A(G378), .B1(new_n1213), .B2(new_n1241), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1286), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1329), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1277), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1353), .A2(new_n1306), .A3(new_n1286), .ZN(new_n1354));
  AND3_X1   g1154(.A1(new_n1347), .A2(new_n1352), .A3(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1347), .B1(new_n1352), .B2(new_n1354), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1355), .A2(new_n1356), .ZN(G402));
endmodule


