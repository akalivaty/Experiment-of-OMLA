

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595;

  INV_X1 U326 ( .A(n585), .ZN(n594) );
  XNOR2_X1 U327 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n389) );
  XNOR2_X1 U328 ( .A(n390), .B(n389), .ZN(n411) );
  XNOR2_X1 U329 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n376) );
  XNOR2_X1 U330 ( .A(n377), .B(n376), .ZN(n542) );
  INV_X1 U331 ( .A(n471), .ZN(n450) );
  INV_X1 U332 ( .A(G218GAT), .ZN(n452) );
  XNOR2_X1 U333 ( .A(n452), .B(KEYINPUT62), .ZN(n453) );
  XNOR2_X1 U334 ( .A(n454), .B(n453), .ZN(G1355GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n295) );
  XNOR2_X1 U336 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(n296), .B(G92GAT), .Z(n298) );
  XOR2_X1 U339 ( .A(G50GAT), .B(G162GAT), .Z(n425) );
  XNOR2_X1 U340 ( .A(G134GAT), .B(n425), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n308) );
  XOR2_X1 U342 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n300) );
  NAND2_X1 U343 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U345 ( .A(n301), .B(KEYINPUT78), .Z(n306) );
  XOR2_X1 U346 ( .A(G29GAT), .B(G43GAT), .Z(n303) );
  XNOR2_X1 U347 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n331) );
  XNOR2_X1 U349 ( .A(G36GAT), .B(G190GAT), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n304), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U351 ( .A(n331), .B(n381), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n313) );
  XOR2_X1 U354 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n310) );
  XNOR2_X1 U355 ( .A(G106GAT), .B(G85GAT), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U357 ( .A(G99GAT), .B(n311), .Z(n327) );
  INV_X1 U358 ( .A(n327), .ZN(n312) );
  XOR2_X1 U359 ( .A(n313), .B(n312), .Z(n570) );
  INV_X1 U360 ( .A(n570), .ZN(n556) );
  XNOR2_X1 U361 ( .A(KEYINPUT36), .B(n556), .ZN(n494) );
  XOR2_X1 U362 ( .A(G64GAT), .B(G92GAT), .Z(n315) );
  XNOR2_X1 U363 ( .A(G176GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n385) );
  XOR2_X1 U365 ( .A(KEYINPUT69), .B(n385), .Z(n317) );
  XOR2_X1 U366 ( .A(KEYINPUT71), .B(G148GAT), .Z(n416) );
  XNOR2_X1 U367 ( .A(G120GAT), .B(n416), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n323) );
  XOR2_X1 U369 ( .A(G57GAT), .B(KEYINPUT13), .Z(n319) );
  XNOR2_X1 U370 ( .A(G71GAT), .B(G78GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n346) );
  XOR2_X1 U372 ( .A(n346), .B(KEYINPUT32), .Z(n321) );
  NAND2_X1 U373 ( .A1(G230GAT), .A2(G233GAT), .ZN(n320) );
  XOR2_X1 U374 ( .A(n321), .B(n320), .Z(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n329) );
  XOR2_X1 U376 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n325) );
  XNOR2_X1 U377 ( .A(KEYINPUT31), .B(KEYINPUT74), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n590) );
  INV_X1 U381 ( .A(KEYINPUT41), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n590), .B(n330), .ZN(n563) );
  XOR2_X1 U383 ( .A(n331), .B(KEYINPUT29), .Z(n333) );
  NAND2_X1 U384 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U386 ( .A(G1GAT), .B(KEYINPUT68), .Z(n362) );
  XOR2_X1 U387 ( .A(n334), .B(n362), .Z(n336) );
  XNOR2_X1 U388 ( .A(G50GAT), .B(G36GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n344) );
  XOR2_X1 U390 ( .A(G22GAT), .B(G113GAT), .Z(n338) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(G15GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U393 ( .A(KEYINPUT30), .B(G8GAT), .Z(n340) );
  XNOR2_X1 U394 ( .A(G197GAT), .B(G141GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U396 ( .A(n342), .B(n341), .Z(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n371) );
  NAND2_X1 U398 ( .A1(n563), .A2(n371), .ZN(n345) );
  XNOR2_X1 U399 ( .A(KEYINPUT46), .B(n345), .ZN(n365) );
  XOR2_X1 U400 ( .A(G15GAT), .B(G127GAT), .Z(n435) );
  XNOR2_X1 U401 ( .A(n346), .B(n435), .ZN(n350) );
  INV_X1 U402 ( .A(n350), .ZN(n348) );
  AND2_X1 U403 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  INV_X1 U404 ( .A(n349), .ZN(n347) );
  NAND2_X1 U405 ( .A1(n348), .A2(n347), .ZN(n352) );
  NAND2_X1 U406 ( .A1(n350), .A2(n349), .ZN(n351) );
  NAND2_X1 U407 ( .A1(n352), .A2(n351), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n353), .B(KEYINPUT80), .ZN(n357) );
  XOR2_X1 U409 ( .A(KEYINPUT79), .B(G211GAT), .Z(n355) );
  XNOR2_X1 U410 ( .A(G8GAT), .B(G183GAT), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n378) );
  XOR2_X1 U412 ( .A(n378), .B(KEYINPUT12), .Z(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U414 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n359) );
  XNOR2_X1 U415 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n358) );
  XOR2_X1 U416 ( .A(n359), .B(n358), .Z(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n364) );
  XOR2_X1 U418 ( .A(G22GAT), .B(G155GAT), .Z(n420) );
  XNOR2_X1 U419 ( .A(n362), .B(n420), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U421 ( .A(n369), .B(KEYINPUT112), .Z(n582) );
  NAND2_X1 U422 ( .A1(n365), .A2(n582), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n366), .B(KEYINPUT113), .ZN(n367) );
  NAND2_X1 U424 ( .A1(n367), .A2(n556), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n368), .B(KEYINPUT47), .ZN(n375) );
  INV_X1 U426 ( .A(n369), .ZN(n462) );
  NOR2_X1 U427 ( .A1(n494), .A2(n462), .ZN(n370) );
  XNOR2_X1 U428 ( .A(KEYINPUT45), .B(n370), .ZN(n372) );
  INV_X1 U429 ( .A(n371), .ZN(n541) );
  NAND2_X1 U430 ( .A1(n372), .A2(n541), .ZN(n373) );
  NOR2_X1 U431 ( .A1(n373), .A2(n590), .ZN(n374) );
  NOR2_X1 U432 ( .A1(n375), .A2(n374), .ZN(n377) );
  XOR2_X1 U433 ( .A(G197GAT), .B(KEYINPUT21), .Z(n417) );
  XOR2_X1 U434 ( .A(n378), .B(n417), .Z(n380) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U437 ( .A(n382), .B(n381), .Z(n387) );
  XOR2_X1 U438 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n384) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n434) );
  XNOR2_X1 U441 ( .A(n434), .B(n385), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n518) );
  XOR2_X1 U443 ( .A(KEYINPUT119), .B(n518), .Z(n388) );
  NOR2_X1 U444 ( .A1(n542), .A2(n388), .ZN(n390) );
  XOR2_X1 U445 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n392) );
  XNOR2_X1 U446 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n406) );
  XOR2_X1 U448 ( .A(G148GAT), .B(G155GAT), .Z(n394) );
  XNOR2_X1 U449 ( .A(G127GAT), .B(G162GAT), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U451 ( .A(G57GAT), .B(KEYINPUT1), .Z(n396) );
  XNOR2_X1 U452 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U454 ( .A(n398), .B(n397), .Z(n404) );
  XNOR2_X1 U455 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n399), .B(KEYINPUT2), .ZN(n424) );
  XOR2_X1 U457 ( .A(G85GAT), .B(n424), .Z(n401) );
  NAND2_X1 U458 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U460 ( .A(G29GAT), .B(n402), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U463 ( .A(KEYINPUT84), .B(G134GAT), .Z(n408) );
  XNOR2_X1 U464 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U466 ( .A(G113GAT), .B(n409), .ZN(n447) );
  XNOR2_X1 U467 ( .A(n410), .B(n447), .ZN(n514) );
  NAND2_X1 U468 ( .A1(n411), .A2(n514), .ZN(n413) );
  INV_X1 U469 ( .A(KEYINPUT65), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n457) );
  INV_X1 U471 ( .A(n457), .ZN(n451) );
  XOR2_X1 U472 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n415) );
  XNOR2_X1 U473 ( .A(G211GAT), .B(KEYINPUT22), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n433) );
  XOR2_X1 U475 ( .A(G106GAT), .B(G218GAT), .Z(n419) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U478 ( .A(n421), .B(n420), .Z(n431) );
  XOR2_X1 U479 ( .A(G204GAT), .B(G78GAT), .Z(n423) );
  XNOR2_X1 U480 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n429) );
  XOR2_X1 U482 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(n433), .B(n432), .Z(n474) );
  XOR2_X1 U488 ( .A(n435), .B(n434), .Z(n437) );
  XNOR2_X1 U489 ( .A(G43GAT), .B(G99GAT), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U491 ( .A(KEYINPUT86), .B(G176GAT), .Z(n439) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U494 ( .A(n441), .B(n440), .Z(n446) );
  XOR2_X1 U495 ( .A(KEYINPUT85), .B(G183GAT), .Z(n443) );
  XNOR2_X1 U496 ( .A(G190GAT), .B(G71GAT), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n444), .B(KEYINPUT20), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n521) );
  NAND2_X1 U501 ( .A1(n474), .A2(n521), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n449), .B(KEYINPUT26), .ZN(n471) );
  NAND2_X1 U503 ( .A1(n451), .A2(n450), .ZN(n585) );
  NOR2_X1 U504 ( .A1(n494), .A2(n585), .ZN(n454) );
  XOR2_X1 U505 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n456) );
  XNOR2_X1 U506 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n455) );
  XOR2_X1 U507 ( .A(n456), .B(n455), .Z(n461) );
  NOR2_X1 U508 ( .A1(n474), .A2(n457), .ZN(n458) );
  XNOR2_X1 U509 ( .A(n458), .B(KEYINPUT55), .ZN(n459) );
  NOR2_X1 U510 ( .A1(n521), .A2(n459), .ZN(n577) );
  INV_X1 U511 ( .A(n577), .ZN(n581) );
  NOR2_X1 U512 ( .A1(n556), .A2(n581), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  INV_X1 U514 ( .A(n514), .ZN(n560) );
  NAND2_X1 U515 ( .A1(n556), .A2(n369), .ZN(n465) );
  XNOR2_X1 U516 ( .A(KEYINPUT82), .B(KEYINPUT16), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n463), .B(KEYINPUT83), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n465), .B(n464), .ZN(n481) );
  XOR2_X1 U519 ( .A(n518), .B(KEYINPUT91), .Z(n466) );
  XNOR2_X1 U520 ( .A(KEYINPUT27), .B(n466), .ZN(n470) );
  XNOR2_X1 U521 ( .A(n474), .B(KEYINPUT28), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT67), .ZN(n525) );
  INV_X1 U523 ( .A(n525), .ZN(n537) );
  OR2_X1 U524 ( .A1(n470), .A2(n537), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n514), .A2(n468), .ZN(n544) );
  XNOR2_X1 U526 ( .A(n544), .B(KEYINPUT92), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n469), .A2(n521), .ZN(n480) );
  NOR2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n559) );
  NOR2_X1 U529 ( .A1(n521), .A2(n518), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT93), .B(n472), .Z(n473) );
  NOR2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT25), .B(n475), .Z(n476) );
  NOR2_X1 U533 ( .A1(n559), .A2(n476), .ZN(n477) );
  NOR2_X1 U534 ( .A1(n560), .A2(n477), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT94), .B(n478), .Z(n479) );
  NAND2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n496) );
  NAND2_X1 U537 ( .A1(n481), .A2(n496), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT95), .B(n482), .Z(n512) );
  NOR2_X1 U539 ( .A1(n541), .A2(n590), .ZN(n483) );
  XNOR2_X1 U540 ( .A(KEYINPUT75), .B(n483), .ZN(n498) );
  NOR2_X1 U541 ( .A1(n512), .A2(n498), .ZN(n491) );
  NAND2_X1 U542 ( .A1(n560), .A2(n491), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(n484), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n487) );
  INV_X1 U546 ( .A(n518), .ZN(n531) );
  NAND2_X1 U547 ( .A1(n491), .A2(n531), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  INV_X1 U551 ( .A(n521), .ZN(n543) );
  NAND2_X1 U552 ( .A1(n491), .A2(n543), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U554 ( .A1(n537), .A2(n491), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n492), .B(KEYINPUT98), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G22GAT), .B(n493), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n501) );
  NOR2_X1 U558 ( .A1(n494), .A2(n369), .ZN(n495) );
  NAND2_X1 U559 ( .A1(n496), .A2(n495), .ZN(n497) );
  XOR2_X1 U560 ( .A(KEYINPUT37), .B(n497), .Z(n528) );
  OR2_X1 U561 ( .A1(n498), .A2(n528), .ZN(n499) );
  XOR2_X1 U562 ( .A(KEYINPUT38), .B(n499), .Z(n508) );
  NAND2_X1 U563 ( .A1(n560), .A2(n508), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U565 ( .A(G29GAT), .B(n502), .Z(G1328GAT) );
  NAND2_X1 U566 ( .A1(n508), .A2(n531), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n503), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U568 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n507) );
  XOR2_X1 U569 ( .A(G43GAT), .B(KEYINPUT101), .Z(n505) );
  NAND2_X1 U570 ( .A1(n508), .A2(n543), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(G1330GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n510) );
  NAND2_X1 U574 ( .A1(n508), .A2(n537), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  XNOR2_X1 U577 ( .A(n563), .B(KEYINPUT104), .ZN(n576) );
  NAND2_X1 U578 ( .A1(n541), .A2(n576), .ZN(n529) );
  NOR2_X1 U579 ( .A1(n512), .A2(n529), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n513), .B(KEYINPUT105), .ZN(n524) );
  NOR2_X1 U581 ( .A1(n514), .A2(n524), .ZN(n516) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n517), .Z(G1332GAT) );
  NOR2_X1 U585 ( .A1(n518), .A2(n524), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1333GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n524), .ZN(n522) );
  XOR2_X1 U589 ( .A(KEYINPUT108), .B(n522), .Z(n523) );
  XNOR2_X1 U590 ( .A(G71GAT), .B(n523), .ZN(G1334GAT) );
  NOR2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1335GAT) );
  NOR2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n560), .A2(n538), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(n530), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n538), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n543), .A2(n538), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n533), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n535) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U604 ( .A(KEYINPUT109), .B(n536), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1339GAT) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U608 ( .A1(n542), .A2(n545), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n371), .A2(n551), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U612 ( .A1(n551), .A2(n576), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n550) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n553) );
  INV_X1 U617 ( .A(n551), .ZN(n555) );
  NOR2_X1 U618 ( .A1(n582), .A2(n555), .ZN(n552) );
  XOR2_X1 U619 ( .A(n553), .B(n552), .Z(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT114), .B(n554), .ZN(G1342GAT) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n558) );
  XNOR2_X1 U622 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U625 ( .A1(n542), .A2(n561), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n371), .A2(n569), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n565) );
  NAND2_X1 U629 ( .A1(n569), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(n566), .ZN(G1345GAT) );
  XOR2_X1 U632 ( .A(G155GAT), .B(KEYINPUT117), .Z(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n369), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1346GAT) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(KEYINPUT118), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1347GAT) );
  NAND2_X1 U638 ( .A1(n577), .A2(n371), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G169GAT), .B(n575), .ZN(G1348GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1350GAT) );
  NAND2_X1 U649 ( .A1(n371), .A2(n594), .ZN(n589) );
  XOR2_X1 U650 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n587) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(G1352GAT) );
  XOR2_X1 U654 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n592) );
  NAND2_X1 U655 ( .A1(n594), .A2(n590), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(G204GAT), .B(n593), .Z(G1353GAT) );
  NAND2_X1 U658 ( .A1(n594), .A2(n369), .ZN(n595) );
  XNOR2_X1 U659 ( .A(n595), .B(G211GAT), .ZN(G1354GAT) );
endmodule

