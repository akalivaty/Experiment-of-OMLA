//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0007(.A(G97), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n213), .A2(new_n214), .B1(new_n202), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g0016(.A1(G77), .A2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n218), .B1(new_n208), .B2(new_n219), .C1(new_n209), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT67), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n216), .B(new_n217), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G116), .ZN(new_n224));
  INV_X1    g0024(.A(G270), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n223), .B1(new_n222), .B2(new_n221), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  NAND2_X1  g0029(.A1(new_n206), .A2(G50), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(G250), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n227), .A2(G13), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n235), .B(new_n237), .C1(new_n219), .C2(new_n220), .ZN(new_n238));
  AOI22_X1  g0038(.A1(new_n231), .A2(new_n234), .B1(KEYINPUT0), .B2(new_n238), .ZN(new_n239));
  OAI211_X1 g0039(.A(new_n229), .B(new_n239), .C1(KEYINPUT0), .C2(new_n238), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(G361));
  XOR2_X1   g0041(.A(G238), .B(G244), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n214), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G264), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n225), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n201), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT69), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(new_n213), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(G107), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(new_n224), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  OAI21_X1  g0058(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G150), .ZN(new_n261));
  XOR2_X1   g0061(.A(KEYINPUT8), .B(G58), .Z(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n259), .B(new_n261), .C1(new_n263), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n232), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT71), .B(G1), .ZN(new_n270));
  INV_X1    g0070(.A(G13), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n270), .A2(new_n271), .A3(new_n233), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n267), .A2(new_n269), .B1(new_n213), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT71), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n269), .B1(new_n278), .B2(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G50), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT9), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n264), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G222), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n289), .B1(new_n290), .B2(new_n287), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT73), .B1(new_n295), .B2(new_n232), .ZN(new_n296));
  INV_X1    g0096(.A(new_n232), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT73), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(new_n294), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G41), .A2(G45), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(new_n274), .A3(G274), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT72), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n270), .B2(new_n302), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n294), .A2(KEYINPUT70), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT70), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(G33), .A3(G41), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n310), .A3(new_n297), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n276), .A2(G1), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n313));
  OAI211_X1 g0113(.A(KEYINPUT72), .B(new_n303), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n307), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G226), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n305), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G200), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n283), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n282), .A2(KEYINPUT9), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n305), .A2(G190), .A3(new_n316), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n319), .A2(new_n320), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n283), .A2(new_n323), .A3(new_n318), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT10), .B1(new_n325), .B2(new_n321), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n317), .A2(G179), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT74), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n317), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n281), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n278), .A2(G13), .A3(G20), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n278), .A2(G33), .ZN(new_n335));
  INV_X1    g0135(.A(new_n269), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(G116), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n272), .A2(new_n224), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n224), .A2(G20), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n269), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G283), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n233), .C1(G33), .C2(new_n208), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT20), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  AND4_X1   g0143(.A1(KEYINPUT20), .A2(new_n342), .A3(new_n269), .A4(new_n339), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n337), .B(new_n338), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  OAI211_X1 g0147(.A(G257), .B(new_n288), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  OAI211_X1 g0148(.A(G264), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n285), .A2(G303), .A3(new_n286), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n300), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT5), .B(G41), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n278), .A2(new_n353), .A3(G45), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(G270), .A3(new_n311), .ZN(new_n355));
  INV_X1    g0155(.A(G45), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n275), .B2(new_n277), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n311), .A2(new_n357), .A3(G274), .A4(new_n353), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n345), .A2(new_n359), .A3(G169), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT21), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n360), .A2(KEYINPUT84), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT84), .B1(new_n360), .B2(new_n361), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n359), .A2(KEYINPUT21), .A3(G169), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n352), .A2(G179), .A3(new_n355), .A4(new_n358), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n345), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n359), .A2(G200), .ZN(new_n369));
  INV_X1    g0169(.A(new_n345), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n369), .B(new_n370), .C1(new_n371), .C2(new_n359), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n364), .A2(KEYINPUT85), .A3(new_n368), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n360), .A2(new_n361), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT84), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n360), .A2(KEYINPUT84), .A3(new_n361), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n368), .A3(new_n377), .A4(new_n372), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT85), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT19), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT82), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT82), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT19), .ZN(new_n385));
  AOI22_X1  g0185(.A1(G97), .A2(new_n265), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n233), .B(G68), .C1(new_n346), .C2(new_n347), .ZN(new_n388));
  AND2_X1   g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n383), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n390), .A2(new_n233), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n210), .A2(G87), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n387), .B(new_n388), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n393), .A2(new_n269), .B1(new_n272), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n334), .A2(new_n336), .A3(new_n335), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n396), .A2(new_n394), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G274), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n278), .A2(G45), .A3(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n400), .A2(new_n311), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n235), .B1(new_n270), .B2(new_n356), .ZN(new_n402));
  OAI211_X1 g0202(.A(G244), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n403));
  OAI211_X1 g0203(.A(G238), .B(new_n288), .C1(new_n346), .C2(new_n347), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n264), .C2(new_n224), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n401), .A2(new_n402), .B1(new_n405), .B2(new_n300), .ZN(new_n406));
  INV_X1    g0206(.A(G179), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n300), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n402), .A2(new_n400), .A3(new_n311), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n330), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n398), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT83), .B1(new_n411), .B2(new_n371), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT83), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n406), .A2(new_n415), .A3(G190), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(G200), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n272), .A2(new_n394), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n334), .A2(new_n335), .A3(G87), .A4(new_n336), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n392), .B1(new_n390), .B2(new_n233), .ZN(new_n421));
  INV_X1    g0221(.A(new_n388), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n421), .A2(new_n422), .A3(new_n386), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n419), .B(new_n420), .C1(new_n423), .C2(new_n336), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n413), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT23), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n427), .A2(new_n233), .A3(G107), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT23), .B1(new_n209), .B2(G20), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n233), .B(G87), .C1(new_n346), .C2(new_n347), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT22), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT22), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n287), .A2(new_n433), .A3(new_n233), .A4(G87), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n265), .A2(G116), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT24), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT24), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(new_n439), .A3(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n396), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n441), .A2(new_n269), .B1(G107), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT86), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n272), .A2(new_n444), .A3(new_n209), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT86), .B1(new_n334), .B2(G107), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT25), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT25), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(G257), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n452));
  OAI211_X1 g0252(.A(G250), .B(new_n288), .C1(new_n346), .C2(new_n347), .ZN(new_n453));
  INV_X1    g0253(.A(G294), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n264), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n300), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n354), .A2(G264), .A3(new_n311), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n358), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G200), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n354), .A2(new_n399), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n460), .A2(new_n311), .B1(new_n455), .B2(new_n300), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G190), .A3(new_n457), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n443), .A2(new_n451), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n432), .A2(new_n434), .ZN(new_n464));
  INV_X1    g0264(.A(new_n430), .ZN(new_n465));
  AND4_X1   g0265(.A1(new_n439), .A2(new_n464), .A3(new_n436), .A4(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n439), .B1(new_n435), .B2(new_n436), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n269), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n442), .A2(G107), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n451), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n456), .A2(G179), .A3(new_n358), .A4(new_n457), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT87), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n458), .A2(G169), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(new_n472), .A3(new_n471), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n470), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n463), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT81), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT7), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n285), .A2(new_n479), .A3(new_n233), .A4(new_n286), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n346), .A2(new_n347), .A3(G20), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n482));
  OAI211_X1 g0282(.A(G107), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n260), .A2(G77), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G97), .A2(G107), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT6), .B1(new_n210), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n487));
  OAI21_X1  g0287(.A(G20), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n489), .A2(new_n269), .B1(new_n208), .B2(new_n272), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n442), .A2(G97), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n354), .A2(G257), .A3(new_n311), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT80), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n354), .A2(KEYINPUT80), .A3(G257), .A4(new_n311), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(G244), .B(new_n288), .C1(new_n346), .C2(new_n347), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n287), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n341), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n300), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n497), .A2(new_n407), .A3(new_n358), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n492), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n495), .A2(new_n496), .B1(new_n311), .B2(new_n460), .ZN(new_n507));
  AOI21_X1  g0307(.A(G169), .B1(new_n507), .B2(new_n504), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n478), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n497), .A2(new_n358), .A3(new_n504), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n330), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n511), .A2(KEYINPUT81), .A3(new_n505), .A4(new_n492), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n510), .A2(new_n371), .ZN(new_n513));
  INV_X1    g0313(.A(G200), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n507), .B2(new_n504), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n492), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n509), .A2(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n381), .A2(new_n426), .A3(new_n477), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G58), .A2(G68), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n203), .A2(new_n205), .A3(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n287), .A2(new_n482), .A3(G20), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT77), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n346), .A2(new_n347), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT77), .B1(new_n285), .B2(new_n286), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n233), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n523), .B1(new_n527), .B2(new_n479), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT16), .B(new_n522), .C1(new_n528), .C2(new_n202), .ZN(new_n529));
  OAI211_X1 g0329(.A(G68), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n522), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT16), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n336), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n334), .A2(new_n263), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n279), .B2(new_n263), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G87), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n537), .B(KEYINPUT79), .ZN(new_n538));
  OAI211_X1 g0338(.A(G226), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n539));
  OAI211_X1 g0339(.A(G223), .B(new_n288), .C1(new_n346), .C2(new_n347), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n300), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n307), .A2(G232), .A3(new_n314), .A4(new_n311), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n543), .A3(new_n304), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G200), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n544), .A2(new_n371), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n534), .A2(new_n536), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT17), .ZN(new_n548));
  INV_X1    g0348(.A(new_n536), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n529), .B2(new_n533), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT17), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n545), .A4(new_n546), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n534), .A2(new_n536), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n544), .A2(G169), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n407), .B2(new_n544), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(KEYINPUT18), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT18), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n544), .A2(G169), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n544), .A2(new_n407), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n558), .B1(new_n561), .B2(new_n550), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n565));
  OAI221_X1 g0365(.A(new_n565), .B1(new_n209), .B2(new_n287), .C1(new_n291), .C2(new_n215), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n300), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n315), .A2(G244), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(G190), .A4(new_n304), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n569), .B(KEYINPUT75), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n262), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n266), .B2(new_n394), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n269), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n272), .A2(new_n290), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n279), .A2(G77), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n567), .A2(new_n304), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n568), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G200), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n570), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(G169), .B1(new_n578), .B2(new_n568), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n567), .A2(new_n568), .A3(new_n407), .A4(new_n304), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n576), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G226), .B(new_n288), .C1(new_n346), .C2(new_n347), .ZN(new_n587));
  OAI211_X1 g0387(.A(G232), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n588));
  INV_X1    g0388(.A(new_n389), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n300), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n307), .A2(G238), .A3(new_n314), .A4(new_n311), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n304), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT13), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT13), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n591), .A2(new_n592), .A3(new_n595), .A4(new_n304), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(new_n371), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n265), .A2(G77), .B1(new_n260), .B2(G50), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n233), .B2(G68), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n269), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n601), .B(KEYINPUT11), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n272), .A2(new_n202), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n279), .A2(G68), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n514), .B1(new_n594), .B2(new_n596), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n598), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n597), .A2(G169), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT14), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(KEYINPUT76), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n594), .A2(G179), .A3(new_n596), .ZN(new_n613));
  INV_X1    g0413(.A(new_n611), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n597), .A2(G169), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n608), .B1(new_n616), .B2(new_n606), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n586), .A2(new_n617), .ZN(new_n618));
  NOR4_X1   g0418(.A1(new_n333), .A2(new_n519), .A3(new_n564), .A4(new_n618), .ZN(G372));
  NOR3_X1   g0419(.A1(new_n333), .A2(new_n564), .A3(new_n618), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n476), .A2(new_n364), .A3(new_n368), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n424), .A2(KEYINPUT88), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n393), .A2(new_n269), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT88), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(new_n419), .A4(new_n420), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n413), .B1(new_n626), .B2(new_n418), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n518), .A2(new_n621), .A3(new_n463), .A4(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n398), .A2(new_n408), .A3(new_n412), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n511), .A2(new_n505), .A3(new_n492), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n509), .A2(new_n512), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT26), .B1(new_n635), .B2(new_n425), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n629), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n620), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n332), .ZN(new_n639));
  OR3_X1    g0439(.A1(new_n582), .A2(KEYINPUT89), .A3(new_n584), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT89), .B1(new_n582), .B2(new_n584), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n608), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n606), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n614), .B1(new_n597), .B2(G169), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n330), .B(new_n611), .C1(new_n594), .C2(new_n596), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n646), .B2(new_n613), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n553), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n563), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n639), .B1(new_n649), .B2(new_n327), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n638), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT90), .ZN(G369));
  NOR2_X1   g0452(.A1(new_n271), .A2(G20), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OR3_X1    g0454(.A1(new_n270), .A2(new_n654), .A3(KEYINPUT27), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT27), .B1(new_n270), .B2(new_n654), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(G213), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n370), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n373), .B2(new_n380), .ZN(new_n662));
  AOI211_X1 g0462(.A(new_n370), .B(new_n660), .C1(new_n364), .C2(new_n368), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G330), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n470), .A2(new_n659), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n477), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n476), .B2(new_n660), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n659), .B1(new_n364), .B2(new_n368), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n477), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n476), .B2(new_n659), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n671), .A2(new_n674), .ZN(G399));
  NOR2_X1   g0475(.A1(new_n237), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n392), .A2(new_n224), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(G1), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n230), .B2(new_n677), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n497), .A2(new_n358), .A3(new_n504), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n352), .A2(new_n355), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n471), .A2(new_n411), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n683), .A2(KEYINPUT30), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n497), .A2(new_n684), .A3(new_n358), .A4(new_n504), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n406), .A2(new_n461), .A3(G179), .A4(new_n457), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(G179), .B1(new_n461), .B2(new_n457), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n510), .A2(new_n691), .A3(new_n359), .A4(new_n411), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n686), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT31), .B1(new_n693), .B2(new_n659), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT91), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n659), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT91), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n516), .A2(new_n517), .ZN(new_n704));
  AND4_X1   g0504(.A1(new_n476), .A2(new_n635), .A3(new_n463), .A4(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(new_n381), .A3(new_n426), .A4(new_n660), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n665), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n637), .A2(new_n660), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n426), .A2(new_n633), .A3(new_n509), .A4(new_n512), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT26), .B1(new_n627), .B2(new_n631), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n629), .A2(new_n711), .A3(new_n712), .A4(new_n413), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n710), .B1(new_n713), .B2(new_n660), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n707), .A2(new_n709), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n682), .B1(new_n715), .B2(G1), .ZN(G364));
  NOR2_X1   g0516(.A1(G13), .A2(G33), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT94), .Z(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n664), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n653), .A2(G45), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n677), .A2(G1), .A3(new_n723), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n254), .A2(new_n356), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT93), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n725), .A2(new_n726), .B1(new_n356), .B2(new_n231), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n524), .B1(new_n346), .B2(new_n347), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n285), .A2(KEYINPUT77), .A3(new_n286), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n237), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n727), .B(new_n732), .C1(new_n726), .C2(new_n725), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n287), .A2(new_n236), .ZN(new_n734));
  XNOR2_X1  g0534(.A(G355), .B(KEYINPUT92), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n733), .B1(G116), .B2(new_n236), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT95), .B(G169), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n297), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n721), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n724), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(G20), .A2(G179), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT96), .Z(new_n744));
  NOR2_X1   g0544(.A1(new_n514), .A2(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g0546(.A(KEYINPUT33), .B(G317), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n514), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G322), .A2(new_n750), .B1(new_n751), .B2(G326), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G179), .A2(G200), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(G20), .A3(new_n371), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n287), .B1(new_n755), .B2(G329), .ZN(new_n756));
  INV_X1    g0556(.A(G303), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n233), .A2(G179), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n756), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n753), .A2(G190), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(G294), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G283), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n758), .A2(new_n745), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n752), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n744), .A2(new_n371), .A3(new_n514), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n748), .B(new_n766), .C1(G311), .C2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT97), .Z(new_n769));
  INV_X1    g0569(.A(new_n765), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n751), .A2(G50), .B1(G107), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G87), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n771), .B1(new_n772), .B2(new_n759), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n762), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n208), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n755), .A2(G159), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n777), .B1(KEYINPUT32), .B2(new_n778), .C1(new_n746), .C2(new_n202), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G77), .B2(new_n767), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(KEYINPUT32), .ZN(new_n781));
  INV_X1    g0581(.A(new_n287), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n750), .B2(G58), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n774), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n769), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT98), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n722), .B(new_n742), .C1(new_n786), .C2(new_n739), .ZN(new_n787));
  INV_X1    g0587(.A(new_n666), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n664), .A2(new_n665), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n788), .A2(new_n724), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n790), .ZN(G396));
  NOR2_X1   g0591(.A1(new_n577), .A2(new_n660), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n640), .A2(new_n641), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n586), .B2(new_n792), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n708), .A2(new_n794), .ZN(new_n795));
  AND3_X1   g0595(.A1(new_n640), .A2(new_n641), .A3(new_n792), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n792), .B1(new_n581), .B2(new_n585), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n637), .A2(new_n660), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(new_n707), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n707), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n801), .A2(new_n724), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n751), .ZN(new_n804));
  INV_X1    g0604(.A(G137), .ZN(new_n805));
  INV_X1    g0605(.A(G150), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n804), .A2(new_n805), .B1(new_n746), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G159), .B2(new_n767), .ZN(new_n808));
  INV_X1    g0608(.A(new_n750), .ZN(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT99), .B(G143), .Z(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n808), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT34), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n759), .A2(new_n213), .B1(new_n765), .B2(new_n202), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n730), .B(new_n814), .C1(G58), .C2(new_n762), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n813), .B(new_n815), .C1(new_n816), .C2(new_n754), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n804), .A2(new_n757), .ZN(new_n818));
  INV_X1    g0618(.A(new_n767), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n819), .A2(new_n224), .B1(new_n746), .B2(new_n764), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n782), .B1(new_n754), .B2(new_n822), .C1(new_n765), .C2(new_n772), .ZN(new_n823));
  INV_X1    g0623(.A(new_n759), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n776), .B(new_n823), .C1(G107), .C2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n821), .B(new_n825), .C1(new_n454), .C2(new_n809), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n817), .B1(new_n818), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n740), .A2(new_n717), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n827), .A2(new_n740), .B1(new_n290), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n718), .B2(new_n798), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n803), .B1(new_n724), .B2(new_n830), .ZN(G384));
  NOR2_X1   g0631(.A1(new_n486), .A2(new_n487), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT35), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n233), .B(new_n232), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n834), .B(G116), .C1(new_n833), .C2(new_n832), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT36), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n520), .A2(G77), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n230), .A2(new_n837), .B1(G50), .B2(new_n202), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(new_n271), .A3(new_n270), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT100), .ZN(new_n841));
  INV_X1    g0641(.A(new_n647), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n659), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT103), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n521), .A2(G20), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n260), .A2(G159), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n482), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n481), .ZN(new_n849));
  AOI21_X1  g0649(.A(G20), .B1(new_n728), .B2(new_n729), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(KEYINPUT7), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n532), .B(new_n847), .C1(new_n851), .C2(G68), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n531), .A2(new_n532), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n269), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n657), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n855), .A2(new_n549), .B1(new_n556), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n857), .A2(new_n858), .A3(new_n547), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n522), .B1(new_n528), .B2(new_n202), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(KEYINPUT16), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n851), .A2(G68), .ZN(new_n865));
  INV_X1    g0665(.A(new_n863), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n522), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(new_n867), .A3(new_n269), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n657), .B1(new_n868), .B2(new_n536), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n561), .B1(new_n868), .B2(new_n536), .ZN(new_n870));
  INV_X1    g0670(.A(new_n547), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n860), .B1(new_n872), .B2(new_n858), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n564), .A2(new_n869), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n866), .B1(new_n865), .B2(new_n522), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n847), .B(new_n863), .C1(new_n851), .C2(G68), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n876), .A2(new_n877), .A3(new_n336), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n856), .B1(new_n878), .B2(new_n549), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n556), .B1(new_n878), .B2(new_n549), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(new_n547), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n859), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n879), .B1(new_n553), .B2(new_n563), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT39), .B1(new_n875), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n869), .A2(new_n871), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n858), .B1(new_n887), .B2(new_n880), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n874), .B(KEYINPUT38), .C1(new_n888), .C2(new_n859), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n858), .B1(new_n857), .B2(new_n547), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n859), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n554), .A2(new_n856), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n553), .B2(new_n563), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n883), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n844), .B1(new_n886), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n883), .B1(new_n882), .B2(new_n884), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n890), .B1(new_n898), .B2(new_n889), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(KEYINPUT103), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n843), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n557), .A2(new_n562), .A3(new_n657), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n585), .A2(new_n659), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n799), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n647), .A2(new_n659), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT101), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n606), .A2(new_n659), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n617), .A2(new_n909), .B1(new_n647), .B2(new_n659), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n910), .B2(new_n907), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n875), .A2(new_n885), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n901), .A2(new_n902), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n620), .B1(new_n709), .B2(new_n714), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n650), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n694), .A2(new_n695), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n706), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n911), .A3(new_n798), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n920), .B1(new_n923), .B2(new_n913), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n920), .B1(new_n889), .B2(new_n895), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n925), .A2(new_n798), .A3(new_n911), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n620), .A2(new_n922), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n927), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(G330), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n919), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n278), .A2(new_n653), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n841), .B1(new_n932), .B2(new_n933), .ZN(G367));
  OAI21_X1  g0734(.A(new_n518), .B1(new_n517), .B2(new_n660), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n631), .A2(new_n660), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n635), .B1(new_n937), .B2(new_n476), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n660), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n673), .A2(new_n935), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT42), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n660), .B1(new_n622), .B2(new_n625), .ZN(new_n942));
  MUX2_X1   g0742(.A(new_n627), .B(new_n413), .S(new_n942), .Z(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n939), .A2(new_n941), .B1(KEYINPUT43), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n670), .A2(new_n937), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT104), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n948), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n676), .B(KEYINPUT41), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n937), .A2(new_n674), .A3(KEYINPUT105), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT105), .B1(new_n937), .B2(new_n674), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n937), .A2(new_n674), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT44), .Z(new_n960));
  NAND3_X1  g0760(.A1(new_n954), .A2(KEYINPUT45), .A3(new_n955), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT106), .B1(new_n962), .B2(new_n671), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n671), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n958), .A2(new_n960), .A3(new_n670), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n966), .B2(KEYINPUT106), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n669), .A2(new_n672), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n673), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n666), .A2(KEYINPUT107), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n666), .A2(KEYINPUT107), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n666), .A2(KEYINPUT107), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n971), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n715), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n967), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n953), .B1(new_n978), .B2(new_n715), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n723), .A2(G1), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT108), .Z(new_n981));
  OAI211_X1 g0781(.A(new_n950), .B(new_n951), .C1(new_n979), .C2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n770), .A2(G77), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n809), .B2(new_n806), .C1(new_n804), .C2(new_n811), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n782), .B1(new_n824), .B2(G58), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n202), .B2(new_n775), .C1(new_n805), .C2(new_n754), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(G159), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n988), .B2(new_n746), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G50), .B2(new_n767), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n809), .A2(new_n757), .B1(new_n991), .B2(new_n754), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n767), .A2(G283), .B1(G107), .B2(new_n762), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n454), .B2(new_n746), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n730), .B1(new_n804), .B2(new_n822), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n765), .A2(new_n208), .ZN(new_n996));
  NOR4_X1   g0796(.A1(new_n992), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n824), .A2(G116), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT46), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n990), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT47), .Z(new_n1001));
  AOI21_X1  g0801(.A(new_n724), .B1(new_n1001), .B2(new_n740), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n732), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n741), .B1(new_n236), .B2(new_n394), .C1(new_n249), .C2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(new_n720), .C2(new_n944), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT109), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n982), .A2(new_n1006), .ZN(G387));
  INV_X1    g0807(.A(KEYINPUT112), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n750), .A2(G317), .B1(new_n767), .B2(G303), .ZN(new_n1009));
  INV_X1    g0809(.A(G322), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1009), .B1(new_n822), .B2(new_n746), .C1(new_n1010), .C2(new_n804), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT48), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n764), .B2(new_n775), .C1(new_n454), .C2(new_n759), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n755), .A2(G326), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n731), .B1(G116), .B2(new_n770), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n213), .A2(new_n809), .B1(new_n804), .B2(new_n988), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n775), .A2(new_n394), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n754), .A2(new_n806), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n1021), .A2(new_n730), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n759), .A2(new_n290), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1020), .A2(new_n1023), .A3(new_n996), .A4(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n202), .B2(new_n819), .C1(new_n263), .C2(new_n746), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1019), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n724), .B1(new_n1027), .B2(new_n740), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n732), .B1(new_n245), .B2(new_n356), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n262), .A2(new_n213), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n678), .B1(new_n1030), .B2(KEYINPUT50), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(new_n356), .C1(KEYINPUT50), .C2(new_n1030), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G68), .B2(G77), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n679), .A2(new_n734), .B1(G107), .B2(new_n236), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT111), .Z(new_n1036));
  OAI21_X1  g0836(.A(new_n741), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n669), .A2(new_n720), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1028), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n975), .A2(new_n981), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(KEYINPUT110), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT110), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n975), .A2(new_n1042), .A3(new_n981), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1039), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n975), .A2(new_n715), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1045), .A2(new_n676), .A3(new_n976), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1008), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1044), .A2(new_n1008), .A3(new_n1046), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(G393));
  NAND3_X1  g0850(.A1(new_n964), .A2(new_n965), .A3(new_n981), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n937), .A2(new_n721), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n287), .B1(new_n770), .B2(G107), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n764), .B2(new_n759), .C1(new_n1010), .C2(new_n754), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT114), .Z(new_n1055));
  OAI22_X1  g0855(.A1(new_n819), .A2(new_n454), .B1(new_n746), .B2(new_n757), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G311), .A2(new_n750), .B1(new_n751), .B2(G317), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT52), .Z(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(new_n224), .C2(new_n775), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G150), .A2(new_n751), .B1(new_n750), .B2(G159), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT113), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT51), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(KEYINPUT51), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n824), .A2(G68), .B1(new_n770), .B2(G87), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n731), .C1(new_n290), .C2(new_n775), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n819), .A2(new_n263), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n746), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1066), .B(new_n1067), .C1(G50), .C2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1063), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n811), .A2(new_n754), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1060), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n724), .B1(new_n1072), .B2(new_n740), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n741), .B1(new_n208), .B2(new_n236), .C1(new_n257), .C2(new_n1003), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1052), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n677), .B1(new_n967), .B2(new_n977), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n966), .A2(new_n976), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(KEYINPUT115), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(KEYINPUT115), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1051), .B(new_n1075), .C1(new_n1079), .C2(new_n1080), .ZN(G390));
  INV_X1    g0881(.A(new_n843), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n912), .A2(new_n1082), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT103), .B1(new_n1084), .B2(new_n899), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n886), .A2(new_n844), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n843), .B1(new_n889), .B2(new_n895), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n713), .A2(new_n660), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n904), .B1(new_n1090), .B2(new_n794), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1089), .B1(new_n1091), .B2(new_n911), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n696), .B(new_n702), .C1(new_n519), .C2(new_n659), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n794), .A2(new_n665), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1094), .A2(new_n911), .A3(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1087), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n922), .A2(new_n911), .A3(new_n1095), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n981), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n224), .A2(new_n809), .B1(new_n804), .B2(new_n764), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n765), .A2(new_n202), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n775), .A2(new_n290), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n782), .B1(new_n754), .B2(new_n454), .C1(new_n759), .C2(new_n772), .ZN(new_n1105));
  NOR4_X1   g0905(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n208), .B2(new_n819), .C1(new_n209), .C2(new_n746), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n755), .A2(G125), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n824), .A2(G150), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n809), .A2(new_n816), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(G128), .C2(new_n751), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n287), .B1(new_n765), .B2(new_n213), .C1(new_n775), .C2(new_n988), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n767), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1112), .B(new_n1115), .C1(new_n805), .C2(new_n746), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1107), .B1(new_n1108), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1117), .A2(new_n740), .B1(new_n263), .B2(new_n828), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n718), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1100), .A2(new_n1101), .B1(new_n724), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n911), .B1(new_n922), .B2(new_n1095), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1096), .A2(new_n1122), .A3(new_n1091), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n911), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n905), .C1(new_n1098), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n922), .A2(new_n911), .A3(new_n1095), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n798), .A2(G330), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n703), .B2(new_n706), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(new_n1131), .B2(new_n911), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1125), .B1(new_n1132), .B2(new_n905), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1124), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n917), .B(new_n650), .C1(new_n665), .C2(new_n928), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1100), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1087), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n897), .A2(new_n900), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1092), .B1(new_n1140), .B2(new_n1083), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1141), .B2(new_n1098), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n905), .B1(new_n1098), .B2(new_n1126), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT116), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1127), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1135), .B1(new_n1145), .B2(new_n1124), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n677), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1121), .B1(new_n1138), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(G378));
  INV_X1    g0949(.A(KEYINPUT56), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n282), .A2(new_n657), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n333), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT55), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n333), .A2(new_n1151), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1153), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1150), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1157), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(KEYINPUT56), .A3(new_n1155), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n924), .A2(G330), .A3(new_n926), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n914), .B1(new_n1119), .B2(new_n843), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n902), .ZN(new_n1164));
  AND4_X1   g0964(.A1(new_n902), .A2(new_n901), .A3(new_n915), .A4(new_n1162), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1161), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1162), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n916), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1163), .A2(new_n902), .A3(new_n1162), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1168), .A2(new_n1169), .A3(new_n1160), .A4(new_n1158), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1135), .A2(KEYINPUT120), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1135), .A2(KEYINPUT120), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n1100), .C2(new_n1137), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1171), .A2(new_n1174), .A3(KEYINPUT57), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT121), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1171), .A2(new_n1174), .A3(KEYINPUT121), .A4(KEYINPUT57), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n677), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1158), .A2(new_n1160), .A3(new_n717), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n828), .A2(new_n213), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n819), .A2(new_n805), .B1(new_n746), .B2(new_n816), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n751), .A2(G125), .B1(G150), .B2(new_n762), .ZN(new_n1187));
  INV_X1    g0987(.A(G128), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n809), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1186), .B(new_n1189), .C1(new_n824), .C2(new_n1114), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT59), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G41), .B1(new_n755), .B2(G124), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G33), .B1(new_n770), .B2(G159), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n209), .A2(new_n809), .B1(new_n804), .B2(new_n224), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G41), .B(new_n1024), .C1(G283), .C2(new_n755), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n730), .C1(new_n202), .C2(new_n775), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n765), .A2(new_n201), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n819), .A2(new_n394), .B1(new_n746), .B2(new_n208), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G41), .B1(new_n731), .B2(G33), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1194), .B(new_n1202), .C1(G50), .C2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n724), .B1(new_n1204), .B2(new_n740), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1184), .A2(new_n1185), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT118), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT118), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1184), .A2(new_n1208), .A3(new_n1185), .A4(new_n1205), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(KEYINPUT119), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT119), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1171), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1211), .A2(new_n1213), .B1(new_n1214), .B2(new_n1101), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1183), .A2(new_n1216), .ZN(G375));
  OR2_X1    g1017(.A1(new_n911), .A2(new_n718), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n828), .A2(new_n202), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n764), .A2(new_n809), .B1(new_n804), .B2(new_n454), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n983), .B(new_n782), .C1(new_n208), .C2(new_n759), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1220), .A2(new_n1021), .A3(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n819), .A2(new_n209), .B1(new_n746), .B2(new_n224), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(new_n757), .C2(new_n754), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT123), .Z(new_n1226));
  NOR2_X1   g1026(.A1(new_n759), .A2(new_n988), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G132), .A2(new_n751), .B1(new_n750), .B2(G137), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n767), .A2(G150), .B1(new_n1068), .B2(new_n1114), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n730), .B1(G50), .B2(new_n762), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1198), .B1(G128), .B2(new_n755), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1226), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n724), .B1(new_n1233), .B2(new_n740), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1218), .A2(new_n1219), .A3(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1123), .B1(new_n1144), .B2(new_n1127), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n981), .B(KEYINPUT122), .Z(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1235), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT124), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1134), .A2(new_n1237), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT124), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n1235), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1135), .B(new_n1124), .C1(new_n1128), .C2(new_n1133), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1137), .A2(new_n952), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(G381));
  AOI21_X1  g1047(.A(new_n1215), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1148), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(G387), .A2(G381), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1048), .A2(new_n787), .A3(new_n790), .A4(new_n1049), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(G390), .A2(G384), .A3(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .ZN(G407));
  OAI211_X1 g1054(.A(G407), .B(G213), .C1(G343), .C2(new_n1249), .ZN(G409));
  INV_X1    g1055(.A(new_n1049), .ZN(new_n1256));
  OAI21_X1  g1056(.A(G396), .B1(new_n1256), .B2(new_n1047), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G390), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT115), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1078), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1260), .A2(new_n1264), .A3(new_n1051), .A4(new_n1075), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1259), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(G387), .ZN(new_n1267));
  INV_X1    g1067(.A(G387), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1259), .A2(new_n1265), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1245), .A2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1145), .A2(KEYINPUT60), .A3(new_n1135), .A4(new_n1124), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1137), .A3(new_n1273), .A4(new_n676), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1242), .B1(new_n1241), .B2(new_n1235), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1235), .ZN(new_n1276));
  AOI211_X1 g1076(.A(KEYINPUT124), .B(new_n1276), .C1(new_n1134), .C2(new_n1237), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1274), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(G384), .B(KEYINPUT125), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G384), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1244), .A2(new_n1282), .A3(new_n1274), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1280), .A2(KEYINPUT126), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT126), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1237), .B1(new_n1174), .B2(new_n952), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1148), .B(new_n1210), .C1(new_n1287), .C2(new_n1214), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n658), .A2(G213), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1286), .B(new_n1290), .C1(new_n1248), .C2(new_n1148), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1142), .A2(new_n1146), .B1(KEYINPUT120), .B2(new_n1135), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1293), .A2(new_n1172), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n676), .B1(new_n1294), .B2(KEYINPUT57), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1296));
  OAI21_X1  g1096(.A(G378), .B1(new_n1296), .B2(new_n1215), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1290), .A4(new_n1286), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1292), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(G375), .B2(G378), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1285), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1280), .A2(KEYINPUT126), .A3(new_n1283), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1289), .B1(new_n1306), .B2(G2897), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1307), .B1(new_n1306), .B2(G2897), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1304), .A2(new_n1305), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1280), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1283), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n658), .A2(G213), .A3(G2897), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1309), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1301), .B1(new_n1303), .B2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1270), .B1(new_n1300), .B2(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1259), .A2(new_n1265), .A3(new_n1268), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1268), .B1(new_n1259), .B2(new_n1265), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1286), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1286), .A2(new_n1308), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1290), .B1(new_n1248), .B2(new_n1148), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT63), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1291), .A2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1320), .A2(new_n1321), .A3(new_n1324), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1317), .A2(new_n1327), .ZN(G405));
  OAI211_X1 g1128(.A(new_n1297), .B(new_n1249), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1248), .A2(new_n1148), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1250), .A2(new_n1330), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1270), .B(new_n1329), .C1(new_n1331), .C2(new_n1312), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1329), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1312), .B1(new_n1297), .B2(new_n1249), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1320), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1332), .A2(new_n1335), .ZN(G402));
endmodule


