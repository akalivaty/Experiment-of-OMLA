//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT82), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT2), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT76), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT76), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n209), .A3(KEYINPUT2), .ZN(new_n210));
  AND2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n206), .A2(KEYINPUT75), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT75), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G155gat), .B2(G162gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n206), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n207), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G155gat), .B(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G211gat), .ZN(new_n226));
  INV_X1    g025(.A(G218gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G211gat), .A2(G218gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(KEYINPUT73), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(G197gat), .A2(G204gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G197gat), .ZN(new_n239));
  INV_X1    g038(.A(G204gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n241), .A2(new_n234), .B1(new_n232), .B2(new_n229), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n230), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT29), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n225), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n245));
  INV_X1    g044(.A(G228gat), .ZN(new_n246));
  INV_X1    g045(.A(G233gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n243), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n214), .A2(new_n218), .B1(new_n222), .B2(new_n223), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT29), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n205), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n250), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n219), .A2(new_n252), .A3(new_n224), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(KEYINPUT29), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(KEYINPUT82), .A3(new_n248), .A4(new_n245), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n228), .A2(new_n229), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT81), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n242), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n263), .B2(new_n242), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n237), .A2(KEYINPUT81), .A3(new_n262), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n254), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n251), .B1(new_n267), .B2(new_n252), .ZN(new_n268));
  OAI22_X1  g067(.A1(new_n268), .A2(new_n255), .B1(new_n246), .B2(new_n247), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT31), .B(G50gat), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n261), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(new_n261), .B2(new_n269), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n204), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n261), .A2(new_n269), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n270), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n261), .A2(new_n269), .A3(new_n271), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n203), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT65), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(G169gat), .A3(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OR3_X1    g083(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n284), .A2(new_n285), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT27), .B(G183gat), .ZN(new_n292));
  INV_X1    g091(.A(G190gat), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT28), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT27), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G183gat), .ZN(new_n298));
  AND4_X1   g097(.A1(KEYINPUT28), .A2(new_n296), .A3(new_n298), .A4(new_n293), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n290), .B(new_n291), .C1(new_n294), .C2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n291), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  INV_X1    g108(.A(G169gat), .ZN(new_n310));
  INV_X1    g109(.A(G176gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT23), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n284), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT25), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n312), .A2(new_n309), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n302), .A2(new_n303), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .A4(new_n284), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G134gat), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n320), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n325));
  INV_X1    g124(.A(G120gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(G113gat), .ZN(new_n327));
  INV_X1    g126(.A(G113gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(G120gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n328), .B2(G120gat), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT70), .B1(new_n326), .B2(G113gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n328), .A3(G120gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n326), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n332), .A2(new_n333), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n320), .A2(G127gat), .ZN(new_n338));
  INV_X1    g137(.A(G127gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G134gat), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n338), .A2(new_n340), .A3(new_n325), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n324), .A2(new_n330), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n337), .A2(new_n341), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n338), .A2(new_n340), .A3(new_n323), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n320), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G113gat), .B(G120gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n345), .B(new_n346), .C1(KEYINPUT1), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n300), .A2(new_n314), .A3(new_n349), .A4(new_n318), .ZN(new_n350));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT64), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n343), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT33), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT71), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT71), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  XNOR2_X1  g157(.A(G15gat), .B(G43gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n353), .B2(KEYINPUT32), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n356), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT34), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n343), .A2(new_n350), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(new_n351), .ZN(new_n367));
  AOI211_X1 g166(.A(KEYINPUT34), .B(new_n352), .C1(new_n343), .C2(new_n350), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n353), .B(KEYINPUT32), .C1(new_n354), .C2(new_n361), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n363), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n363), .B2(new_n370), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n279), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT29), .ZN(new_n377));
  AND4_X1   g176(.A1(new_n317), .A2(new_n284), .A3(new_n309), .A4(new_n312), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(new_n284), .A3(new_n315), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n316), .A2(new_n378), .B1(new_n380), .B2(KEYINPUT25), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n377), .B1(new_n381), .B2(new_n300), .ZN(new_n382));
  AND4_X1   g181(.A1(new_n375), .A2(new_n300), .A3(new_n314), .A4(new_n318), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n257), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n319), .B1(KEYINPUT29), .B2(new_n376), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n375), .A3(new_n300), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n250), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(KEYINPUT74), .B(new_n257), .C1(new_n382), .C2(new_n383), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT30), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n389), .A2(new_n390), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n393), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n396), .B(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n219), .A2(new_n224), .A3(new_n348), .A4(new_n344), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n251), .A2(new_n342), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n401), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n349), .B1(new_n251), .B2(new_n252), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n410), .B(new_n411), .C1(new_n412), .C2(new_n258), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n407), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n225), .A2(new_n349), .A3(KEYINPUT4), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n404), .B1(new_n251), .B2(new_n342), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n411), .B1(new_n412), .B2(new_n258), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT77), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n405), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(new_n349), .A3(new_n253), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT77), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n420), .A2(new_n422), .A3(new_n423), .A4(new_n411), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n411), .ZN(new_n426));
  INV_X1    g225(.A(new_n401), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n251), .A2(new_n342), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n216), .A2(G155gat), .A3(G162gat), .ZN(new_n432));
  INV_X1    g231(.A(G155gat), .ZN(new_n433));
  INV_X1    g232(.A(G162gat), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT75), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n206), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n209), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n438), .A2(new_n212), .A3(new_n211), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n439), .B2(new_n210), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n222), .A2(new_n223), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n349), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n401), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(KEYINPUT78), .A3(new_n426), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n410), .B1(new_n431), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n414), .B1(new_n425), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT0), .ZN(new_n448));
  XNOR2_X1  g247(.A(G57gat), .B(G85gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  AOI21_X1  g249(.A(KEYINPUT6), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n450), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT78), .B1(new_n443), .B2(new_n426), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n430), .B(new_n411), .C1(new_n442), .C2(new_n401), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT5), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n419), .B2(new_n424), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n452), .B1(new_n456), .B2(new_n414), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT6), .B(new_n452), .C1(new_n456), .C2(new_n414), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT80), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT80), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n451), .B2(new_n457), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n374), .B(new_n400), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n363), .A2(new_n370), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n367), .A2(new_n368), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n363), .B(new_n370), .C1(new_n367), .C2(new_n368), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(new_n399), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n425), .A2(new_n445), .ZN(new_n471));
  INV_X1    g270(.A(new_n414), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n450), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n446), .A2(new_n450), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n459), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n279), .A2(KEYINPUT35), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n470), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n369), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(KEYINPUT36), .A3(new_n371), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n483), .A3(new_n468), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n446), .A2(new_n474), .A3(new_n450), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n457), .B2(new_n451), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n394), .A2(KEYINPUT37), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n395), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n385), .A2(KEYINPUT83), .A3(new_n386), .A4(new_n250), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n490), .A2(KEYINPUT37), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n384), .A2(new_n387), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT38), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n489), .A2(new_n494), .B1(new_n397), .B2(new_n393), .ZN(new_n495));
  INV_X1    g294(.A(new_n397), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n496), .A2(KEYINPUT37), .B1(new_n395), .B2(new_n488), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT38), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT84), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n389), .A2(KEYINPUT37), .A3(new_n390), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n489), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT38), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n495), .A3(new_n499), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n406), .A2(new_n422), .A3(new_n408), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n426), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n443), .A2(new_n426), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n505), .A2(new_n508), .A3(new_n426), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n510), .A2(KEYINPUT40), .A3(new_n450), .A4(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n450), .B2(new_n446), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n511), .A2(new_n450), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT40), .B1(new_n514), .B2(new_n510), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n279), .B1(new_n516), .B2(new_n399), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n485), .B1(new_n504), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n462), .B1(new_n477), .B2(new_n461), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n279), .B1(new_n519), .B2(new_n399), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n464), .A2(new_n479), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n522));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G8gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n527), .A2(G1gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n529));
  INV_X1    g328(.A(G1gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT16), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n526), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n526), .A3(new_n532), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT88), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n537), .A2(new_n538), .A3(new_n533), .ZN(new_n539));
  XOR2_X1   g338(.A(G43gat), .B(G50gat), .Z(new_n540));
  INV_X1    g339(.A(G29gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n542));
  INV_X1    g341(.A(G36gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n541), .B2(KEYINPUT14), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(G29gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n540), .B1(new_n547), .B2(KEYINPUT15), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(KEYINPUT15), .B2(new_n547), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(KEYINPUT15), .A3(new_n540), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n536), .A2(new_n539), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n538), .B1(new_n537), .B2(new_n533), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n534), .A2(KEYINPUT88), .A3(new_n535), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n553), .A2(new_n554), .B1(new_n549), .B2(new_n550), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n525), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n549), .A2(KEYINPUT17), .A3(new_n550), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n558), .A2(new_n534), .A3(new_n535), .A4(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n551), .B1(new_n536), .B2(new_n539), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT18), .A4(new_n523), .ZN(new_n562));
  XNOR2_X1  g361(.A(G169gat), .B(G197gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT86), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n564), .B(KEYINPUT86), .ZN(new_n569));
  INV_X1    g368(.A(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n563), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n571), .A3(new_n563), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT12), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n576));
  INV_X1    g375(.A(new_n574), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(new_n572), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n556), .A2(new_n562), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n561), .A3(new_n523), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT18), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT90), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT90), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n583), .A2(new_n556), .A3(new_n562), .ZN(new_n588));
  INV_X1    g387(.A(new_n579), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n521), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT91), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n597), .A2(new_n601), .A3(new_n598), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n599), .B(KEYINPUT91), .C1(new_n594), .C2(new_n595), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT20), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n553), .A2(new_n554), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G134gat), .B(G162gat), .Z(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT96), .ZN(new_n625));
  OR2_X1    g424(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n626));
  NAND2_X1  g425(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n627));
  INV_X1    g426(.A(G85gat), .ZN(new_n628));
  INV_X1    g427(.A(G92gat), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G99gat), .A2(G106gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(KEYINPUT8), .A2(new_n631), .B1(new_n628), .B2(new_n629), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(G99gat), .A2(G106gat), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n634), .A2(new_n631), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT94), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n626), .A2(new_n627), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n628), .A2(new_n629), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n635), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n631), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT94), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n638), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n636), .A3(new_n631), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n643), .A2(new_n630), .A3(new_n632), .A4(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n641), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n558), .A2(new_n559), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT95), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n558), .A2(new_n652), .A3(new_n649), .A4(new_n559), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n551), .A2(new_n648), .B1(KEYINPUT41), .B2(new_n622), .ZN(new_n655));
  XOR2_X1   g454(.A(G190gat), .B(G218gat), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n654), .B2(new_n655), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n625), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n624), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n664), .A3(new_n658), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT98), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n641), .B1(new_n633), .B2(new_n639), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n645), .A2(new_n646), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n605), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n642), .A2(new_n647), .A3(new_n604), .A4(new_n603), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT10), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n648), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT97), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n669), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n675), .A2(KEYINPUT97), .A3(new_n676), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n672), .A2(new_n673), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n669), .ZN(new_n683));
  XNOR2_X1  g482(.A(G120gat), .B(G148gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(G176gat), .B(G204gat), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n684), .B(new_n685), .Z(new_n686));
  NAND3_X1  g485(.A1(new_n681), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n669), .B1(new_n675), .B2(new_n676), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n683), .ZN(new_n690));
  INV_X1    g489(.A(new_n686), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n620), .A2(new_n667), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n593), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n519), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(new_n530), .ZN(G1324gat));
  NOR2_X1   g500(.A1(new_n698), .A2(new_n400), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT16), .B(G8gat), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n526), .B2(new_n702), .ZN(new_n705));
  MUX2_X1   g504(.A(new_n704), .B(new_n705), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g505(.A(new_n485), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n698), .B2(new_n707), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n469), .A2(G15gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n698), .B2(new_n709), .ZN(G1326gat));
  INV_X1    g509(.A(new_n279), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n698), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT43), .B(G22gat), .Z(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(new_n693), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n620), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n666), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n593), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n541), .A3(new_n519), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n464), .A2(new_n479), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n518), .A2(new_n520), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n666), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT44), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n521), .B2(new_n666), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n587), .A2(new_n729), .A3(new_n590), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n587), .B2(new_n590), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G29gat), .B1(new_n735), .B2(new_n699), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n736), .ZN(G1328gat));
  NOR3_X1   g536(.A1(new_n718), .A2(G36gat), .A3(new_n400), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT46), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n735), .A2(new_n400), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(KEYINPUT101), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n740), .B2(KEYINPUT101), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(G1329gat));
  NAND4_X1  g542(.A1(new_n725), .A2(new_n727), .A3(new_n485), .A4(new_n734), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G43gat), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n469), .A2(G43gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n593), .A2(new_n717), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(KEYINPUT47), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n747), .B(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n751), .B2(new_n745), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(KEYINPUT104), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n754), .B(new_n749), .C1(new_n751), .C2(new_n745), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n748), .B1(new_n753), .B2(new_n755), .ZN(G1330gat));
  INV_X1    g555(.A(G50gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n719), .A2(new_n757), .A3(new_n279), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n735), .A2(new_n711), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n757), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT48), .B1(new_n758), .B2(KEYINPUT105), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI221_X1 g561(.A(new_n758), .B1(KEYINPUT105), .B2(KEYINPUT48), .C1(new_n759), .C2(new_n757), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(G1331gat));
  NAND2_X1  g563(.A1(new_n722), .A2(new_n723), .ZN(new_n765));
  NOR4_X1   g564(.A1(new_n620), .A2(new_n732), .A3(new_n667), .A4(new_n715), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n699), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g568(.A(new_n767), .B(KEYINPUT106), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n400), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  AND2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n771), .B2(new_n772), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n770), .B2(new_n707), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n469), .A2(G71gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n770), .A2(new_n711), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT107), .B(G78gat), .Z(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1335gat));
  NAND2_X1  g582(.A1(new_n733), .A2(new_n620), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n715), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n728), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n699), .ZN(new_n787));
  INV_X1    g586(.A(new_n784), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT51), .B1(new_n724), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  NOR4_X1   g589(.A1(new_n521), .A2(new_n790), .A3(new_n666), .A4(new_n784), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n519), .A2(new_n628), .A3(new_n693), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT108), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n787), .B1(new_n792), .B2(new_n794), .ZN(G1336gat));
  NOR3_X1   g594(.A1(new_n400), .A2(G92gat), .A3(new_n715), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n789), .B2(new_n791), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n725), .A2(new_n727), .A3(new_n399), .A4(new_n785), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G92gat), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT109), .B(new_n796), .C1(new_n789), .C2(new_n791), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT52), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n797), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n797), .A2(new_n808), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n809), .A2(new_n810), .A3(new_n801), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n806), .A2(new_n807), .A3(new_n812), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n786), .B2(new_n707), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n469), .A2(G99gat), .A3(new_n715), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n792), .B2(new_n815), .ZN(G1338gat));
  NAND4_X1  g615(.A1(new_n725), .A2(new_n727), .A3(new_n279), .A4(new_n785), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G106gat), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n711), .A2(new_n715), .A3(G106gat), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT112), .Z(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n789), .B2(new_n791), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n818), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n818), .B2(new_n825), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n821), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n818), .A2(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT114), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n818), .A2(new_n822), .A3(new_n825), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n830), .A2(new_n831), .B1(KEYINPUT53), .B2(new_n820), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n828), .A2(new_n832), .ZN(G1339gat));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n686), .B1(new_n688), .B2(new_n834), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n675), .A2(KEYINPUT97), .A3(new_n676), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT97), .B1(new_n675), .B2(new_n676), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n836), .A2(new_n837), .A3(new_n669), .ZN(new_n838));
  INV_X1    g637(.A(new_n669), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT54), .B1(new_n677), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT55), .B(new_n835), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n840), .B1(new_n680), .B2(new_n679), .ZN(new_n844));
  INV_X1    g643(.A(new_n835), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n842), .A2(new_n687), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n840), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n681), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT55), .A4(new_n835), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n732), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n552), .A2(new_n555), .A3(new_n525), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n523), .B1(new_n560), .B2(new_n561), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n574), .B(new_n573), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n587), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n693), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n667), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n666), .A2(new_n856), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n847), .A2(new_n860), .A3(new_n861), .A4(new_n851), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n665), .A3(new_n661), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n842), .A2(new_n851), .A3(new_n687), .A4(new_n846), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT116), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n620), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n694), .A2(new_n733), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n699), .B(new_n279), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n372), .A2(new_n373), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n400), .A3(new_n870), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n871), .A2(G113gat), .A3(new_n733), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n470), .ZN(new_n874));
  OAI21_X1  g673(.A(G113gat), .B1(new_n874), .B2(new_n592), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n873), .B1(new_n872), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(G1340gat));
  OAI21_X1  g677(.A(G120gat), .B1(new_n874), .B2(new_n715), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n693), .A2(new_n326), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT118), .Z(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n871), .B2(new_n881), .ZN(G1341gat));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n874), .A2(new_n620), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n339), .ZN(new_n885));
  INV_X1    g684(.A(new_n620), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n339), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n883), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  OAI221_X1 g688(.A(KEYINPUT119), .B1(new_n871), .B2(new_n887), .C1(new_n884), .C2(new_n339), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1342gat));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n870), .ZN(new_n892));
  NOR4_X1   g691(.A1(new_n892), .A2(G134gat), .A3(new_n399), .A4(new_n666), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n874), .B2(new_n666), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1343gat));
  INV_X1    g697(.A(G141gat), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n864), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n681), .A2(new_n683), .A3(new_n686), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n849), .A2(new_n835), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n843), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(KEYINPUT120), .A3(new_n851), .A4(new_n842), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n905), .A3(new_n591), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n667), .B1(new_n906), .B2(new_n858), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(new_n866), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n908), .A2(new_n620), .B1(new_n694), .B2(new_n733), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n711), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n699), .A2(new_n485), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n400), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n711), .B1(new_n867), .B2(new_n868), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT57), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n899), .B1(new_n917), .B2(new_n591), .ZN(new_n918));
  INV_X1    g717(.A(new_n913), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n912), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n592), .A2(G141gat), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g721(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n910), .A2(new_n732), .A3(new_n915), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n925), .A2(G141gat), .B1(new_n920), .B2(new_n921), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT58), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n918), .A2(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1344gat));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929));
  AOI211_X1 g728(.A(new_n929), .B(G148gat), .C1(new_n920), .C2(new_n693), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n916), .B2(new_n715), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n711), .A2(KEYINPUT57), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n863), .A2(new_n864), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n907), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n935), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n592), .B1(new_n864), .B2(new_n900), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n938), .A2(new_n905), .B1(new_n693), .B2(new_n857), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n937), .B(KEYINPUT122), .C1(new_n939), .C2(new_n667), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n620), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n696), .A2(new_n592), .A3(new_n697), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n933), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n913), .A2(new_n914), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n912), .A2(new_n929), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(new_n693), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n930), .B1(new_n948), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g748(.A(G155gat), .B1(new_n916), .B2(new_n620), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n920), .A2(new_n433), .A3(new_n886), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1346gat));
  OAI21_X1  g751(.A(G162gat), .B1(new_n916), .B2(new_n666), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n911), .A2(new_n434), .A3(new_n400), .A4(new_n667), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n919), .B2(new_n954), .ZN(G1347gat));
  NAND2_X1  g754(.A1(new_n867), .A2(new_n868), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n374), .A2(new_n399), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n519), .B1(new_n959), .B2(KEYINPUT123), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(KEYINPUT123), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n310), .A3(new_n732), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT124), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n519), .A2(new_n400), .ZN(new_n965));
  INV_X1    g764(.A(new_n469), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n711), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n957), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n310), .B1(new_n968), .B2(new_n591), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n964), .A2(new_n969), .ZN(G1348gat));
  NAND3_X1  g769(.A1(new_n962), .A2(new_n311), .A3(new_n693), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n957), .A2(new_n715), .A3(new_n967), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(new_n311), .ZN(G1349gat));
  NAND3_X1  g772(.A1(new_n962), .A2(new_n292), .A3(new_n886), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n620), .A3(new_n967), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(new_n295), .ZN(new_n976));
  XOR2_X1   g775(.A(KEYINPUT125), .B(KEYINPUT60), .Z(new_n977));
  XNOR2_X1  g776(.A(new_n976), .B(new_n977), .ZN(G1350gat));
  AOI21_X1  g777(.A(new_n293), .B1(new_n968), .B2(new_n667), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n979), .B(KEYINPUT61), .Z(new_n980));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n293), .A3(new_n667), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1351gat));
  NAND2_X1  g781(.A1(new_n941), .A2(new_n942), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(new_n932), .ZN(new_n984));
  INV_X1    g783(.A(new_n944), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n965), .A2(new_n707), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n988), .A2(new_n239), .A3(new_n592), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n919), .A2(new_n986), .ZN(new_n990));
  AOI21_X1  g789(.A(G197gat), .B1(new_n990), .B2(new_n732), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n989), .A2(new_n991), .ZN(G1352gat));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n993));
  AOI21_X1  g792(.A(G204gat), .B1(new_n993), .B2(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n990), .A2(new_n693), .A3(new_n994), .ZN(new_n995));
  OR3_X1    g794(.A1(new_n995), .A2(new_n993), .A3(KEYINPUT62), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n993), .B2(KEYINPUT62), .ZN(new_n997));
  NOR4_X1   g796(.A1(new_n943), .A2(new_n944), .A3(new_n715), .A4(new_n986), .ZN(new_n998));
  OAI211_X1 g797(.A(new_n996), .B(new_n997), .C1(new_n240), .C2(new_n998), .ZN(G1353gat));
  NAND3_X1  g798(.A1(new_n990), .A2(new_n226), .A3(new_n886), .ZN(new_n1000));
  OAI211_X1 g799(.A(KEYINPUT63), .B(G211gat), .C1(new_n988), .C2(new_n620), .ZN(new_n1001));
  INV_X1    g800(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n945), .A2(new_n886), .A3(new_n987), .ZN(new_n1003));
  AOI21_X1  g802(.A(KEYINPUT63), .B1(new_n1003), .B2(G211gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1000), .B1(new_n1002), .B2(new_n1004), .ZN(G1354gat));
  NAND3_X1  g804(.A1(new_n990), .A2(new_n227), .A3(new_n667), .ZN(new_n1006));
  NOR4_X1   g805(.A1(new_n943), .A2(new_n944), .A3(new_n666), .A4(new_n986), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1006), .B1(new_n1007), .B2(new_n227), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g809(.A(new_n1006), .B(KEYINPUT127), .C1(new_n1007), .C2(new_n227), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1355gat));
endmodule


