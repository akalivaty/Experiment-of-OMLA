//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G217), .ZN(new_n190));
  NOR3_X1   g004(.A1(new_n189), .A2(new_n190), .A3(G953), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  INV_X1    g006(.A(G122), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT86), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT86), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G122), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(new_n193), .B2(G116), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT87), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(new_n192), .A3(G122), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT86), .B(G122), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n203), .B(new_n198), .C1(new_n204), .C2(new_n192), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n197), .B1(new_n192), .B2(G122), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT65), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G128), .B(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n215), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT65), .B(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n208), .A2(new_n209), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n207), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT88), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n207), .A2(new_n223), .A3(new_n220), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT13), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(G128), .ZN(new_n228));
  OAI211_X1 g042(.A(G134), .B(new_n228), .C1(new_n217), .C2(new_n226), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n208), .A2(new_n209), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n208), .A2(new_n209), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n216), .B(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n191), .B1(new_n225), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n207), .A2(new_n223), .A3(new_n220), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n223), .B1(new_n207), .B2(new_n220), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n232), .B(new_n191), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n187), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G478), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT15), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n242));
  INV_X1    g056(.A(new_n191), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(G902), .B1(new_n244), .B2(new_n236), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(KEYINPUT89), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT89), .ZN(new_n247));
  AOI211_X1 g061(.A(new_n247), .B(G902), .C1(new_n244), .C2(new_n236), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n241), .B1(new_n249), .B2(new_n240), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT85), .ZN(new_n251));
  INV_X1    g065(.A(G475), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n187), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G237), .ZN(new_n256));
  INV_X1    g070(.A(G237), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  OAI211_X1 g072(.A(G214), .B(new_n254), .C1(new_n256), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n227), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(G237), .ZN(new_n262));
  AOI21_X1  g076(.A(G953), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(G143), .A3(G214), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT18), .A2(G131), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n260), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G125), .ZN(new_n267));
  INV_X1    g081(.A(G140), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(G125), .A2(G140), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G146), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n259), .A2(new_n227), .ZN(new_n274));
  AOI21_X1  g088(.A(G143), .B1(new_n263), .B2(G214), .ZN(new_n275));
  OAI21_X1  g089(.A(G131), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT18), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n266), .B(new_n273), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(G113), .B(G122), .Z(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT83), .ZN(new_n280));
  INV_X1    g094(.A(G104), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT17), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n260), .A2(new_n284), .A3(new_n264), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n276), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT16), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n269), .B2(new_n270), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n268), .A3(G125), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n272), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(G125), .A2(G140), .ZN(new_n292));
  NOR2_X1   g106(.A1(G125), .A2(G140), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT16), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(G146), .A3(new_n289), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(KEYINPUT73), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n294), .A2(new_n297), .A3(G146), .A4(new_n289), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT17), .B(G131), .C1(new_n274), .C2(new_n275), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n278), .B(new_n282), .C1(new_n286), .C2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n280), .B(G104), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n277), .B(new_n284), .C1(new_n260), .C2(new_n264), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n266), .A2(new_n273), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT19), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n271), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n269), .A2(KEYINPUT19), .A3(new_n270), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n295), .B1(new_n310), .B2(G146), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n276), .B2(new_n285), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n303), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n302), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n302), .A2(new_n313), .A3(KEYINPUT84), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n253), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT20), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n251), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n302), .A2(new_n313), .A3(KEYINPUT84), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT84), .B1(new_n302), .B2(new_n313), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT85), .B(KEYINPUT20), .C1(new_n323), .C2(new_n253), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n253), .A2(KEYINPUT20), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n314), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n254), .A2(G952), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(G234), .B2(G237), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT21), .B(G898), .Z(new_n331));
  NAND2_X1  g145(.A1(G234), .A2(G237), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(G902), .A3(G953), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n330), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n278), .B1(new_n286), .B2(new_n301), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n303), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n302), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n187), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G475), .ZN(new_n339));
  AND4_X1   g153(.A1(new_n250), .A2(new_n327), .A3(new_n334), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n271), .A2(new_n272), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n295), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G119), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G128), .ZN(new_n345));
  INV_X1    g159(.A(G128), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G119), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT24), .B(G110), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT23), .B1(new_n344), .B2(G128), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n346), .A3(G119), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n345), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n350), .B1(new_n355), .B2(G110), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT74), .B1(new_n343), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n351), .A2(new_n353), .B1(new_n344), .B2(G128), .ZN(new_n358));
  INV_X1    g172(.A(G110), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n358), .A2(new_n359), .B1(new_n348), .B2(new_n349), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n360), .A2(new_n342), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n348), .A2(new_n349), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n296), .A2(new_n363), .A3(new_n298), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT72), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n355), .A2(new_n365), .A3(G110), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT72), .B1(new_n358), .B2(new_n359), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI22_X1  g182(.A1(new_n357), .A2(new_n362), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n254), .A2(G221), .A3(G234), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT22), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(G137), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n343), .A2(new_n356), .A3(KEYINPUT74), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n361), .B1(new_n360), .B2(new_n342), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(new_n372), .C1(new_n364), .C2(new_n368), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n190), .B1(G234), .B2(new_n187), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G902), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n374), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT75), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n374), .A2(new_n378), .A3(new_n187), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT25), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n374), .A2(new_n378), .A3(new_n386), .A4(new_n187), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n379), .A3(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n383), .A2(KEYINPUT76), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT76), .B1(new_n383), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(G101), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n263), .A2(G210), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n398));
  INV_X1    g212(.A(G137), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n399), .A2(KEYINPUT11), .A3(G134), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(new_n214), .B2(G137), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n211), .A2(new_n213), .A3(new_n399), .ZN(new_n402));
  AND2_X1   g216(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n403));
  NOR2_X1   g217(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n401), .A2(new_n284), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n284), .B1(new_n401), .B2(new_n406), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n272), .A2(G143), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n227), .A2(G146), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OR2_X1    g225(.A1(KEYINPUT0), .A2(G128), .ZN(new_n412));
  NAND2_X1  g226(.A1(KEYINPUT0), .A2(G128), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT0), .A4(G128), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n414), .A2(KEYINPUT66), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT66), .B1(new_n414), .B2(new_n415), .ZN(new_n417));
  OAI22_X1  g231(.A1(new_n407), .A2(new_n408), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(G116), .B(G119), .Z(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT2), .B(G113), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n401), .A2(new_n406), .A3(new_n284), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n402), .B1(G134), .B2(new_n399), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G131), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n411), .A2(new_n346), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n227), .A2(KEYINPUT1), .A3(G146), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n346), .A2(KEYINPUT1), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n409), .A3(new_n410), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n423), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n418), .A2(new_n422), .A3(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n415), .B(new_n414), .C1(new_n407), .C2(new_n408), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n422), .B1(new_n433), .B2(new_n431), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n398), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n418), .A2(new_n422), .A3(new_n431), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT28), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n397), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n414), .A2(new_n415), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n402), .A2(new_n405), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n399), .A2(KEYINPUT11), .A3(G134), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n218), .B2(new_n399), .ZN(new_n444));
  OAI21_X1  g258(.A(G131), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n441), .B1(new_n445), .B2(new_n423), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n423), .A2(new_n425), .A3(new_n430), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n440), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n418), .A2(KEYINPUT30), .A3(new_n431), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n421), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n450), .A2(new_n397), .A3(new_n436), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n392), .B1(new_n439), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT70), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n422), .B1(new_n418), .B2(new_n431), .ZN(new_n454));
  OAI211_X1 g268(.A(KEYINPUT71), .B(KEYINPUT28), .C1(new_n432), .C2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n397), .A2(new_n392), .ZN(new_n456));
  INV_X1    g270(.A(new_n454), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n437), .B1(new_n457), .B2(new_n436), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT71), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n436), .B2(new_n437), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n455), .B(new_n456), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n461), .A2(new_n187), .ZN(new_n462));
  INV_X1    g276(.A(new_n398), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n421), .B1(new_n446), .B2(new_n447), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(new_n436), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n436), .A2(new_n437), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n396), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n450), .A2(new_n397), .A3(new_n436), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT70), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n392), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n453), .A2(new_n462), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n450), .A2(new_n396), .A3(new_n436), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT31), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n397), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT31), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n450), .A2(new_n477), .A3(new_n396), .A4(new_n436), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(G472), .A2(G902), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT32), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT32), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n479), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n391), .B1(new_n473), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G469), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(KEYINPUT80), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(KEYINPUT80), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT3), .B1(new_n281), .B2(G107), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n209), .A3(G104), .ZN(new_n494));
  INV_X1    g308(.A(G101), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n281), .A2(G107), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n492), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n209), .A2(G104), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n281), .A2(G107), .ZN(new_n499));
  OAI21_X1  g313(.A(G101), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(new_n430), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT78), .ZN(new_n503));
  AOI21_X1  g317(.A(G128), .B1(new_n409), .B2(new_n410), .ZN(new_n504));
  INV_X1    g318(.A(new_n427), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(G143), .B(G146), .ZN(new_n507));
  OAI211_X1 g321(.A(KEYINPUT78), .B(new_n427), .C1(new_n507), .C2(G128), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n429), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n502), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n407), .A2(new_n408), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n490), .B(new_n491), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n501), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n430), .B2(new_n501), .ZN(new_n514));
  INV_X1    g328(.A(new_n511), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT80), .A4(new_n489), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT4), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n518), .A3(G101), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT77), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(KEYINPUT77), .A3(new_n518), .A4(G101), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n517), .B2(G101), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n521), .A2(new_n522), .B1(new_n497), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT66), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n441), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n414), .A2(KEYINPUT66), .A3(new_n415), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT79), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n497), .A2(new_n500), .A3(KEYINPUT10), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n501), .A2(new_n430), .A3(KEYINPUT79), .A4(KEYINPUT10), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT10), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n513), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n529), .A2(new_n535), .A3(new_n537), .A4(new_n511), .ZN(new_n538));
  XNOR2_X1  g352(.A(G110), .B(G140), .ZN(new_n539));
  INV_X1    g353(.A(G227), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(G953), .ZN(new_n541));
  XOR2_X1   g355(.A(new_n539), .B(new_n541), .Z(new_n542));
  NAND4_X1  g356(.A1(new_n512), .A2(new_n516), .A3(new_n538), .A4(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n529), .A2(new_n535), .A3(new_n537), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n515), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n542), .B1(new_n546), .B2(new_n538), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n488), .B(new_n187), .C1(new_n544), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(G469), .A2(G902), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n512), .A2(new_n516), .A3(new_n538), .ZN(new_n550));
  INV_X1    g364(.A(new_n542), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n546), .A2(new_n538), .A3(new_n542), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(G469), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n548), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G221), .B1(new_n189), .B2(G902), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G214), .B1(G237), .B2(G902), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n521), .A2(new_n522), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n523), .A2(new_n497), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n421), .A3(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n419), .A2(new_n420), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT5), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n344), .A3(G116), .ZN(new_n564));
  OAI211_X1 g378(.A(G113), .B(new_n564), .C1(new_n419), .C2(new_n563), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n501), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G110), .B(G122), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT81), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n569), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n561), .A2(new_n571), .A3(new_n566), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(KEYINPUT6), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n441), .A2(G125), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n574), .B1(G125), .B2(new_n430), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n254), .A2(G224), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT82), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n575), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT6), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n567), .A2(new_n579), .A3(new_n569), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n565), .A2(new_n562), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n497), .A2(new_n500), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n566), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n569), .A2(KEYINPUT8), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n569), .A2(KEYINPUT8), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(new_n572), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n576), .A2(KEYINPUT7), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n575), .B(new_n590), .Z(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G210), .B1(G237), .B2(G902), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n581), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n593), .B1(new_n581), .B2(new_n592), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n558), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n557), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n340), .A2(new_n487), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  INV_X1    g414(.A(new_n482), .ZN(new_n601));
  INV_X1    g415(.A(G472), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n479), .B2(new_n187), .ZN(new_n603));
  INV_X1    g417(.A(new_n334), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n390), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n383), .A2(KEYINPUT76), .A3(new_n388), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n598), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n238), .A2(new_n247), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n245), .A2(KEYINPUT89), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n239), .A3(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n233), .A2(new_n237), .A3(KEYINPUT33), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n244), .B2(new_n236), .ZN(new_n616));
  OAI211_X1 g430(.A(G478), .B(new_n187), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n327), .A2(new_n339), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  NAND3_X1  g435(.A1(new_n611), .A2(new_n240), .A3(new_n612), .ZN(new_n622));
  INV_X1    g436(.A(new_n241), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n622), .A2(new_n623), .B1(G475), .B2(new_n338), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n325), .B1(new_n321), .B2(new_n322), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT90), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(KEYINPUT90), .B(new_n325), .C1(new_n321), .C2(new_n322), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n320), .A3(new_n324), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n609), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT91), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(G9));
  NOR2_X1   g450(.A1(new_n601), .A2(new_n603), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n369), .B(KEYINPUT92), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n373), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n380), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n641), .A2(new_n388), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n340), .A2(new_n598), .A3(new_n637), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT37), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n359), .ZN(G12));
  INV_X1    g460(.A(new_n558), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n581), .A2(new_n592), .ZN(new_n648));
  INV_X1    g462(.A(new_n593), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n647), .B1(new_n650), .B2(new_n594), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n330), .B1(new_n333), .B2(G900), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n631), .A2(KEYINPUT93), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n557), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n642), .B1(new_n473), .B2(new_n486), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n624), .A2(new_n630), .A3(new_n651), .A4(new_n652), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT93), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT94), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n652), .B(KEYINPUT39), .Z(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n555), .A2(new_n556), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT96), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(KEYINPUT96), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n666), .B1(new_n665), .B2(new_n667), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n457), .A2(new_n397), .A3(new_n436), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n187), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n397), .B1(new_n450), .B2(new_n436), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n479), .A2(new_n484), .A3(new_n481), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n484), .B1(new_n479), .B2(new_n481), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT95), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g493(.A(KEYINPUT95), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n643), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n327), .A2(new_n339), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n622), .A2(new_n623), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n595), .A2(new_n596), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT38), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n670), .A2(new_n558), .A3(new_n681), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  NAND3_X1  g503(.A1(new_n618), .A2(new_n598), .A3(new_n652), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n470), .B1(new_n469), .B2(new_n392), .ZN(new_n691));
  AOI211_X1 g505(.A(KEYINPUT70), .B(KEYINPUT29), .C1(new_n467), .C2(new_n468), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n602), .B1(new_n693), .B2(new_n462), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n675), .A2(new_n676), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n643), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n272), .ZN(G48));
  INV_X1    g512(.A(new_n538), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n524), .A2(new_n528), .B1(new_n513), .B2(new_n536), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n511), .B1(new_n700), .B2(new_n535), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n551), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n543), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n488), .B1(new_n703), .B2(new_n187), .ZN(new_n704));
  AOI211_X1 g518(.A(G469), .B(G902), .C1(new_n702), .C2(new_n543), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n651), .A3(new_n556), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n487), .A2(new_n334), .A3(new_n618), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n487), .A2(new_n631), .A3(new_n334), .A4(new_n708), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  NAND3_X1  g527(.A1(new_n340), .A2(new_n655), .A3(new_n708), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  NAND2_X1  g529(.A1(new_n475), .A2(new_n478), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT28), .B1(new_n432), .B2(new_n454), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n438), .A2(KEYINPUT71), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n396), .B1(new_n719), .B2(new_n455), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n481), .B1(new_n716), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT97), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n603), .ZN(new_n724));
  OAI211_X1 g538(.A(KEYINPUT97), .B(new_n481), .C1(new_n716), .C2(new_n720), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n383), .A2(new_n388), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT98), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT98), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n383), .A2(new_n729), .A3(new_n388), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n250), .B1(new_n339), .B2(new_n327), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n334), .A4(new_n708), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT99), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NOR3_X1   g550(.A1(new_n726), .A2(new_n707), .A3(new_n642), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT100), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n613), .A2(new_n617), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n738), .A2(new_n682), .A3(new_n739), .A4(new_n652), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n738), .B1(new_n618), .B2(new_n652), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  NAND3_X1  g557(.A1(new_n650), .A2(new_n558), .A3(new_n594), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n557), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n472), .A2(G472), .B1(new_n483), .B2(new_n485), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n746), .A2(new_n747), .A3(new_n731), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n745), .B(new_n748), .C1(new_n740), .C2(new_n741), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n608), .B(new_n745), .C1(new_n694), .C2(new_n695), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n682), .A2(new_n739), .A3(new_n652), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT100), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n618), .A2(new_n738), .A3(new_n652), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT102), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n284), .ZN(G33));
  INV_X1    g572(.A(new_n652), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n750), .A2(new_n632), .A3(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT103), .B(G134), .Z(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G36));
  NAND3_X1  g576(.A1(new_n327), .A2(new_n739), .A3(new_n339), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT105), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n327), .A2(new_n739), .A3(KEYINPUT43), .A4(new_n339), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n763), .A2(KEYINPUT105), .A3(new_n764), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n637), .A2(new_n642), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT106), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n744), .B1(new_n774), .B2(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n552), .A2(new_n553), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n552), .A2(KEYINPUT45), .A3(new_n553), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(G469), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n549), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n549), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n548), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n556), .A3(new_n663), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n786), .B1(new_n773), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n775), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  AND3_X1   g604(.A1(new_n785), .A2(KEYINPUT47), .A3(new_n556), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT47), .B1(new_n785), .B2(new_n556), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n746), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n751), .A2(new_n744), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(new_n608), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT107), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  NAND3_X1  g611(.A1(new_n706), .A2(new_n647), .A3(new_n556), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n686), .B1(new_n798), .B2(KEYINPUT113), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n770), .A2(new_n329), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n732), .ZN(new_n801));
  AOI211_X1 g615(.A(new_n799), .B(new_n801), .C1(KEYINPUT113), .C2(new_n798), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT50), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n679), .A2(new_n680), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n558), .A2(new_n706), .A3(new_n685), .A4(new_n556), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n608), .A3(new_n329), .A4(new_n805), .ZN(new_n806));
  OR3_X1    g620(.A1(new_n806), .A2(new_n682), .A3(new_n739), .ZN(new_n807));
  INV_X1    g621(.A(new_n556), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n792), .B(new_n791), .C1(new_n808), .C2(new_n706), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n801), .A2(new_n809), .A3(new_n744), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n726), .A2(new_n642), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n800), .A2(new_n805), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n803), .A2(new_n807), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n803), .A2(KEYINPUT51), .A3(new_n807), .A4(new_n813), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n682), .A2(new_n651), .A3(new_n683), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n681), .A2(new_n654), .A3(new_n652), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n751), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n598), .A3(new_n655), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n659), .A2(new_n742), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n752), .A2(new_n753), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n697), .B1(new_n827), .B2(new_n737), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(KEYINPUT52), .A3(new_n659), .A4(new_n820), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n825), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(KEYINPUT111), .A3(new_n824), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  INV_X1    g647(.A(new_n760), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n756), .A2(new_n834), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n746), .A2(new_n707), .A3(new_n391), .A4(new_n604), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n684), .A2(new_n707), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n726), .A2(new_n604), .A3(new_n731), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n836), .A2(new_n618), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n746), .A2(new_n642), .A3(new_n707), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n836), .A2(new_n631), .B1(new_n840), .B2(new_n340), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n811), .B(new_n745), .C1(new_n740), .C2(new_n741), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n745), .A2(new_n630), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n683), .A2(new_n759), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n655), .A3(new_n339), .A4(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n839), .A2(new_n841), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n835), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n327), .A2(new_n683), .A3(new_n339), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT108), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n327), .A2(new_n683), .A3(KEYINPUT108), .A4(new_n339), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n609), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n250), .A2(new_n327), .A3(new_n334), .A4(new_n339), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n651), .A2(new_n556), .A3(new_n555), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n724), .A2(new_n482), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n642), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT109), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n850), .A2(new_n851), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n610), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT109), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n644), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n857), .A2(new_n861), .A3(new_n599), .A4(new_n619), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT110), .B1(new_n847), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n835), .A2(new_n862), .A3(new_n846), .A4(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n832), .B(new_n833), .C1(new_n864), .C2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n709), .A2(new_n734), .A3(new_n712), .A4(new_n714), .ZN(new_n868));
  INV_X1    g682(.A(new_n845), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n756), .A3(new_n834), .A4(new_n842), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n865), .B1(new_n871), .B2(new_n862), .ZN(new_n872));
  INV_X1    g686(.A(new_n835), .ZN(new_n873));
  INV_X1    g687(.A(new_n846), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n863), .A3(KEYINPUT110), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n825), .A2(new_n829), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT112), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n825), .A2(KEYINPUT112), .A3(new_n829), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n872), .A2(new_n875), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n867), .B(KEYINPUT54), .C1(new_n833), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n746), .A2(new_n731), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n812), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT48), .Z(new_n884));
  NOR2_X1   g698(.A1(new_n801), .A2(new_n707), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n328), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n682), .A2(new_n739), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n806), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n871), .A2(new_n862), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n832), .A2(KEYINPUT53), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n890), .B(new_n891), .C1(new_n880), .C2(KEYINPUT53), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n881), .A2(new_n886), .A3(new_n888), .A4(new_n892), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n818), .A2(new_n893), .B1(G952), .B2(G953), .ZN(new_n894));
  NOR4_X1   g708(.A1(new_n763), .A2(new_n731), .A3(new_n647), .A4(new_n808), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n706), .B(KEYINPUT49), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n804), .A3(new_n686), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(G75));
  NAND2_X1  g712(.A1(new_n573), .A2(new_n580), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n578), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT114), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT112), .B1(new_n825), .B2(new_n829), .ZN(new_n906));
  INV_X1    g720(.A(new_n879), .ZN(new_n907));
  OAI22_X1  g721(.A1(new_n864), .A2(new_n866), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n833), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n187), .B1(new_n909), .B2(new_n890), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G210), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n905), .B1(new_n911), .B2(new_n903), .ZN(new_n912));
  AOI211_X1 g726(.A(KEYINPUT56), .B(new_n904), .C1(new_n910), .C2(G210), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n254), .A2(G952), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G51));
  NAND2_X1  g729(.A1(new_n872), .A2(new_n875), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n878), .A2(new_n879), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT53), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND4_X1   g732(.A1(KEYINPUT53), .A2(new_n889), .A3(new_n831), .A4(new_n830), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT54), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n892), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n549), .A2(KEYINPUT57), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n549), .A2(KEYINPUT57), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n703), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n780), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n910), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n914), .B1(new_n925), .B2(new_n927), .ZN(G54));
  INV_X1    g742(.A(new_n914), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n909), .A2(new_n890), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(new_n323), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n323), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT115), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n931), .A2(KEYINPUT115), .A3(new_n323), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G60));
  NOR2_X1   g751(.A1(new_n614), .A2(new_n616), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n920), .B2(new_n892), .ZN(new_n939));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT59), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n939), .A2(KEYINPUT116), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT116), .B1(new_n939), .B2(new_n942), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n881), .B2(new_n892), .ZN(new_n945));
  INV_X1    g759(.A(new_n938), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n929), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(G63));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  XOR2_X1   g763(.A(KEYINPUT118), .B(KEYINPUT60), .Z(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT119), .ZN(new_n951));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n951), .B(new_n952), .Z(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n918), .B2(new_n919), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n374), .A2(new_n378), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n914), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n640), .B(new_n953), .C1(new_n918), .C2(new_n919), .ZN(new_n957));
  AOI211_X1 g771(.A(KEYINPUT117), .B(new_n949), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n953), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n909), .B2(new_n890), .ZN(new_n960));
  INV_X1    g774(.A(new_n955), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n929), .B(new_n957), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT117), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT61), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n958), .A2(new_n964), .ZN(G66));
  INV_X1    g779(.A(KEYINPUT121), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n254), .B1(new_n331), .B2(G224), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n862), .A2(new_n868), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT120), .Z(new_n969));
  AOI211_X1 g783(.A(new_n966), .B(new_n967), .C1(new_n969), .C2(new_n254), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n966), .B2(new_n967), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n899), .B1(G898), .B2(new_n254), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n971), .B(new_n973), .ZN(G69));
  NAND2_X1  g788(.A1(new_n448), .A2(new_n449), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(new_n310), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n795), .B1(new_n775), .B2(new_n788), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n665), .A2(new_n667), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT40), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n980), .A2(new_n558), .A3(new_n681), .A4(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n687), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n659), .A2(new_n822), .A3(new_n742), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n978), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n688), .A2(KEYINPUT62), .A3(new_n659), .A4(new_n828), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n487), .B1(new_n858), .B2(new_n618), .ZN(new_n989));
  OR3_X1    g803(.A1(new_n989), .A2(new_n979), .A3(new_n744), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n977), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT123), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT123), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n977), .A2(new_n988), .A3(new_n993), .A4(new_n990), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n976), .B1(new_n995), .B2(new_n254), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT124), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n819), .A2(new_n882), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(new_n786), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n835), .A2(new_n985), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n977), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(KEYINPUT126), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n977), .A2(new_n1004), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1005));
  AOI21_X1  g819(.A(G953), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n254), .A2(G900), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n976), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT124), .ZN(new_n1009));
  AOI21_X1  g823(.A(G953), .B1(new_n992), .B2(new_n994), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n976), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n997), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n254), .B1(G227), .B2(G900), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT125), .Z(new_n1014));
  XNOR2_X1  g828(.A(new_n1012), .B(new_n1014), .ZN(G72));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  NAND2_X1  g831(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1017), .B1(new_n1018), .B2(new_n969), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n914), .B1(new_n1019), .B2(new_n451), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1017), .B1(new_n995), .B2(new_n969), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n673), .ZN(new_n1022));
  INV_X1    g836(.A(new_n673), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1023), .A2(new_n468), .A3(new_n1017), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n867), .B(new_n1024), .C1(new_n833), .C2(new_n880), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1020), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(KEYINPUT127), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT127), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1020), .A2(new_n1028), .A3(new_n1022), .A4(new_n1025), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(G57));
endmodule


