

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U321 ( .A(n319), .B(KEYINPUT8), .ZN(n320) );
  XOR2_X1 U322 ( .A(n546), .B(KEYINPUT28), .Z(n511) );
  XOR2_X1 U323 ( .A(KEYINPUT62), .B(n584), .Z(n289) );
  XOR2_X1 U324 ( .A(G218GAT), .B(KEYINPUT10), .Z(n290) );
  XNOR2_X1 U325 ( .A(n422), .B(n290), .ZN(n423) );
  XNOR2_X1 U326 ( .A(n321), .B(n320), .ZN(n415) );
  XOR2_X1 U327 ( .A(KEYINPUT123), .B(n568), .Z(n581) );
  XNOR2_X1 U328 ( .A(n424), .B(n423), .ZN(n537) );
  XOR2_X1 U329 ( .A(n382), .B(n381), .Z(n487) );
  XOR2_X1 U330 ( .A(G57GAT), .B(G148GAT), .Z(n292) );
  XNOR2_X1 U331 ( .A(G1GAT), .B(G120GAT), .ZN(n291) );
  XNOR2_X1 U332 ( .A(n292), .B(n291), .ZN(n308) );
  XOR2_X1 U333 ( .A(G85GAT), .B(G162GAT), .Z(n294) );
  XNOR2_X1 U334 ( .A(G29GAT), .B(G141GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n299) );
  XNOR2_X1 U336 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n295), .B(KEYINPUT3), .ZN(n353) );
  XOR2_X1 U338 ( .A(n353), .B(KEYINPUT94), .Z(n297) );
  NAND2_X1 U339 ( .A1(G225GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U341 ( .A(n299), .B(n298), .Z(n306) );
  XOR2_X1 U342 ( .A(G127GAT), .B(KEYINPUT0), .Z(n301) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(G134GAT), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n373) );
  XOR2_X1 U345 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n303) );
  XNOR2_X1 U346 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U348 ( .A(n373), .B(n304), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U350 ( .A(n308), .B(n307), .Z(n544) );
  INV_X1 U351 ( .A(n544), .ZN(n564) );
  XOR2_X1 U352 ( .A(G113GAT), .B(G197GAT), .Z(n310) );
  XOR2_X1 U353 ( .A(G169GAT), .B(G8GAT), .Z(n384) );
  XOR2_X1 U354 ( .A(G15GAT), .B(G1GAT), .Z(n426) );
  XNOR2_X1 U355 ( .A(n384), .B(n426), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U357 ( .A(G141GAT), .B(G22GAT), .Z(n361) );
  XOR2_X1 U358 ( .A(n311), .B(n361), .Z(n316) );
  XOR2_X1 U359 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n313) );
  NAND2_X1 U360 ( .A1(G229GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U362 ( .A(KEYINPUT72), .B(n314), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n326) );
  XOR2_X1 U364 ( .A(G43GAT), .B(G29GAT), .Z(n318) );
  XNOR2_X1 U365 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n321) );
  XOR2_X1 U367 ( .A(G36GAT), .B(KEYINPUT71), .Z(n319) );
  XOR2_X1 U368 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n323) );
  XNOR2_X1 U369 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U371 ( .A(n415), .B(n324), .Z(n325) );
  XNOR2_X1 U372 ( .A(n326), .B(n325), .ZN(n569) );
  XOR2_X1 U373 ( .A(KEYINPUT73), .B(n569), .Z(n504) );
  INV_X1 U374 ( .A(n504), .ZN(n551) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n359) );
  XNOR2_X1 U378 ( .A(G176GAT), .B(G92GAT), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n329), .B(G64GAT), .ZN(n383) );
  XNOR2_X1 U380 ( .A(n359), .B(n383), .ZN(n342) );
  XOR2_X1 U381 ( .A(G99GAT), .B(G85GAT), .Z(n418) );
  XOR2_X1 U382 ( .A(G57GAT), .B(KEYINPUT13), .Z(n425) );
  XOR2_X1 U383 ( .A(n418), .B(n425), .Z(n331) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U386 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n333) );
  XNOR2_X1 U387 ( .A(KEYINPUT76), .B(KEYINPUT78), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U389 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U390 ( .A(G120GAT), .B(G71GAT), .Z(n369) );
  XOR2_X1 U391 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n337) );
  XNOR2_X1 U392 ( .A(G204GAT), .B(KEYINPUT32), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n369), .B(n338), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n573) );
  NOR2_X1 U397 ( .A1(n551), .A2(n573), .ZN(n460) );
  XOR2_X1 U398 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n344) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(KEYINPUT92), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U401 ( .A(KEYINPUT93), .B(KEYINPUT88), .Z(n346) );
  XNOR2_X1 U402 ( .A(KEYINPUT91), .B(KEYINPUT89), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U404 ( .A(n348), .B(n347), .Z(n358) );
  XNOR2_X1 U405 ( .A(G211GAT), .B(G218GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n349), .B(KEYINPUT21), .ZN(n350) );
  XOR2_X1 U407 ( .A(n350), .B(KEYINPUT90), .Z(n352) );
  XNOR2_X1 U408 ( .A(G197GAT), .B(G204GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n390) );
  XOR2_X1 U410 ( .A(n353), .B(KEYINPUT22), .Z(n355) );
  NAND2_X1 U411 ( .A1(G228GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n390), .B(n356), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n360) );
  XOR2_X1 U415 ( .A(n360), .B(n359), .Z(n363) );
  XOR2_X1 U416 ( .A(KEYINPUT79), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U417 ( .A(n361), .B(n419), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n546) );
  XOR2_X1 U419 ( .A(KEYINPUT85), .B(G176GAT), .Z(n365) );
  XNOR2_X1 U420 ( .A(G169GAT), .B(G15GAT), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n377) );
  XOR2_X1 U422 ( .A(KEYINPUT64), .B(G99GAT), .Z(n367) );
  XNOR2_X1 U423 ( .A(G43GAT), .B(G190GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U425 ( .A(n369), .B(n368), .Z(n371) );
  NAND2_X1 U426 ( .A1(G227GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U428 ( .A(n372), .B(KEYINPUT87), .Z(n375) );
  XNOR2_X1 U429 ( .A(n373), .B(KEYINPUT20), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n377), .B(n376), .ZN(n382) );
  XOR2_X1 U432 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n379) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U435 ( .A(KEYINPUT19), .B(n380), .Z(n394) );
  INV_X1 U436 ( .A(n394), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U438 ( .A(G190GAT), .B(KEYINPUT81), .Z(n408) );
  XNOR2_X1 U439 ( .A(n385), .B(n408), .ZN(n389) );
  XOR2_X1 U440 ( .A(KEYINPUT82), .B(KEYINPUT95), .Z(n387) );
  NAND2_X1 U441 ( .A1(G226GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U443 ( .A(n389), .B(n388), .Z(n392) );
  XNOR2_X1 U444 ( .A(G36GAT), .B(n390), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U446 ( .A(n394), .B(n393), .Z(n449) );
  INV_X1 U447 ( .A(n449), .ZN(n541) );
  NOR2_X1 U448 ( .A1(n487), .A2(n541), .ZN(n395) );
  NOR2_X1 U449 ( .A1(n546), .A2(n395), .ZN(n396) );
  XOR2_X1 U450 ( .A(KEYINPUT25), .B(n396), .Z(n400) );
  XOR2_X1 U451 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n398) );
  NAND2_X1 U452 ( .A1(n546), .A2(n487), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n398), .B(n397), .ZN(n565) );
  XNOR2_X1 U454 ( .A(KEYINPUT27), .B(n541), .ZN(n402) );
  NOR2_X1 U455 ( .A1(n565), .A2(n402), .ZN(n399) );
  NOR2_X1 U456 ( .A1(n400), .A2(n399), .ZN(n401) );
  NOR2_X1 U457 ( .A1(n564), .A2(n401), .ZN(n406) );
  NOR2_X1 U458 ( .A1(n544), .A2(n402), .ZN(n403) );
  XOR2_X1 U459 ( .A(KEYINPUT96), .B(n403), .Z(n509) );
  NAND2_X1 U460 ( .A1(n487), .A2(n511), .ZN(n404) );
  NOR2_X1 U461 ( .A1(n509), .A2(n404), .ZN(n405) );
  NOR2_X1 U462 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U463 ( .A(KEYINPUT98), .B(n407), .ZN(n457) );
  XOR2_X1 U464 ( .A(G92GAT), .B(n408), .Z(n410) );
  NAND2_X1 U465 ( .A1(G232GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U467 ( .A(KEYINPUT65), .B(KEYINPUT80), .Z(n412) );
  XNOR2_X1 U468 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n417) );
  XNOR2_X1 U471 ( .A(n415), .B(G106GAT), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n424) );
  XOR2_X1 U473 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n421) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U476 ( .A(n425), .B(G78GAT), .Z(n428) );
  XNOR2_X1 U477 ( .A(n426), .B(G155GAT), .ZN(n427) );
  XNOR2_X1 U478 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U479 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n430) );
  XNOR2_X1 U480 ( .A(G64GAT), .B(KEYINPUT83), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U482 ( .A(n432), .B(n431), .Z(n434) );
  XNOR2_X1 U483 ( .A(G22GAT), .B(G211GAT), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U485 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n436) );
  NAND2_X1 U486 ( .A1(G231GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U488 ( .A(n438), .B(n437), .Z(n443) );
  XOR2_X1 U489 ( .A(G71GAT), .B(G127GAT), .Z(n440) );
  XNOR2_X1 U490 ( .A(G8GAT), .B(G183GAT), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U492 ( .A(n441), .B(KEYINPUT12), .ZN(n442) );
  XNOR2_X1 U493 ( .A(n443), .B(n442), .ZN(n577) );
  INV_X1 U494 ( .A(n577), .ZN(n558) );
  NOR2_X1 U495 ( .A1(n537), .A2(n558), .ZN(n444) );
  XOR2_X1 U496 ( .A(KEYINPUT16), .B(n444), .Z(n445) );
  NOR2_X1 U497 ( .A1(n457), .A2(n445), .ZN(n472) );
  NAND2_X1 U498 ( .A1(n460), .A2(n472), .ZN(n446) );
  XNOR2_X1 U499 ( .A(KEYINPUT99), .B(n446), .ZN(n454) );
  NAND2_X1 U500 ( .A1(n564), .A2(n454), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n447), .B(KEYINPUT34), .ZN(n448) );
  XNOR2_X1 U502 ( .A(G1GAT), .B(n448), .ZN(G1324GAT) );
  NAND2_X1 U503 ( .A1(n449), .A2(n454), .ZN(n450) );
  XNOR2_X1 U504 ( .A(G8GAT), .B(n450), .ZN(G1325GAT) );
  XOR2_X1 U505 ( .A(G15GAT), .B(KEYINPUT35), .Z(n452) );
  INV_X1 U506 ( .A(n487), .ZN(n549) );
  NAND2_X1 U507 ( .A1(n454), .A2(n549), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(G1326GAT) );
  XNOR2_X1 U509 ( .A(G22GAT), .B(KEYINPUT100), .ZN(n456) );
  INV_X1 U510 ( .A(n511), .ZN(n453) );
  NAND2_X1 U511 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n456), .B(n455), .ZN(G1327GAT) );
  XNOR2_X1 U513 ( .A(KEYINPUT101), .B(KEYINPUT39), .ZN(n463) );
  INV_X1 U514 ( .A(n537), .ZN(n561) );
  XNOR2_X1 U515 ( .A(n561), .B(KEYINPUT36), .ZN(n583) );
  NOR2_X1 U516 ( .A1(n583), .A2(n457), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n458), .A2(n558), .ZN(n459) );
  XNOR2_X1 U518 ( .A(KEYINPUT37), .B(n459), .ZN(n484) );
  NAND2_X1 U519 ( .A1(n460), .A2(n484), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT38), .ZN(n469) );
  NOR2_X1 U521 ( .A1(n544), .A2(n469), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U523 ( .A(G29GAT), .B(n464), .Z(G1328GAT) );
  NOR2_X1 U524 ( .A1(n469), .A2(n541), .ZN(n465) );
  XOR2_X1 U525 ( .A(G36GAT), .B(n465), .Z(G1329GAT) );
  XNOR2_X1 U526 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n487), .A2(n469), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U529 ( .A(G43GAT), .B(n468), .Z(G1330GAT) );
  XNOR2_X1 U530 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n511), .A2(n469), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(G1331GAT) );
  XOR2_X1 U533 ( .A(n573), .B(KEYINPUT41), .Z(n530) );
  INV_X1 U534 ( .A(n530), .ZN(n555) );
  NOR2_X1 U535 ( .A1(n569), .A2(n555), .ZN(n483) );
  NAND2_X1 U536 ( .A1(n472), .A2(n483), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n544), .A2(n479), .ZN(n474) );
  XNOR2_X1 U538 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n473) );
  XNOR2_X1 U539 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U540 ( .A(G57GAT), .B(n475), .Z(G1332GAT) );
  NOR2_X1 U541 ( .A1(n541), .A2(n479), .ZN(n476) );
  XOR2_X1 U542 ( .A(G64GAT), .B(n476), .Z(G1333GAT) );
  NOR2_X1 U543 ( .A1(n487), .A2(n479), .ZN(n478) );
  XNOR2_X1 U544 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n477) );
  XNOR2_X1 U545 ( .A(n478), .B(n477), .ZN(G1334GAT) );
  NOR2_X1 U546 ( .A1(n511), .A2(n479), .ZN(n481) );
  XNOR2_X1 U547 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n480) );
  XNOR2_X1 U548 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U549 ( .A(G78GAT), .B(n482), .ZN(G1335GAT) );
  NAND2_X1 U550 ( .A1(n484), .A2(n483), .ZN(n490) );
  NOR2_X1 U551 ( .A1(n544), .A2(n490), .ZN(n485) );
  XOR2_X1 U552 ( .A(G85GAT), .B(n485), .Z(G1336GAT) );
  NOR2_X1 U553 ( .A1(n541), .A2(n490), .ZN(n486) );
  XOR2_X1 U554 ( .A(G92GAT), .B(n486), .Z(G1337GAT) );
  NOR2_X1 U555 ( .A1(n487), .A2(n490), .ZN(n489) );
  XNOR2_X1 U556 ( .A(G99GAT), .B(KEYINPUT107), .ZN(n488) );
  XNOR2_X1 U557 ( .A(n489), .B(n488), .ZN(G1338GAT) );
  NOR2_X1 U558 ( .A1(n511), .A2(n490), .ZN(n491) );
  XOR2_X1 U559 ( .A(KEYINPUT44), .B(n491), .Z(n492) );
  XNOR2_X1 U560 ( .A(G106GAT), .B(n492), .ZN(G1339GAT) );
  INV_X1 U561 ( .A(n569), .ZN(n493) );
  NOR2_X1 U562 ( .A1(n493), .A2(n555), .ZN(n495) );
  XNOR2_X1 U563 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n494) );
  XNOR2_X1 U564 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U565 ( .A(n496), .B(KEYINPUT108), .ZN(n498) );
  NOR2_X1 U566 ( .A1(n537), .A2(n577), .ZN(n497) );
  NAND2_X1 U567 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U568 ( .A(n499), .B(KEYINPUT47), .ZN(n507) );
  NOR2_X1 U569 ( .A1(n583), .A2(n558), .ZN(n500) );
  XNOR2_X1 U570 ( .A(n500), .B(KEYINPUT45), .ZN(n502) );
  INV_X1 U571 ( .A(n573), .ZN(n501) );
  NAND2_X1 U572 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U573 ( .A(n503), .B(KEYINPUT110), .ZN(n505) );
  NOR2_X1 U574 ( .A1(n505), .A2(n504), .ZN(n506) );
  NOR2_X1 U575 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n508), .B(KEYINPUT48), .ZN(n542) );
  NOR2_X1 U577 ( .A1(n509), .A2(n542), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n525), .A2(n549), .ZN(n510) );
  XNOR2_X1 U579 ( .A(KEYINPUT111), .B(n510), .ZN(n512) );
  NAND2_X1 U580 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U581 ( .A(KEYINPUT112), .B(n513), .ZN(n521) );
  NOR2_X1 U582 ( .A1(n551), .A2(n521), .ZN(n514) );
  XNOR2_X1 U583 ( .A(G113GAT), .B(n514), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n515), .B(KEYINPUT113), .ZN(G1340GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n555), .ZN(n517) );
  XNOR2_X1 U586 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n516) );
  XNOR2_X1 U587 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U588 ( .A(G120GAT), .B(n518), .ZN(G1341GAT) );
  NOR2_X1 U589 ( .A1(n521), .A2(n558), .ZN(n519) );
  XOR2_X1 U590 ( .A(KEYINPUT50), .B(n519), .Z(n520) );
  XNOR2_X1 U591 ( .A(G127GAT), .B(n520), .ZN(G1342GAT) );
  NOR2_X1 U592 ( .A1(n521), .A2(n561), .ZN(n523) );
  XNOR2_X1 U593 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n522) );
  XNOR2_X1 U594 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U595 ( .A(G134GAT), .B(n524), .Z(G1343GAT) );
  XOR2_X1 U596 ( .A(G141GAT), .B(KEYINPUT117), .Z(n529) );
  INV_X1 U597 ( .A(n565), .ZN(n526) );
  NAND2_X1 U598 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(n527), .Z(n538) );
  NAND2_X1 U600 ( .A1(n538), .A2(n569), .ZN(n528) );
  XNOR2_X1 U601 ( .A(n529), .B(n528), .ZN(G1344GAT) );
  XNOR2_X1 U602 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n534) );
  XOR2_X1 U603 ( .A(G148GAT), .B(KEYINPUT118), .Z(n532) );
  NAND2_X1 U604 ( .A1(n530), .A2(n538), .ZN(n531) );
  XNOR2_X1 U605 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U606 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  XOR2_X1 U607 ( .A(G155GAT), .B(KEYINPUT119), .Z(n536) );
  NAND2_X1 U608 ( .A1(n577), .A2(n538), .ZN(n535) );
  XNOR2_X1 U609 ( .A(n536), .B(n535), .ZN(G1346GAT) );
  NAND2_X1 U610 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U611 ( .A(n539), .B(KEYINPUT120), .ZN(n540) );
  XNOR2_X1 U612 ( .A(G162GAT), .B(n540), .ZN(G1347GAT) );
  NOR2_X1 U613 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n543), .B(KEYINPUT54), .ZN(n567) );
  NAND2_X1 U615 ( .A1(n567), .A2(n544), .ZN(n545) );
  NOR2_X1 U616 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U617 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n547) );
  XNOR2_X1 U618 ( .A(n548), .B(n547), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n560) );
  NOR2_X1 U620 ( .A1(n551), .A2(n560), .ZN(n552) );
  XOR2_X1 U621 ( .A(G169GAT), .B(n552), .Z(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n554) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n553) );
  XNOR2_X1 U624 ( .A(n554), .B(n553), .ZN(n557) );
  NOR2_X1 U625 ( .A1(n555), .A2(n560), .ZN(n556) );
  XOR2_X1 U626 ( .A(n557), .B(n556), .Z(G1349GAT) );
  NOR2_X1 U627 ( .A1(n558), .A2(n560), .ZN(n559) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n559), .Z(G1350GAT) );
  NOR2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U630 ( .A(KEYINPUT58), .B(n562), .Z(n563) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NOR2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U635 ( .A1(n581), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n579) );
  NAND2_X1 U643 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  INV_X1 U646 ( .A(n581), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n289), .ZN(G1355GAT) );
endmodule

