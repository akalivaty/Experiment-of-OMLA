//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n205), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT64), .Z(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n208), .B(new_n222), .C1(new_n225), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G68), .Z(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G274), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  OAI211_X1 g0052(.A(G1), .B(G13), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n248), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n250), .B1(new_n254), .B2(new_n211), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G222), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n258), .B1(new_n202), .B2(new_n256), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G190), .ZN(new_n264));
  INV_X1    g0064(.A(new_n263), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G200), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT10), .ZN(new_n269));
  INV_X1    g0069(.A(G200), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n269), .B1(new_n271), .B2(KEYINPUT70), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n223), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n224), .A2(G33), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT67), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT8), .B(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT66), .ZN(new_n279));
  XOR2_X1   g0079(.A(KEYINPUT8), .B(G58), .Z(new_n280));
  INV_X1    g0080(.A(KEYINPUT66), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n277), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n284), .A2(new_n286), .B1(new_n201), .B2(new_n224), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n275), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n275), .B1(new_n247), .B2(G20), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(G50), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(KEYINPUT9), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT9), .B1(new_n288), .B2(new_n292), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT69), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n295), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT69), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n273), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT71), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n273), .A2(new_n300), .A3(KEYINPUT71), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n297), .A2(new_n293), .A3(new_n266), .A4(new_n264), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n303), .A2(new_n304), .B1(KEYINPUT10), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n288), .A2(new_n292), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G169), .B2(new_n263), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n265), .A2(G179), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n277), .A2(new_n202), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n286), .A2(new_n210), .B1(new_n224), .B2(G68), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n275), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n314), .A2(KEYINPUT11), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(KEYINPUT11), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT72), .B1(new_n289), .B2(G68), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT12), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n291), .A2(G68), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G33), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n323), .A2(new_n325), .A3(G232), .A4(G1698), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n323), .A2(new_n325), .A3(G226), .A4(new_n257), .ZN(new_n327));
  INV_X1    g0127(.A(G97), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n327), .C1(new_n251), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n262), .ZN(new_n330));
  INV_X1    g0130(.A(G274), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n248), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n254), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(G238), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT13), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT13), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(G179), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n336), .B2(new_n338), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n338), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n337), .B1(new_n330), .B2(new_n334), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n342), .B(G169), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n322), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(G200), .B1(new_n344), .B2(new_n345), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n336), .A2(G190), .A3(new_n338), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n317), .A2(new_n321), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n323), .A2(new_n325), .A3(G226), .A4(G1698), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n323), .A2(new_n325), .A3(G223), .A4(new_n257), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G87), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n262), .ZN(new_n357));
  INV_X1    g0157(.A(G179), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n253), .A2(G232), .A3(new_n248), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n359), .A2(new_n250), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n250), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n262), .B2(new_n356), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n363), .B2(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n323), .A2(new_n325), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT7), .B1(new_n365), .B2(new_n224), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  AOI211_X1 g0167(.A(new_n367), .B(G20), .C1(new_n323), .C2(new_n325), .ZN(new_n368));
  OAI21_X1  g0168(.A(G68), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n216), .A2(new_n218), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G58), .A2(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n285), .A2(G159), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT16), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n367), .B1(new_n256), .B2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n365), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n218), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n377), .B1(new_n380), .B2(new_n374), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(new_n381), .A3(new_n275), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n282), .A2(new_n279), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n291), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n383), .B2(new_n289), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n364), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G190), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n357), .A2(new_n390), .A3(new_n360), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n363), .B2(G200), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n382), .A2(new_n386), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT17), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n291), .A2(G77), .ZN(new_n396));
  INV_X1    g0196(.A(new_n289), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n202), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n280), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n400));
  XOR2_X1   g0200(.A(KEYINPUT15), .B(G87), .Z(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n276), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n399), .B1(new_n403), .B2(new_n275), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n365), .A2(G107), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n259), .B2(new_n219), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n365), .A2(new_n217), .A3(G1698), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n262), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT68), .ZN(new_n409));
  INV_X1    g0209(.A(G244), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n250), .B(new_n409), .C1(new_n254), .C2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n250), .B1(new_n254), .B2(new_n410), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT68), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n404), .B1(new_n340), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n413), .A2(new_n411), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(new_n358), .A3(new_n408), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(G190), .A3(new_n408), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(G200), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n404), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n352), .A2(new_n389), .A3(new_n395), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n311), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n323), .A2(new_n325), .A3(G257), .A4(new_n257), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n323), .A2(new_n325), .A3(G264), .A4(G1698), .ZN(new_n426));
  INV_X1    g0226(.A(G303), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n425), .B(new_n426), .C1(new_n427), .C2(new_n256), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n262), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT5), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT77), .B1(new_n430), .B2(G41), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT77), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(new_n252), .A3(KEYINPUT5), .ZN(new_n433));
  INV_X1    g0233(.A(G45), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(G1), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(G41), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n431), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n437), .A2(new_n331), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(G270), .A3(new_n253), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n429), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G200), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n251), .A2(KEYINPUT74), .A3(G1), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n397), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n275), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT74), .B1(new_n251), .B2(G1), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n443), .A2(G116), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G116), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n397), .A2(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n274), .A2(new_n223), .B1(G20), .B2(new_n447), .ZN(new_n449));
  AOI21_X1  g0249(.A(G20), .B1(G33), .B2(G283), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(G33), .B2(new_n328), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT20), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT20), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n446), .B(new_n448), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n441), .B(new_n455), .C1(new_n390), .C2(new_n440), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n440), .A2(new_n454), .A3(G169), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT21), .ZN(new_n459));
  AND4_X1   g0259(.A1(G179), .A2(new_n429), .A3(new_n438), .A4(new_n439), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n458), .A2(new_n459), .B1(new_n460), .B2(new_n454), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n437), .A2(new_n331), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n437), .A2(new_n253), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(G270), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n340), .B1(new_n465), .B2(new_n429), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT78), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT21), .A4(new_n454), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT78), .B1(new_n458), .B2(new_n459), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n461), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n457), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n323), .A2(new_n325), .A3(G244), .A4(new_n257), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n323), .A2(new_n325), .A3(G250), .A4(G1698), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT76), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n256), .A2(KEYINPUT76), .A3(G250), .A4(G1698), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n475), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G283), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n251), .A2(new_n481), .B1(KEYINPUT75), .B2(KEYINPUT4), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n473), .B2(new_n474), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n262), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n462), .B1(new_n464), .B2(G257), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n340), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n358), .A3(new_n486), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n289), .A2(G97), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n328), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G107), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n378), .B2(new_n379), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n328), .A2(G107), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT73), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT6), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(KEYINPUT73), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n497), .B(new_n498), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n328), .A2(G107), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(KEYINPUT73), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n224), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n286), .A2(new_n202), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n496), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n494), .B1(new_n510), .B2(new_n444), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n488), .A2(new_n489), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n497), .A2(new_n498), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT73), .B(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n509), .B1(new_n515), .B2(G20), .ZN(new_n516));
  OAI21_X1  g0316(.A(G107), .B1(new_n366), .B2(new_n368), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n493), .B1(new_n518), .B2(new_n275), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n485), .A2(G190), .A3(new_n486), .ZN(new_n520));
  INV_X1    g0320(.A(G257), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n438), .B1(new_n521), .B2(new_n463), .ZN(new_n522));
  INV_X1    g0322(.A(new_n484), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(new_n475), .A3(new_n478), .A4(new_n479), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n522), .B1(new_n524), .B2(new_n262), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n519), .B(new_n520), .C1(new_n525), .C2(new_n270), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n495), .A2(KEYINPUT23), .A3(G20), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT23), .B1(new_n495), .B2(G20), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G116), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n527), .A2(new_n528), .B1(G20), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n323), .A2(new_n325), .A3(new_n224), .A4(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT22), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT22), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n256), .A2(new_n533), .A3(new_n224), .A4(G87), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n535), .A2(KEYINPUT24), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(KEYINPUT24), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n275), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n256), .A2(G250), .A3(new_n257), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n256), .A2(G257), .A3(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G294), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n262), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n437), .A2(G264), .A3(new_n253), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n438), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT25), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n289), .B2(G107), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n397), .A2(KEYINPUT25), .A3(new_n495), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n547), .A2(G107), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n543), .A2(G190), .A3(new_n438), .A4(new_n544), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n538), .A2(new_n546), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n512), .A2(new_n526), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n224), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n212), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n323), .A2(new_n325), .A3(new_n224), .A4(G68), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n276), .B2(new_n328), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n275), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n401), .A2(new_n289), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n566), .C1(new_n402), .C2(new_n492), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n435), .A2(G274), .ZN(new_n568));
  OAI21_X1  g0368(.A(G250), .B1(new_n434), .B2(G1), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n262), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n323), .A2(new_n325), .A3(G238), .A4(new_n257), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n323), .A2(new_n325), .A3(G244), .A4(G1698), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(new_n529), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n570), .B1(new_n573), .B2(new_n262), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n358), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n567), .B(new_n575), .C1(G169), .C2(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n262), .ZN(new_n577));
  INV_X1    g0377(.A(new_n570), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G200), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n443), .A2(G87), .A3(new_n444), .A4(new_n445), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n564), .A2(new_n566), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n574), .A2(G190), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n275), .B1(new_n535), .B2(KEYINPUT24), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT24), .ZN(new_n587));
  AOI211_X1 g0387(.A(new_n587), .B(new_n530), .C1(new_n532), .C2(new_n534), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n551), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n545), .A2(new_n340), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n543), .A2(new_n358), .A3(new_n438), .A4(new_n544), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  NOR4_X1   g0393(.A1(new_n424), .A2(new_n472), .A3(new_n554), .A4(new_n593), .ZN(G372));
  INV_X1    g0394(.A(new_n424), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n512), .A2(new_n526), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n461), .A2(new_n592), .A3(new_n469), .A4(new_n468), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT80), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n598), .A2(new_n564), .A3(new_n566), .A4(new_n581), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n565), .B1(new_n563), .B2(new_n275), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n598), .B1(new_n600), .B2(new_n581), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n574), .A2(G190), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n574), .A2(new_n270), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n574), .A2(G169), .ZN(new_n606));
  AOI211_X1 g0406(.A(G179), .B(new_n570), .C1(new_n573), .C2(new_n262), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n602), .A2(new_n605), .B1(new_n608), .B2(new_n567), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n596), .A2(new_n597), .A3(new_n553), .A4(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n576), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n564), .A2(new_n566), .A3(new_n581), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT80), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n600), .A2(new_n598), .A3(new_n581), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(new_n580), .A3(new_n583), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n576), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n512), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n576), .A2(new_n584), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT26), .B1(new_n512), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n610), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n595), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n624));
  INV_X1    g0424(.A(new_n304), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT71), .B1(new_n273), .B2(new_n300), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n369), .A2(new_n375), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n444), .B1(new_n628), .B2(new_n377), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n385), .B1(new_n629), .B2(new_n376), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n388), .B1(new_n630), .B2(new_n364), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n387), .A2(KEYINPUT18), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n348), .A2(new_n418), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n630), .A2(new_n394), .A3(new_n392), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n393), .A2(KEYINPUT17), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n351), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n633), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n310), .B1(new_n627), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n623), .A2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(G13), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(G20), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n247), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n455), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n472), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n470), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT81), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n649), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT82), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n589), .A2(new_n649), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n553), .A2(new_n592), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n471), .A2(new_n649), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n657), .B2(new_n650), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(G399));
  INV_X1    g0469(.A(KEYINPUT83), .ZN(new_n670));
  INV_X1    g0470(.A(new_n206), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(G41), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n206), .A2(KEYINPUT83), .A3(new_n252), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n557), .A2(new_n212), .A3(new_n447), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n675), .A2(new_n247), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n226), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n675), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT28), .Z(new_n680));
  NOR2_X1   g0480(.A1(new_n554), .A2(new_n593), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n471), .A3(new_n457), .A4(new_n650), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n429), .A2(G179), .A3(new_n438), .A4(new_n439), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT84), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n543), .A2(new_n544), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n579), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n525), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n684), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n487), .A2(new_n687), .A3(new_n579), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(KEYINPUT84), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n685), .A2(KEYINPUT84), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n691), .A2(KEYINPUT30), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n574), .A2(G179), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n487), .A2(new_n440), .A3(new_n545), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n690), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n683), .B1(new_n697), .B2(new_n649), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n682), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(new_n683), .A3(new_n649), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT26), .B1(new_n512), .B2(new_n616), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n485), .A2(new_n358), .A3(new_n486), .ZN(new_n705));
  AOI21_X1  g0505(.A(G169), .B1(new_n485), .B2(new_n486), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n706), .A3(new_n519), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(new_n585), .A3(new_n618), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n704), .A2(new_n708), .A3(new_n576), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT85), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n704), .A2(new_n708), .A3(KEYINPUT85), .A4(new_n576), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n610), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT86), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n713), .A2(new_n714), .A3(new_n650), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n713), .B2(new_n650), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT29), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n622), .A2(new_n650), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n703), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n680), .B1(new_n721), .B2(G1), .ZN(G364));
  AOI21_X1  g0522(.A(new_n247), .B1(new_n643), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n675), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n656), .B(new_n726), .C1(G330), .C2(new_n654), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n671), .A2(new_n365), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n728), .A2(G355), .B1(new_n447), .B2(new_n671), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT87), .Z(new_n730));
  NOR2_X1   g0530(.A1(new_n671), .A2(new_n256), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n245), .A2(new_n434), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT88), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n732), .B(new_n734), .C1(new_n434), .C2(new_n228), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(KEYINPUT88), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n730), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n223), .B1(G20), .B2(new_n340), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n725), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n224), .A2(new_n390), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n358), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G322), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n224), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n746), .ZN(new_n750));
  INV_X1    g0550(.A(G311), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n747), .A2(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n358), .A2(new_n270), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n745), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n256), .B1(new_n755), .B2(G326), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n270), .A2(G179), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n753), .A2(new_n749), .ZN(new_n759));
  XOR2_X1   g0559(.A(KEYINPUT33), .B(G317), .Z(new_n760));
  OAI221_X1 g0560(.A(new_n756), .B1(new_n481), .B2(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n745), .A2(new_n757), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n752), .B(new_n761), .C1(G303), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT89), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(new_n749), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT90), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT90), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G329), .ZN(new_n772));
  INV_X1    g0572(.A(G294), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n766), .A2(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n224), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n764), .B(new_n772), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n775), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G97), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT32), .B1(new_n770), .B2(new_n777), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n759), .A2(new_n218), .B1(new_n750), .B2(new_n202), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G50), .B2(new_n755), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n758), .A2(new_n495), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n256), .B1(new_n762), .B2(new_n212), .ZN(new_n785));
  INV_X1    g0585(.A(new_n747), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n784), .B(new_n785), .C1(G58), .C2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n780), .A2(new_n781), .A3(new_n783), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n776), .B1(new_n778), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT91), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n741), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n789), .B2(new_n790), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n744), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n740), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n654), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n727), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  INV_X1    g0598(.A(new_n759), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G143), .A2(new_n786), .B1(new_n799), .B2(G150), .ZN(new_n800));
  INV_X1    g0600(.A(G137), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n800), .B1(new_n801), .B2(new_n754), .C1(new_n777), .C2(new_n750), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT34), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n802), .A2(new_n803), .B1(new_n779), .B2(G58), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n256), .B1(new_n758), .B2(new_n218), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G50), .B2(new_n763), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n804), .B(new_n806), .C1(new_n803), .C2(new_n802), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n770), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n770), .A2(new_n751), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n365), .B1(new_n762), .B2(new_n495), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n747), .A2(new_n773), .B1(new_n758), .B2(new_n212), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n811), .B(new_n812), .C1(G303), .C2(new_n755), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n759), .A2(new_n481), .B1(new_n750), .B2(new_n447), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT93), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n780), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n807), .A2(new_n809), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n741), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n741), .A2(new_n738), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT92), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n726), .B1(new_n821), .B2(new_n202), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n404), .A2(new_n650), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT94), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n415), .A2(new_n824), .A3(new_n417), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n415), .B2(new_n417), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n421), .B(new_n823), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n415), .A2(new_n417), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n649), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n818), .B(new_n822), .C1(new_n830), .C2(new_n739), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n718), .A2(new_n829), .A3(new_n827), .ZN(new_n832));
  INV_X1    g0632(.A(new_n421), .ZN(new_n833));
  INV_X1    g0633(.A(new_n825), .ZN(new_n834));
  INV_X1    g0634(.A(new_n826), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND4_X1   g0636(.A1(new_n468), .A2(new_n461), .A3(new_n469), .A4(new_n592), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n609), .A2(new_n553), .A3(new_n512), .A4(new_n526), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n609), .A2(new_n707), .A3(new_n618), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(new_n621), .A3(new_n576), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n650), .B(new_n836), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT95), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n622), .A2(KEYINPUT95), .A3(new_n650), .A4(new_n836), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n703), .B1(new_n832), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT98), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n703), .A2(new_n832), .A3(new_n846), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n725), .B1(new_n849), .B2(KEYINPUT96), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(KEYINPUT96), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n848), .B1(new_n851), .B2(KEYINPUT97), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n851), .A2(KEYINPUT97), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n831), .B1(new_n852), .B2(new_n853), .ZN(G384));
  OAI21_X1  g0654(.A(G77), .B1(new_n216), .B2(new_n218), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n855), .A2(new_n226), .B1(G50), .B2(new_n218), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(G1), .A3(new_n642), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(G116), .A3(new_n225), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(KEYINPUT35), .B2(new_n515), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n857), .B1(new_n860), .B2(KEYINPUT36), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(KEYINPUT36), .B2(new_n860), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n863), .B(new_n393), .C1(new_n630), .C2(new_n647), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT99), .B1(new_n630), .B2(new_n364), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT99), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n387), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n864), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n382), .A2(new_n386), .A3(new_n392), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n387), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n382), .A2(new_n386), .ZN(new_n871));
  INV_X1    g0671(.A(new_n647), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n863), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT100), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n393), .A2(new_n863), .ZN(new_n876));
  AOI211_X1 g0676(.A(KEYINPUT99), .B(new_n364), .C1(new_n382), .C2(new_n386), .ZN(new_n877));
  INV_X1    g0677(.A(new_n364), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n866), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n876), .B(new_n873), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n871), .A2(new_n878), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n873), .A3(new_n393), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT100), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n647), .B1(new_n382), .B2(new_n386), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n389), .B2(new_n395), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n885), .A4(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n873), .B1(new_n633), .B2(new_n637), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n880), .A2(new_n883), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(KEYINPUT100), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(KEYINPUT102), .A3(KEYINPUT38), .A4(new_n885), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n873), .B1(new_n870), .B2(KEYINPUT101), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n881), .A2(KEYINPUT101), .A3(new_n393), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT37), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n880), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n900), .B2(new_n887), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n895), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n865), .A2(new_n867), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n869), .A2(new_n886), .A3(KEYINPUT37), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n905), .A2(new_n906), .B1(new_n882), .B2(KEYINPUT37), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n887), .B1(new_n907), .B2(new_n884), .ZN(new_n908));
  INV_X1    g0708(.A(new_n885), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n888), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT39), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n348), .A2(new_n649), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n825), .A2(new_n826), .A3(new_n649), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n844), .B2(new_n845), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n322), .A2(new_n649), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n348), .A2(new_n351), .A3(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n322), .B(new_n649), .C1(new_n343), .C2(new_n347), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n918), .A2(new_n911), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n633), .A2(new_n872), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n915), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n717), .A2(new_n595), .A3(new_n720), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n640), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n927), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n595), .A2(new_n703), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n901), .B1(new_n890), .B2(new_n894), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n920), .A2(new_n921), .B1(new_n827), .B2(new_n829), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n699), .A2(new_n933), .A3(new_n700), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT40), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n934), .B1(new_n910), .B2(new_n888), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n932), .A2(new_n936), .B1(new_n937), .B2(KEYINPUT40), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n931), .B1(new_n938), .B2(new_n702), .ZN(new_n939));
  INV_X1    g0739(.A(new_n701), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n595), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n939), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n930), .A2(new_n942), .B1(new_n247), .B2(new_n643), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n943), .A2(KEYINPUT103), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n930), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n943), .B2(KEYINPUT103), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n862), .B1(new_n944), .B2(new_n946), .ZN(G367));
  AOI21_X1  g0747(.A(KEYINPUT46), .B1(new_n763), .B2(G116), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT109), .Z(new_n949));
  NAND3_X1  g0749(.A1(new_n763), .A2(KEYINPUT46), .A3(G116), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n365), .C1(new_n328), .C2(new_n758), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n754), .A2(new_n751), .B1(new_n750), .B2(new_n481), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n773), .A2(new_n759), .B1(new_n747), .B2(new_n427), .ZN(new_n953));
  NOR4_X1   g0753(.A1(new_n949), .A2(new_n951), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(G317), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n954), .B1(new_n495), .B2(new_n775), .C1(new_n955), .C2(new_n770), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G143), .A2(new_n755), .B1(new_n786), .B2(G150), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n775), .B2(new_n218), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(KEYINPUT110), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n771), .A2(G137), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(KEYINPUT110), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n256), .B1(new_n762), .B2(new_n216), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n759), .A2(new_n777), .B1(new_n758), .B2(new_n202), .ZN(new_n963));
  INV_X1    g0763(.A(new_n750), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n962), .B(new_n963), .C1(G50), .C2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n960), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n956), .B1(new_n959), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT47), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n792), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n968), .B2(new_n967), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n237), .A2(new_n731), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n743), .B1(new_n671), .B2(new_n401), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n726), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n609), .B1(new_n602), .B2(new_n650), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n611), .B(new_n649), .C1(new_n601), .C2(new_n599), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n970), .B(new_n973), .C1(new_n795), .C2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n596), .B1(new_n519), .B2(new_n650), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n707), .A2(new_n649), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n668), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(KEYINPUT44), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT44), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n668), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n668), .A2(new_n980), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT45), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT45), .B1(new_n668), .B2(new_n980), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n982), .A2(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n663), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n667), .A2(KEYINPUT107), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n662), .A2(new_n666), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n991), .B(new_n992), .Z(new_n993));
  INV_X1    g0793(.A(KEYINPUT108), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n656), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n993), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n721), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n721), .B1(new_n990), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n674), .B(KEYINPUT41), .Z(new_n999));
  AOI21_X1  g0799(.A(new_n724), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT105), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n1003));
  NAND3_X1  g0803(.A1(new_n974), .A2(new_n975), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n667), .A2(new_n980), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n512), .B1(new_n978), .B2(new_n592), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n650), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1002), .B1(KEYINPUT106), .B2(new_n1004), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n663), .A2(new_n980), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1004), .A2(KEYINPUT106), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n977), .B1(new_n1000), .B2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n662), .A2(new_n740), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n755), .A2(G322), .B1(new_n964), .B2(G303), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n751), .B2(new_n759), .C1(new_n955), .C2(new_n747), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n481), .B2(new_n775), .C1(new_n773), .C2(new_n762), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT49), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n365), .B1(new_n758), .B2(new_n447), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n771), .B2(G326), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G50), .A2(new_n786), .B1(new_n964), .B2(G68), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n202), .B2(new_n762), .C1(new_n777), .C2(new_n754), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n758), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n365), .B(new_n1029), .C1(G97), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n771), .A2(G150), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n779), .A2(new_n401), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n383), .A2(new_n799), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n792), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n728), .A2(new_n676), .B1(new_n495), .B2(new_n671), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n233), .A2(G45), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT111), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n278), .A2(G50), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  AOI211_X1 g0841(.A(G45), .B(new_n676), .C1(G68), .C2(G77), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n732), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT112), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1037), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n726), .B(new_n1036), .C1(new_n742), .C2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n996), .A2(new_n724), .B1(new_n1017), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n997), .A2(new_n675), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n996), .A2(new_n721), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(G393));
  OAI221_X1 g0850(.A(new_n742), .B1(new_n328), .B2(new_n206), .C1(new_n242), .C2(new_n732), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n725), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n771), .A2(G143), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n754), .A2(new_n284), .B1(new_n747), .B2(new_n777), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n779), .A2(G77), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n256), .B1(new_n758), .B2(new_n212), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n210), .A2(new_n759), .B1(new_n762), .B2(new_n218), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n280), .C2(new_n964), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n754), .A2(new_n955), .B1(new_n747), .B2(new_n751), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  OAI22_X1  g0862(.A1(new_n762), .A2(new_n481), .B1(new_n750), .B2(new_n773), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1062), .A2(new_n256), .A3(new_n784), .A4(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n775), .A2(new_n447), .B1(new_n427), .B2(new_n759), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(new_n748), .C2(new_n770), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1060), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT114), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n792), .B1(new_n1069), .B2(KEYINPUT114), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1052), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n795), .B2(new_n980), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n990), .B2(new_n723), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n990), .A2(new_n997), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(new_n674), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n990), .A2(new_n997), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G390));
  INV_X1    g0879(.A(new_n914), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n922), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n917), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n903), .A2(new_n912), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n830), .B1(new_n715), .B2(new_n716), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n916), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1081), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n895), .A2(new_n902), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n1080), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1083), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n940), .A2(G330), .A3(new_n933), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1083), .B(new_n1090), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n699), .A2(G330), .A3(new_n700), .A4(new_n830), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1081), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n917), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n713), .A2(new_n650), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT86), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n713), .A2(new_n714), .A3(new_n650), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n916), .B1(new_n1101), .B2(new_n830), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1097), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n928), .A2(new_n640), .A3(new_n931), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1094), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1092), .A2(new_n1093), .A3(new_n1106), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n675), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1092), .A2(new_n724), .A3(new_n1093), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n725), .B1(new_n820), .B2(new_n383), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n762), .A2(new_n284), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT53), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n256), .B1(new_n1113), .B2(new_n754), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT54), .B(G143), .Z(new_n1117));
  AOI22_X1  g0917(.A1(new_n964), .A2(new_n1117), .B1(new_n1030), .B2(G50), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n808), .B2(new_n747), .C1(new_n801), .C2(new_n759), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1116), .B(new_n1119), .C1(new_n1115), .C2(new_n1114), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n771), .A2(G125), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(new_n777), .C2(new_n775), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n770), .A2(new_n773), .B1(new_n218), .B2(new_n758), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(KEYINPUT117), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n365), .B1(new_n762), .B2(new_n212), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT116), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n759), .A2(new_n495), .B1(new_n750), .B2(new_n328), .ZN(new_n1127));
  OR2_X1    g0927(.A1(new_n1127), .A2(KEYINPUT115), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(KEYINPUT115), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G283), .A2(new_n755), .B1(new_n786), .B2(G116), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1126), .B(new_n1131), .C1(G77), .C2(new_n779), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1123), .A2(KEYINPUT117), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1122), .B1(new_n1124), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1112), .B1(new_n1135), .B2(new_n741), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n913), .B2(new_n739), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1110), .A2(new_n1111), .A3(new_n1137), .ZN(G378));
  INV_X1    g0938(.A(new_n1105), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1109), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1080), .B1(new_n903), .B2(new_n912), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n923), .A2(new_n925), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT40), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n934), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1087), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n911), .A2(new_n935), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1144), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n307), .A2(new_n872), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n306), .A2(new_n310), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n310), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1151), .B1(new_n627), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1150), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1152), .B1(new_n306), .B2(new_n310), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n627), .A2(new_n1154), .A3(new_n1151), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n1149), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1146), .A2(G330), .A3(new_n1148), .A4(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n938), .B2(new_n702), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1143), .A2(KEYINPUT120), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1161), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n927), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT120), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1143), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1140), .A2(new_n1164), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n674), .B1(new_n1140), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n256), .A2(G41), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G50), .B(new_n1176), .C1(new_n251), .C2(new_n252), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n251), .B(new_n252), .C1(new_n758), .C2(new_n777), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G132), .A2(new_n799), .B1(new_n763), .B2(new_n1117), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n747), .A2(new_n1113), .B1(new_n750), .B2(new_n801), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G125), .B2(new_n755), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(new_n775), .C2(new_n284), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1178), .B(new_n1184), .C1(G124), .C2(new_n771), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1177), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n758), .A2(new_n216), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G77), .B2(new_n763), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1176), .B(new_n1189), .C1(new_n770), .C2(new_n481), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT118), .Z(new_n1191));
  AOI22_X1  g0991(.A1(new_n799), .A2(G97), .B1(new_n964), .B2(new_n401), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n495), .B2(new_n747), .C1(new_n447), .C2(new_n754), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G68), .B2(new_n779), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(KEYINPUT58), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1187), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT58), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n741), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n726), .B1(new_n821), .B2(new_n210), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n1160), .C2(new_n739), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1169), .A2(new_n1164), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n724), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1175), .A2(new_n1203), .ZN(G375));
  NOR2_X1   g1004(.A1(new_n1104), .A2(new_n723), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT121), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n725), .B1(new_n820), .B2(G68), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT122), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n799), .A2(new_n1117), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n284), .B2(new_n750), .C1(new_n777), .C2(new_n762), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n754), .A2(new_n808), .B1(new_n747), .B2(new_n801), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1210), .A2(new_n365), .A3(new_n1188), .A4(new_n1211), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n210), .B2(new_n775), .C1(new_n1113), .C2(new_n770), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G97), .A2(new_n763), .B1(new_n786), .B2(G283), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n773), .B2(new_n754), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n365), .B1(new_n758), .B2(new_n202), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n759), .A2(new_n447), .B1(new_n750), .B2(new_n495), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1218), .B(new_n1033), .C1(new_n427), .C2(new_n770), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1213), .A2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1208), .B1(new_n792), .B2(new_n1220), .C1(new_n922), .C2(new_n739), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1205), .B2(KEYINPUT121), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1206), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1104), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(new_n1139), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1107), .A2(new_n999), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(G381));
  NOR3_X1   g1027(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT123), .Z(new_n1229));
  NOR2_X1   g1029(.A1(G375), .A2(G378), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(G390), .A2(G387), .A3(G381), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(G407));
  NAND3_X1  g1032(.A1(new_n1230), .A2(G213), .A3(new_n648), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1234), .A2(G213), .A3(G407), .A4(new_n1235), .ZN(G409));
  NAND2_X1  g1036(.A1(new_n648), .A2(G213), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1175), .A2(G378), .A3(new_n1203), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1165), .A2(new_n927), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1163), .A2(new_n1161), .B1(new_n915), .B2(new_n926), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n724), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1200), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1140), .A2(new_n1169), .A3(new_n999), .A4(new_n1164), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1202), .A2(KEYINPUT125), .A3(new_n999), .A4(new_n1140), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G378), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT126), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1238), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI211_X1 g1049(.A(KEYINPUT126), .B(G378), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1237), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1224), .B2(new_n1139), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1104), .A2(new_n1105), .A3(KEYINPUT60), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(new_n1107), .A3(new_n675), .A4(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1223), .A2(G384), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G384), .B1(new_n1223), .B2(new_n1255), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G2897), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1258), .A2(KEYINPUT127), .B1(new_n1259), .B2(new_n1237), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT127), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1237), .A2(new_n1259), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1258), .A2(KEYINPUT127), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1260), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1251), .B2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1237), .B(new_n1258), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(KEYINPUT62), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1269));
  INV_X1    g1069(.A(G378), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT126), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1238), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1237), .A4(new_n1258), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1266), .A2(new_n1268), .A3(new_n1276), .ZN(new_n1277));
  OR2_X1    g1077(.A1(G387), .A2(new_n1078), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(G393), .B(new_n797), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(new_n1078), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1277), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1274), .A2(KEYINPUT63), .A3(new_n1237), .A4(new_n1258), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1267), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1283), .A2(new_n1266), .A3(new_n1286), .A4(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1285), .A2(new_n1289), .ZN(G405));
  XNOR2_X1  g1090(.A(G375), .B(new_n1270), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1258), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1292), .A2(new_n1283), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1283), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(G402));
endmodule


