

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U548 ( .A1(n515), .A2(G2104), .ZN(n867) );
  NOR2_X2 U549 ( .A1(n785), .A2(n734), .ZN(n735) );
  NOR2_X2 U550 ( .A1(G164), .A2(G1384), .ZN(n758) );
  NOR2_X2 U551 ( .A1(n520), .A2(n519), .ZN(G164) );
  NAND2_X2 U552 ( .A1(n756), .A2(n758), .ZN(n711) );
  INV_X1 U553 ( .A(KEYINPUT28), .ZN(n673) );
  NOR2_X1 U554 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U555 ( .A(n521), .B(KEYINPUT23), .ZN(n522) );
  XNOR2_X1 U556 ( .A(KEYINPUT98), .B(KEYINPUT30), .ZN(n701) );
  XNOR2_X1 U557 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U558 ( .A1(G543), .A2(n535), .ZN(n536) );
  INV_X1 U559 ( .A(KEYINPUT66), .ZN(n521) );
  NOR2_X1 U560 ( .A1(n628), .A2(G651), .ZN(n638) );
  XNOR2_X1 U561 ( .A(n523), .B(n522), .ZN(n525) );
  NOR2_X1 U562 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U563 ( .A(G2105), .ZN(n515) );
  NAND2_X1 U564 ( .A1(G102), .A2(n867), .ZN(n514) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n512) );
  XOR2_X2 U566 ( .A(KEYINPUT17), .B(n512), .Z(n868) );
  NAND2_X1 U567 ( .A1(G138), .A2(n868), .ZN(n513) );
  NAND2_X1 U568 ( .A1(n514), .A2(n513), .ZN(n520) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n871) );
  NAND2_X1 U570 ( .A1(G114), .A2(n871), .ZN(n517) );
  NOR2_X2 U571 ( .A1(G2104), .A2(n515), .ZN(n872) );
  NAND2_X1 U572 ( .A1(G126), .A2(n872), .ZN(n516) );
  NAND2_X1 U573 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U574 ( .A(KEYINPUT85), .B(n518), .Z(n519) );
  NAND2_X1 U575 ( .A1(G101), .A2(n867), .ZN(n523) );
  NAND2_X1 U576 ( .A1(G137), .A2(n868), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n529) );
  NAND2_X1 U578 ( .A1(G113), .A2(n871), .ZN(n527) );
  NAND2_X1 U579 ( .A1(G125), .A2(n872), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n628) );
  INV_X1 U582 ( .A(G651), .ZN(n535) );
  NOR2_X1 U583 ( .A1(n628), .A2(n535), .ZN(n632) );
  NAND2_X1 U584 ( .A1(n632), .A2(G76), .ZN(n530) );
  XNOR2_X1 U585 ( .A(KEYINPUT76), .B(n530), .ZN(n533) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n631) );
  NAND2_X1 U587 ( .A1(n631), .A2(G89), .ZN(n531) );
  XNOR2_X1 U588 ( .A(KEYINPUT4), .B(n531), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U590 ( .A(n534), .B(KEYINPUT5), .ZN(n541) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n536), .Z(n636) );
  NAND2_X1 U592 ( .A1(G63), .A2(n636), .ZN(n538) );
  NAND2_X1 U593 ( .A1(G51), .A2(n638), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U595 ( .A(KEYINPUT6), .B(n539), .Z(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n542), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U599 ( .A1(G64), .A2(n636), .ZN(n544) );
  NAND2_X1 U600 ( .A1(G52), .A2(n638), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n549) );
  NAND2_X1 U602 ( .A1(G90), .A2(n631), .ZN(n546) );
  NAND2_X1 U603 ( .A1(G77), .A2(n632), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U606 ( .A1(n549), .A2(n548), .ZN(G171) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U608 ( .A(G132), .ZN(G219) );
  INV_X1 U609 ( .A(G82), .ZN(G220) );
  NAND2_X1 U610 ( .A1(G88), .A2(n631), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G75), .A2(n632), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G62), .A2(n636), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G50), .A2(n638), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U616 ( .A1(n555), .A2(n554), .ZN(G166) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n556), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U619 ( .A(G223), .ZN(n812) );
  NAND2_X1 U620 ( .A1(n812), .A2(G567), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  NAND2_X1 U622 ( .A1(G56), .A2(n636), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT14), .B(n558), .Z(n564) );
  NAND2_X1 U624 ( .A1(n631), .A2(G81), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U626 ( .A1(G68), .A2(n632), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT13), .B(n562), .Z(n563) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n638), .A2(G43), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n987) );
  INV_X1 U632 ( .A(G860), .ZN(n606) );
  OR2_X1 U633 ( .A1(n987), .A2(n606), .ZN(G153) );
  INV_X1 U634 ( .A(G868), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G92), .A2(n631), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n636), .A2(G66), .ZN(n567) );
  NAND2_X1 U637 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U638 ( .A(KEYINPUT74), .B(n569), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G54), .A2(n638), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G79), .A2(n632), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U642 ( .A(KEYINPUT15), .B(n574), .Z(n992) );
  NAND2_X1 U643 ( .A1(n575), .A2(n992), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G171), .A2(G868), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n578), .B(KEYINPUT75), .ZN(G284) );
  NAND2_X1 U647 ( .A1(G78), .A2(n632), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n579), .B(KEYINPUT72), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G65), .A2(n636), .ZN(n581) );
  NAND2_X1 U650 ( .A1(G53), .A2(n638), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U652 ( .A1(G91), .A2(n631), .ZN(n582) );
  XNOR2_X1 U653 ( .A(KEYINPUT71), .B(n582), .ZN(n583) );
  NOR2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(G299) );
  XNOR2_X1 U656 ( .A(KEYINPUT77), .B(G868), .ZN(n587) );
  NOR2_X1 U657 ( .A1(G286), .A2(n587), .ZN(n589) );
  NOR2_X1 U658 ( .A1(G868), .A2(G299), .ZN(n588) );
  NOR2_X1 U659 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U660 ( .A1(n606), .A2(G559), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n590), .A2(n992), .ZN(n591) );
  XNOR2_X1 U662 ( .A(n591), .B(KEYINPUT16), .ZN(n592) );
  XNOR2_X1 U663 ( .A(KEYINPUT78), .B(n592), .ZN(G148) );
  NOR2_X1 U664 ( .A1(G868), .A2(n987), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G868), .A2(n992), .ZN(n593) );
  NOR2_X1 U666 ( .A1(G559), .A2(n593), .ZN(n594) );
  NOR2_X1 U667 ( .A1(n595), .A2(n594), .ZN(G282) );
  NAND2_X1 U668 ( .A1(G123), .A2(n872), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n596), .B(KEYINPUT18), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n871), .A2(G111), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G99), .A2(n867), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G135), .A2(n868), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n909) );
  XNOR2_X1 U676 ( .A(G2096), .B(n909), .ZN(n604) );
  INV_X1 U677 ( .A(G2100), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(G156) );
  NAND2_X1 U679 ( .A1(G559), .A2(n992), .ZN(n605) );
  XOR2_X1 U680 ( .A(n987), .B(n605), .Z(n650) );
  NAND2_X1 U681 ( .A1(n606), .A2(n650), .ZN(n613) );
  NAND2_X1 U682 ( .A1(G67), .A2(n636), .ZN(n608) );
  NAND2_X1 U683 ( .A1(G93), .A2(n631), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G55), .A2(n638), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G80), .A2(n632), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n652) );
  XOR2_X1 U689 ( .A(n613), .B(n652), .Z(G145) );
  NAND2_X1 U690 ( .A1(n638), .A2(G48), .ZN(n614) );
  XNOR2_X1 U691 ( .A(KEYINPUT82), .B(n614), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n636), .A2(G61), .ZN(n615) );
  XNOR2_X1 U693 ( .A(n615), .B(KEYINPUT80), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G86), .A2(n631), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n632), .A2(G73), .ZN(n618) );
  XOR2_X1 U697 ( .A(KEYINPUT2), .B(n618), .Z(n619) );
  NOR2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U699 ( .A(KEYINPUT81), .B(n621), .Z(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(G305) );
  NAND2_X1 U701 ( .A1(G49), .A2(n638), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U704 ( .A1(n636), .A2(n626), .ZN(n627) );
  XOR2_X1 U705 ( .A(KEYINPUT79), .B(n627), .Z(n630) );
  NAND2_X1 U706 ( .A1(n628), .A2(G87), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U708 ( .A1(G85), .A2(n631), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G72), .A2(n632), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT67), .ZN(n643) );
  NAND2_X1 U712 ( .A1(n636), .A2(G60), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(KEYINPUT68), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G47), .A2(n638), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U716 ( .A(KEYINPUT69), .B(n641), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n644), .B(KEYINPUT70), .ZN(G290) );
  XNOR2_X1 U719 ( .A(G288), .B(KEYINPUT19), .ZN(n646) );
  XNOR2_X1 U720 ( .A(G290), .B(G166), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n652), .B(n647), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n648), .B(G299), .ZN(n649) );
  XNOR2_X1 U724 ( .A(G305), .B(n649), .ZN(n839) );
  XNOR2_X1 U725 ( .A(n839), .B(n650), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n651), .A2(G868), .ZN(n654) );
  OR2_X1 U727 ( .A1(G868), .A2(n652), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n654), .A2(n653), .ZN(G295) );
  NAND2_X1 U729 ( .A1(G2084), .A2(G2078), .ZN(n655) );
  XOR2_X1 U730 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U731 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U732 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n658), .A2(G2072), .ZN(n659) );
  XOR2_X1 U734 ( .A(KEYINPUT83), .B(n659), .Z(G158) );
  XNOR2_X1 U735 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U736 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  NOR2_X1 U737 ( .A1(G220), .A2(G219), .ZN(n660) );
  XNOR2_X1 U738 ( .A(KEYINPUT22), .B(n660), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n661), .A2(G96), .ZN(n662) );
  NOR2_X1 U740 ( .A1(G218), .A2(n662), .ZN(n663) );
  XOR2_X1 U741 ( .A(KEYINPUT84), .B(n663), .Z(n816) );
  NAND2_X1 U742 ( .A1(n816), .A2(G2106), .ZN(n667) );
  NAND2_X1 U743 ( .A1(G108), .A2(G120), .ZN(n664) );
  NOR2_X1 U744 ( .A1(G237), .A2(n664), .ZN(n665) );
  NAND2_X1 U745 ( .A1(G69), .A2(n665), .ZN(n817) );
  NAND2_X1 U746 ( .A1(G567), .A2(n817), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(n819) );
  NAND2_X1 U748 ( .A1(G661), .A2(G483), .ZN(n668) );
  NOR2_X1 U749 ( .A1(n819), .A2(n668), .ZN(n815) );
  NAND2_X1 U750 ( .A1(n815), .A2(G36), .ZN(G176) );
  INV_X1 U751 ( .A(G166), .ZN(G303) );
  AND2_X1 U752 ( .A1(G160), .A2(G40), .ZN(n756) );
  NAND2_X1 U753 ( .A1(G8), .A2(n711), .ZN(n785) );
  INV_X1 U754 ( .A(G299), .ZN(n990) );
  INV_X1 U755 ( .A(n711), .ZN(n695) );
  NAND2_X1 U756 ( .A1(n695), .A2(G2072), .ZN(n669) );
  XOR2_X1 U757 ( .A(KEYINPUT27), .B(n669), .Z(n671) );
  XNOR2_X1 U758 ( .A(G1956), .B(KEYINPUT94), .ZN(n937) );
  NAND2_X1 U759 ( .A1(n711), .A2(n937), .ZN(n670) );
  NAND2_X1 U760 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U761 ( .A(n672), .B(KEYINPUT95), .ZN(n688) );
  NOR2_X1 U762 ( .A1(n990), .A2(n688), .ZN(n674) );
  XNOR2_X1 U763 ( .A(n674), .B(n673), .ZN(n692) );
  INV_X1 U764 ( .A(G1996), .ZN(n837) );
  NOR2_X1 U765 ( .A1(n711), .A2(n837), .ZN(n676) );
  XNOR2_X1 U766 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n675) );
  XNOR2_X1 U767 ( .A(n676), .B(n675), .ZN(n678) );
  NAND2_X1 U768 ( .A1(n711), .A2(G1341), .ZN(n677) );
  NAND2_X1 U769 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U770 ( .A1(n987), .A2(n679), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n992), .A2(n685), .ZN(n684) );
  INV_X1 U772 ( .A(G2067), .ZN(n959) );
  NOR2_X1 U773 ( .A1(n711), .A2(n959), .ZN(n680) );
  XOR2_X1 U774 ( .A(n680), .B(KEYINPUT96), .Z(n682) );
  NAND2_X1 U775 ( .A1(n711), .A2(G1348), .ZN(n681) );
  NAND2_X1 U776 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U777 ( .A1(n684), .A2(n683), .ZN(n687) );
  OR2_X1 U778 ( .A1(n992), .A2(n685), .ZN(n686) );
  NAND2_X1 U779 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n990), .A2(n688), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n694) );
  XNOR2_X1 U783 ( .A(KEYINPUT97), .B(KEYINPUT29), .ZN(n693) );
  XNOR2_X1 U784 ( .A(n694), .B(n693), .ZN(n699) );
  XNOR2_X1 U785 ( .A(G1961), .B(KEYINPUT93), .ZN(n929) );
  NAND2_X1 U786 ( .A1(n711), .A2(n929), .ZN(n697) );
  XNOR2_X1 U787 ( .A(KEYINPUT25), .B(G2078), .ZN(n963) );
  NAND2_X1 U788 ( .A1(n695), .A2(n963), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n704) );
  NAND2_X1 U790 ( .A1(n704), .A2(G171), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n709) );
  NOR2_X1 U792 ( .A1(G1966), .A2(n785), .ZN(n725) );
  NOR2_X1 U793 ( .A1(G2084), .A2(n711), .ZN(n722) );
  NOR2_X1 U794 ( .A1(n725), .A2(n722), .ZN(n700) );
  NAND2_X1 U795 ( .A1(G8), .A2(n700), .ZN(n702) );
  NOR2_X1 U796 ( .A1(n703), .A2(G168), .ZN(n706) );
  NOR2_X1 U797 ( .A1(G171), .A2(n704), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U799 ( .A(KEYINPUT31), .B(n707), .Z(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n721) );
  NAND2_X1 U801 ( .A1(n721), .A2(G286), .ZN(n710) );
  XNOR2_X1 U802 ( .A(n710), .B(KEYINPUT100), .ZN(n718) );
  NOR2_X1 U803 ( .A1(G2090), .A2(n711), .ZN(n712) );
  XNOR2_X1 U804 ( .A(KEYINPUT101), .B(n712), .ZN(n715) );
  NOR2_X1 U805 ( .A1(G1971), .A2(n785), .ZN(n713) );
  NOR2_X1 U806 ( .A1(G166), .A2(n713), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U808 ( .A(KEYINPUT102), .B(n716), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U810 ( .A1(n719), .A2(G8), .ZN(n720) );
  XNOR2_X1 U811 ( .A(n720), .B(KEYINPUT32), .ZN(n777) );
  XOR2_X1 U812 ( .A(KEYINPUT99), .B(n721), .Z(n727) );
  NAND2_X1 U813 ( .A1(n722), .A2(G8), .ZN(n723) );
  XOR2_X1 U814 ( .A(KEYINPUT92), .B(n723), .Z(n724) );
  NOR2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n778) );
  NAND2_X1 U817 ( .A1(G1976), .A2(G288), .ZN(n985) );
  AND2_X1 U818 ( .A1(n778), .A2(n985), .ZN(n728) );
  NAND2_X1 U819 ( .A1(n777), .A2(n728), .ZN(n733) );
  INV_X1 U820 ( .A(n985), .ZN(n731) );
  NOR2_X1 U821 ( .A1(G1976), .A2(G288), .ZN(n737) );
  NOR2_X1 U822 ( .A1(G1971), .A2(G303), .ZN(n729) );
  NOR2_X1 U823 ( .A1(n737), .A2(n729), .ZN(n998) );
  XOR2_X1 U824 ( .A(n998), .B(KEYINPUT103), .Z(n730) );
  OR2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n732) );
  AND2_X1 U826 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U827 ( .A(n735), .B(KEYINPUT64), .ZN(n736) );
  OR2_X1 U828 ( .A1(KEYINPUT33), .A2(n736), .ZN(n776) );
  NAND2_X1 U829 ( .A1(n737), .A2(KEYINPUT33), .ZN(n738) );
  NOR2_X1 U830 ( .A1(n738), .A2(n785), .ZN(n740) );
  XOR2_X1 U831 ( .A(G1981), .B(G305), .Z(n999) );
  INV_X1 U832 ( .A(n999), .ZN(n739) );
  NOR2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n774) );
  NAND2_X1 U834 ( .A1(G95), .A2(n867), .ZN(n742) );
  NAND2_X1 U835 ( .A1(G131), .A2(n868), .ZN(n741) );
  NAND2_X1 U836 ( .A1(n742), .A2(n741), .ZN(n746) );
  NAND2_X1 U837 ( .A1(G107), .A2(n871), .ZN(n744) );
  NAND2_X1 U838 ( .A1(G119), .A2(n872), .ZN(n743) );
  NAND2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n745) );
  OR2_X1 U840 ( .A1(n746), .A2(n745), .ZN(n878) );
  XOR2_X1 U841 ( .A(KEYINPUT89), .B(G1991), .Z(n964) );
  AND2_X1 U842 ( .A1(n878), .A2(n964), .ZN(n755) );
  NAND2_X1 U843 ( .A1(G141), .A2(n868), .ZN(n748) );
  NAND2_X1 U844 ( .A1(G129), .A2(n872), .ZN(n747) );
  NAND2_X1 U845 ( .A1(n748), .A2(n747), .ZN(n751) );
  NAND2_X1 U846 ( .A1(n867), .A2(G105), .ZN(n749) );
  XOR2_X1 U847 ( .A(KEYINPUT38), .B(n749), .Z(n750) );
  NOR2_X1 U848 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U849 ( .A1(n871), .A2(G117), .ZN(n752) );
  NAND2_X1 U850 ( .A1(n753), .A2(n752), .ZN(n861) );
  AND2_X1 U851 ( .A1(n861), .A2(G1996), .ZN(n754) );
  NOR2_X1 U852 ( .A1(n755), .A2(n754), .ZN(n916) );
  INV_X1 U853 ( .A(n756), .ZN(n757) );
  NOR2_X1 U854 ( .A1(n758), .A2(n757), .ZN(n807) );
  INV_X1 U855 ( .A(n807), .ZN(n759) );
  NOR2_X1 U856 ( .A1(n916), .A2(n759), .ZN(n799) );
  XOR2_X1 U857 ( .A(n799), .B(KEYINPUT90), .Z(n771) );
  NAND2_X1 U858 ( .A1(n868), .A2(G140), .ZN(n760) );
  XOR2_X1 U859 ( .A(KEYINPUT87), .B(n760), .Z(n762) );
  NAND2_X1 U860 ( .A1(n867), .A2(G104), .ZN(n761) );
  NAND2_X1 U861 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U862 ( .A(KEYINPUT34), .B(n763), .ZN(n768) );
  NAND2_X1 U863 ( .A1(G116), .A2(n871), .ZN(n765) );
  NAND2_X1 U864 ( .A1(G128), .A2(n872), .ZN(n764) );
  NAND2_X1 U865 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U866 ( .A(n766), .B(KEYINPUT35), .Z(n767) );
  NOR2_X1 U867 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U868 ( .A(KEYINPUT36), .B(n769), .Z(n770) );
  XOR2_X1 U869 ( .A(KEYINPUT88), .B(n770), .Z(n882) );
  XNOR2_X1 U870 ( .A(G2067), .B(KEYINPUT37), .ZN(n796) );
  NOR2_X1 U871 ( .A1(n882), .A2(n796), .ZN(n925) );
  NAND2_X1 U872 ( .A1(n807), .A2(n925), .ZN(n804) );
  NAND2_X1 U873 ( .A1(n771), .A2(n804), .ZN(n772) );
  XOR2_X1 U874 ( .A(KEYINPUT91), .B(n772), .Z(n789) );
  INV_X1 U875 ( .A(n789), .ZN(n773) );
  AND2_X1 U876 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U877 ( .A1(n776), .A2(n775), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n777), .A2(n778), .ZN(n781) );
  NOR2_X1 U879 ( .A1(G2090), .A2(G303), .ZN(n779) );
  NAND2_X1 U880 ( .A1(G8), .A2(n779), .ZN(n780) );
  NAND2_X1 U881 ( .A1(n781), .A2(n780), .ZN(n782) );
  AND2_X1 U882 ( .A1(n782), .A2(n785), .ZN(n787) );
  NOR2_X1 U883 ( .A1(G1981), .A2(G305), .ZN(n783) );
  XOR2_X1 U884 ( .A(n783), .B(KEYINPUT24), .Z(n784) );
  NOR2_X1 U885 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U886 ( .A1(n787), .A2(n786), .ZN(n788) );
  OR2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U889 ( .A(n792), .B(KEYINPUT104), .ZN(n795) );
  XNOR2_X1 U890 ( .A(KEYINPUT86), .B(G1986), .ZN(n793) );
  XNOR2_X1 U891 ( .A(n793), .B(G290), .ZN(n1008) );
  NAND2_X1 U892 ( .A1(n1008), .A2(n807), .ZN(n794) );
  NAND2_X1 U893 ( .A1(n795), .A2(n794), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n882), .A2(n796), .ZN(n922) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n861), .ZN(n918) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n797) );
  NOR2_X1 U897 ( .A1(n964), .A2(n878), .ZN(n910) );
  NOR2_X1 U898 ( .A1(n797), .A2(n910), .ZN(n798) );
  NOR2_X1 U899 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U900 ( .A(KEYINPUT105), .B(n800), .Z(n801) );
  NOR2_X1 U901 ( .A1(n918), .A2(n801), .ZN(n802) );
  XNOR2_X1 U902 ( .A(KEYINPUT39), .B(n802), .ZN(n803) );
  XNOR2_X1 U903 ( .A(n803), .B(KEYINPUT106), .ZN(n805) );
  NAND2_X1 U904 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U905 ( .A1(n922), .A2(n806), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U908 ( .A(KEYINPUT40), .B(n811), .ZN(G329) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n812), .ZN(G217) );
  AND2_X1 U910 ( .A1(G15), .A2(G2), .ZN(n813) );
  NAND2_X1 U911 ( .A1(G661), .A2(n813), .ZN(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n815), .A2(n814), .ZN(G188) );
  XNOR2_X1 U914 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  NOR2_X1 U916 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U917 ( .A(n818), .B(KEYINPUT108), .ZN(G325) );
  XNOR2_X1 U918 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U919 ( .A(G108), .ZN(G238) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  INV_X1 U921 ( .A(G69), .ZN(G235) );
  XOR2_X1 U922 ( .A(KEYINPUT110), .B(n819), .Z(G319) );
  XOR2_X1 U923 ( .A(KEYINPUT42), .B(G2096), .Z(n821) );
  XNOR2_X1 U924 ( .A(G2100), .B(G2678), .ZN(n820) );
  XNOR2_X1 U925 ( .A(n821), .B(n820), .ZN(n825) );
  XOR2_X1 U926 ( .A(KEYINPUT43), .B(G2090), .Z(n823) );
  XNOR2_X1 U927 ( .A(G2067), .B(G2072), .ZN(n822) );
  XNOR2_X1 U928 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U929 ( .A(n825), .B(n824), .Z(n827) );
  XNOR2_X1 U930 ( .A(G2084), .B(G2078), .ZN(n826) );
  XNOR2_X1 U931 ( .A(n827), .B(n826), .ZN(G227) );
  XOR2_X1 U932 ( .A(G1991), .B(G1981), .Z(n829) );
  XNOR2_X1 U933 ( .A(G1966), .B(G1961), .ZN(n828) );
  XNOR2_X1 U934 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U935 ( .A(G1976), .B(G1971), .Z(n831) );
  XNOR2_X1 U936 ( .A(G1986), .B(G1956), .ZN(n830) );
  XNOR2_X1 U937 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U938 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U939 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n834) );
  XNOR2_X1 U940 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U941 ( .A(G2474), .B(n836), .ZN(n838) );
  XNOR2_X1 U942 ( .A(n838), .B(n837), .ZN(G229) );
  XNOR2_X1 U943 ( .A(G171), .B(n987), .ZN(n840) );
  XNOR2_X1 U944 ( .A(n840), .B(n839), .ZN(n842) );
  XNOR2_X1 U945 ( .A(G286), .B(n992), .ZN(n841) );
  XNOR2_X1 U946 ( .A(n842), .B(n841), .ZN(n843) );
  NOR2_X1 U947 ( .A1(G37), .A2(n843), .ZN(n844) );
  XOR2_X1 U948 ( .A(KEYINPUT115), .B(n844), .Z(G397) );
  NAND2_X1 U949 ( .A1(G100), .A2(n867), .ZN(n846) );
  NAND2_X1 U950 ( .A1(G112), .A2(n871), .ZN(n845) );
  NAND2_X1 U951 ( .A1(n846), .A2(n845), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G124), .A2(n872), .ZN(n847) );
  XNOR2_X1 U953 ( .A(n847), .B(KEYINPUT112), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U955 ( .A1(G136), .A2(n868), .ZN(n849) );
  NAND2_X1 U956 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U957 ( .A(KEYINPUT113), .B(n851), .Z(n852) );
  NOR2_X1 U958 ( .A1(n853), .A2(n852), .ZN(G162) );
  NAND2_X1 U959 ( .A1(G118), .A2(n871), .ZN(n855) );
  NAND2_X1 U960 ( .A1(G130), .A2(n872), .ZN(n854) );
  NAND2_X1 U961 ( .A1(n855), .A2(n854), .ZN(n860) );
  NAND2_X1 U962 ( .A1(G106), .A2(n867), .ZN(n857) );
  NAND2_X1 U963 ( .A1(G142), .A2(n868), .ZN(n856) );
  NAND2_X1 U964 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U965 ( .A(KEYINPUT45), .B(n858), .Z(n859) );
  NOR2_X1 U966 ( .A1(n860), .A2(n859), .ZN(n864) );
  XOR2_X1 U967 ( .A(n861), .B(G162), .Z(n862) );
  XNOR2_X1 U968 ( .A(n862), .B(n909), .ZN(n863) );
  XOR2_X1 U969 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U970 ( .A(G160), .B(G164), .ZN(n865) );
  XNOR2_X1 U971 ( .A(n866), .B(n865), .ZN(n884) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n880) );
  NAND2_X1 U973 ( .A1(G103), .A2(n867), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G139), .A2(n868), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G115), .A2(n871), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G127), .A2(n872), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n902) );
  XOR2_X1 U981 ( .A(n878), .B(n902), .Z(n879) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n884), .B(n883), .ZN(n885) );
  NOR2_X1 U985 ( .A1(G37), .A2(n885), .ZN(n886) );
  XNOR2_X1 U986 ( .A(KEYINPUT114), .B(n886), .ZN(G395) );
  XOR2_X1 U987 ( .A(G2451), .B(G2430), .Z(n888) );
  XNOR2_X1 U988 ( .A(G2438), .B(G2443), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n894) );
  XOR2_X1 U990 ( .A(G2435), .B(G2454), .Z(n890) );
  XNOR2_X1 U991 ( .A(G1348), .B(G1341), .ZN(n889) );
  XNOR2_X1 U992 ( .A(n890), .B(n889), .ZN(n892) );
  XOR2_X1 U993 ( .A(G2446), .B(G2427), .Z(n891) );
  XNOR2_X1 U994 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U995 ( .A(n894), .B(n893), .Z(n895) );
  NAND2_X1 U996 ( .A1(G14), .A2(n895), .ZN(n901) );
  NAND2_X1 U997 ( .A1(n901), .A2(G319), .ZN(n898) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n896) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n896), .ZN(n897) );
  NOR2_X1 U1000 ( .A1(n898), .A2(n897), .ZN(n900) );
  NOR2_X1 U1001 ( .A1(G397), .A2(G395), .ZN(n899) );
  NAND2_X1 U1002 ( .A1(n900), .A2(n899), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(G171), .ZN(G301) );
  INV_X1 U1005 ( .A(n901), .ZN(G401) );
  INV_X1 U1006 ( .A(KEYINPUT55), .ZN(n977) );
  XNOR2_X1 U1007 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(G164), .B(G2078), .ZN(n905) );
  XNOR2_X1 U1009 ( .A(G2072), .B(n902), .ZN(n903) );
  XNOR2_X1 U1010 ( .A(n903), .B(KEYINPUT116), .ZN(n904) );
  NAND2_X1 U1011 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1012 ( .A(n906), .B(KEYINPUT118), .ZN(n907) );
  XNOR2_X1 U1013 ( .A(n908), .B(n907), .ZN(n912) );
  NOR2_X1 U1014 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1015 ( .A1(n912), .A2(n911), .ZN(n914) );
  XOR2_X1 U1016 ( .A(G160), .B(G2084), .Z(n913) );
  NOR2_X1 U1017 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1018 ( .A1(n916), .A2(n915), .ZN(n921) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(KEYINPUT51), .B(n919), .ZN(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT52), .B(n926), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n977), .A2(n927), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n928), .A2(G29), .ZN(n984) );
  XNOR2_X1 U1028 ( .A(KEYINPUT123), .B(G5), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(n930), .B(n929), .ZN(n954) );
  XOR2_X1 U1030 ( .A(G1986), .B(G24), .Z(n934) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G22), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G23), .B(G1976), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(n936), .B(n935), .ZN(n952) );
  XOR2_X1 U1037 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n947) );
  XNOR2_X1 U1038 ( .A(n937), .B(G20), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(G19), .B(G1341), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1041 ( .A(G4), .B(KEYINPUT124), .Z(n941) );
  XNOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT59), .ZN(n940) );
  XNOR2_X1 U1043 ( .A(n941), .B(n940), .ZN(n943) );
  XNOR2_X1 U1044 ( .A(G1981), .B(G6), .ZN(n942) );
  NOR2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(n947), .B(n946), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(G21), .B(G1966), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(KEYINPUT126), .B(n948), .ZN(n949) );
  NOR2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1053 ( .A(KEYINPUT61), .B(n955), .Z(n956) );
  NOR2_X1 U1054 ( .A1(G16), .A2(n956), .ZN(n982) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(G34), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(n957), .B(KEYINPUT119), .ZN(n958) );
  XNOR2_X1 U1057 ( .A(G2084), .B(n958), .ZN(n975) );
  XNOR2_X1 U1058 ( .A(G2090), .B(G35), .ZN(n973) );
  XNOR2_X1 U1059 ( .A(G26), .B(n959), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n960), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(G1996), .B(G32), .ZN(n962) );
  XNOR2_X1 U1062 ( .A(G33), .B(G2072), .ZN(n961) );
  NOR2_X1 U1063 ( .A1(n962), .A2(n961), .ZN(n968) );
  XOR2_X1 U1064 ( .A(n963), .B(G27), .Z(n966) );
  XNOR2_X1 U1065 ( .A(n964), .B(G25), .ZN(n965) );
  NOR2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1069 ( .A(KEYINPUT53), .B(n971), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(n977), .B(n976), .ZN(n979) );
  INV_X1 U1073 ( .A(G29), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(G11), .A2(n980), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n1013) );
  XOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .Z(n1011) );
  XNOR2_X1 U1079 ( .A(G171), .B(G1961), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(G1341), .B(n987), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n1006) );
  XNOR2_X1 U1083 ( .A(n990), .B(G1956), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(n991), .B(KEYINPUT121), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G1348), .B(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(G1971), .A2(G303), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G168), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(KEYINPUT57), .ZN(n1002) );
  XOR2_X1 U1093 ( .A(KEYINPUT120), .B(n1002), .Z(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT122), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(n1014), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1101 ( .A(G311), .ZN(G150) );
endmodule

