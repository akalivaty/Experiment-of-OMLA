//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G228gat), .ZN(new_n204));
  INV_X1    g003(.A(G233gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n207), .B1(new_n215), .B2(KEYINPUT29), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT2), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT79), .ZN(new_n219));
  XNOR2_X1  g018(.A(G155gat), .B(G162gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT79), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n221), .A3(KEYINPUT2), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(G141gat), .A3(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(KEYINPUT76), .A2(G141gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(G148gat), .A3(new_n229), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n227), .A2(new_n230), .A3(KEYINPUT78), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT78), .B1(new_n227), .B2(new_n230), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n224), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(G141gat), .A2(G148gat), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(new_n220), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n216), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT85), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n216), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n215), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n233), .A2(new_n207), .A3(new_n238), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT29), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n206), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n206), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n230), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n227), .A2(new_n230), .A3(KEYINPUT78), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n223), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT80), .B1(new_n255), .B2(new_n237), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n257), .A3(new_n238), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n216), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n250), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G78gat), .B(G106gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT31), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n249), .B2(new_n261), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n203), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n267), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(new_n202), .A3(new_n265), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT75), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT23), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(G169gat), .B2(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n274), .B(new_n276), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(KEYINPUT25), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT24), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(G183gat), .A3(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT66), .B(G190gat), .Z(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT27), .B(G183gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(KEYINPUT28), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(KEYINPUT27), .C1(new_n295), .C2(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G183gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT27), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT68), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n290), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n293), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n273), .B1(KEYINPUT70), .B2(KEYINPUT26), .ZN(new_n303));
  AND2_X1   g102(.A1(KEYINPUT70), .A2(KEYINPUT26), .ZN(new_n304));
  OAI22_X1  g103(.A1(new_n303), .A2(new_n304), .B1(new_n279), .B2(new_n280), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT69), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n283), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n289), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT65), .B(G183gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n290), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n287), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n281), .B1(new_n313), .B2(KEYINPUT67), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n290), .A2(new_n311), .B1(new_n284), .B2(new_n286), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n310), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G226gat), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n319), .A2(KEYINPUT29), .B1(new_n320), .B2(new_n205), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n294), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n292), .ZN(new_n323));
  INV_X1    g122(.A(new_n308), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n323), .A2(new_n324), .B1(new_n288), .B2(new_n282), .ZN(new_n325));
  INV_X1    g124(.A(new_n281), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(new_n315), .B2(new_n316), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n312), .A2(new_n316), .A3(new_n287), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT25), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n320), .A2(new_n205), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n321), .A2(new_n245), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n245), .B1(new_n321), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n272), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(G64gat), .ZN(new_n338));
  INV_X1    g137(.A(G92gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n332), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n331), .B1(new_n330), .B2(new_n247), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n215), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(new_n333), .A3(KEYINPUT75), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n336), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n333), .A3(new_n340), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n352), .A2(KEYINPUT35), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(KEYINPUT35), .ZN(new_n354));
  AOI211_X1 g153(.A(new_n271), .B(new_n351), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT88), .ZN(new_n356));
  INV_X1    g155(.A(G113gat), .ZN(new_n357));
  INV_X1    g156(.A(G120gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G113gat), .A2(G120gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(KEYINPUT72), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n360), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT71), .ZN(new_n369));
  INV_X1    g168(.A(G134gat), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n369), .A2(new_n370), .A3(G127gat), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n369), .B2(new_n363), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n359), .A2(new_n362), .A3(new_n360), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n309), .B2(new_n318), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT74), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT74), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n330), .A2(new_n378), .A3(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n323), .A2(new_n324), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n364), .A2(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n380), .A2(new_n329), .A3(new_n381), .A4(new_n289), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT73), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n325), .A2(KEYINPUT73), .A3(new_n381), .A4(new_n329), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n377), .A2(new_n379), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT34), .ZN(new_n387));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n386), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT32), .B1(new_n386), .B2(new_n388), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n386), .B2(new_n388), .ZN(new_n394));
  XOR2_X1   g193(.A(G15gat), .B(G43gat), .Z(new_n395));
  XNOR2_X1  g194(.A(G71gat), .B(G99gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  OAI221_X1 g198(.A(KEYINPUT32), .B1(new_n393), .B2(new_n399), .C1(new_n386), .C2(new_n388), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n391), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n390), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n398), .A2(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n356), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n398), .A2(new_n400), .ZN(new_n406));
  INV_X1    g205(.A(new_n391), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n398), .A3(new_n400), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT88), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n375), .B1(new_n255), .B2(new_n237), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n233), .A2(new_n381), .A3(new_n238), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT81), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n420), .A3(new_n417), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n412), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT82), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n246), .A3(new_n375), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n256), .A2(KEYINPUT4), .A3(new_n381), .A4(new_n258), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n414), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n416), .A4(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n423), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n420), .B1(new_n415), .B2(new_n417), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT81), .B(new_n416), .C1(new_n413), .C2(new_n414), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT5), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AND4_X1   g232(.A1(new_n416), .A2(new_n425), .A3(new_n426), .A4(new_n428), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT82), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n425), .A2(new_n416), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n414), .A2(KEYINPUT4), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n256), .A2(new_n381), .A3(new_n258), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n438), .B1(new_n439), .B2(KEYINPUT4), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n412), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n443));
  XNOR2_X1  g242(.A(G1gat), .B(G29gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G57gat), .B(G85gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n445), .B(new_n446), .Z(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n441), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n430), .B2(new_n435), .ZN(new_n450));
  INV_X1    g249(.A(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT6), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n451), .B1(new_n436), .B2(new_n441), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(KEYINPUT6), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457));
  NOR4_X1   g256(.A1(new_n450), .A2(KEYINPUT84), .A3(new_n457), .A4(new_n451), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n453), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n355), .A2(new_n411), .A3(new_n459), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n401), .A2(new_n404), .A3(new_n271), .ZN(new_n461));
  INV_X1    g260(.A(new_n351), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT90), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT35), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n463), .B2(KEYINPUT35), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n401), .B2(new_n404), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n408), .A2(KEYINPUT36), .A3(new_n409), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n336), .A2(KEYINPUT37), .A3(new_n345), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n344), .A2(new_n333), .A3(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n475), .A2(new_n341), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT37), .B1(new_n334), .B2(new_n335), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n478), .A2(new_n472), .A3(new_n341), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n347), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(new_n453), .C1(new_n456), .C2(new_n458), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n416), .B1(new_n440), .B2(new_n425), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n447), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT39), .B1(new_n415), .B2(new_n417), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(KEYINPUT87), .Z(new_n489));
  OR2_X1    g288(.A1(new_n489), .A2(new_n483), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n487), .A2(KEYINPUT40), .A3(new_n490), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n493), .A2(new_n448), .A3(new_n494), .A4(new_n351), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n271), .B1(new_n482), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n459), .A2(new_n271), .A3(new_n462), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n471), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n467), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G8gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT93), .ZN(new_n503));
  INV_X1    g302(.A(G1gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT16), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  AND4_X1   g307(.A1(new_n501), .A2(new_n505), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n503), .A2(new_n504), .B1(new_n507), .B2(new_n502), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n501), .B1(new_n510), .B2(new_n506), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G71gat), .ZN(new_n514));
  INV_X1    g313(.A(G78gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(G71gat), .A2(G78gat), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n519));
  OAI22_X1  g318(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G57gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G64gat), .ZN(new_n522));
  INV_X1    g321(.A(G64gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G57gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n518), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n520), .B(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n513), .B1(KEYINPUT21), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G183gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n526), .A2(KEYINPUT21), .ZN(new_n529));
  XOR2_X1   g328(.A(G127gat), .B(G155gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n528), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT96), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(KEYINPUT97), .B(G211gat), .Z(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n532), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT91), .B(G29gat), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G36gat), .ZN(new_n541));
  INV_X1    g340(.A(G29gat), .ZN(new_n542));
  INV_X1    g341(.A(G36gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT14), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(G43gat), .A2(G50gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(G43gat), .A2(G50gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT15), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n553), .A3(new_n550), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n541), .A2(new_n548), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT91), .B(G29gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(new_n543), .ZN(new_n557));
  OAI211_X1 g356(.A(KEYINPUT15), .B(new_n551), .C1(new_n557), .C2(new_n547), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT17), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT92), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(new_n558), .A3(KEYINPUT17), .ZN(new_n561));
  XOR2_X1   g360(.A(G99gat), .B(G106gat), .Z(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT8), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n339), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n564), .A2(KEYINPUT99), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT99), .B1(new_n564), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n570));
  NOR2_X1   g369(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g370(.A1(G85gat), .A2(G92gat), .ZN(new_n572));
  OR3_X1    g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n562), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT8), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(G99gat), .B2(G106gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n564), .A2(KEYINPUT99), .A3(new_n566), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n562), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n587));
  INV_X1    g386(.A(new_n576), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n578), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n560), .A2(new_n561), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n555), .A2(new_n558), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n592), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n594), .B1(new_n592), .B2(new_n598), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OR3_X1    g403(.A1(new_n599), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n599), .B2(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n539), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n520), .B(new_n525), .Z(new_n610));
  AND3_X1   g409(.A1(new_n585), .A2(new_n586), .A3(new_n589), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n586), .B1(new_n585), .B2(new_n589), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n578), .A2(new_n526), .A3(new_n590), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(KEYINPUT100), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n591), .A2(new_n616), .A3(new_n610), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT10), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n609), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT102), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n623), .B(new_n609), .C1(new_n618), .C2(new_n620), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n615), .A2(new_n617), .ZN(new_n626));
  INV_X1    g425(.A(new_n609), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G204gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT101), .B(G176gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n621), .A2(new_n628), .A3(new_n633), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n608), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G229gat), .A2(G233gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n513), .A2(new_n597), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n510), .A2(new_n506), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(G8gat), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n510), .A2(new_n501), .A3(new_n506), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT94), .B1(new_n509), .B2(new_n511), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n561), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n559), .A2(KEYINPUT92), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT92), .ZN(new_n649));
  AOI211_X1 g448(.A(new_n649), .B(KEYINPUT17), .C1(new_n555), .C2(new_n558), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n639), .B(new_n640), .C1(new_n647), .C2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n561), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(new_n512), .B2(new_n643), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n560), .A2(new_n656), .A3(new_n646), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n657), .A2(KEYINPUT18), .A3(new_n639), .A4(new_n640), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n512), .B(new_n597), .Z(new_n659));
  XOR2_X1   g458(.A(new_n639), .B(KEYINPUT13), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n654), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G113gat), .B(G141gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT11), .ZN(new_n664));
  INV_X1    g463(.A(G169gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G197gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT12), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n668), .A2(new_n654), .A3(new_n658), .A4(new_n661), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n638), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n500), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n459), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n504), .ZN(G1324gat));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678));
  INV_X1    g477(.A(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n351), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT16), .B(G8gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(G8gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(new_n411), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n675), .A2(G15gat), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT104), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT104), .B1(new_n469), .B2(new_n470), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G15gat), .B1(new_n675), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n688), .A2(new_n693), .ZN(G1326gat));
  INV_X1    g493(.A(new_n271), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n675), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT43), .B(G22gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n607), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n467), .B2(new_n499), .ZN(new_n700));
  INV_X1    g499(.A(new_n539), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n635), .A2(new_n636), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(new_n673), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(new_n459), .A3(new_n540), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT45), .Z(new_n706));
  OAI21_X1  g505(.A(new_n692), .B1(new_n496), .B2(new_n498), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n467), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n607), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n700), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n703), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n540), .B1(new_n713), .B2(new_n459), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n706), .A2(new_n714), .ZN(G1328gat));
  NOR3_X1   g514(.A1(new_n704), .A2(G36gat), .A3(new_n462), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n713), .A2(new_n462), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n718), .A2(KEYINPUT106), .ZN(new_n719));
  OAI21_X1  g518(.A(G36gat), .B1(new_n718), .B2(KEYINPUT106), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(new_n719), .B2(new_n720), .ZN(G1329gat));
  NOR3_X1   g520(.A1(new_n704), .A2(G43gat), .A3(new_n687), .ZN(new_n722));
  INV_X1    g521(.A(new_n691), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n689), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n711), .B1(new_n500), .B2(new_n607), .ZN(new_n725));
  INV_X1    g524(.A(new_n709), .ZN(new_n726));
  AOI211_X1 g525(.A(new_n699), .B(new_n726), .C1(new_n467), .C2(new_n707), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n724), .B(new_n703), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n722), .B1(new_n728), .B2(G43gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(KEYINPUT107), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(KEYINPUT47), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n729), .A2(KEYINPUT107), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n731), .A2(new_n733), .ZN(G1330gat));
  OAI211_X1 g533(.A(KEYINPUT108), .B(G50gat), .C1(new_n713), .C2(new_n695), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n695), .A2(new_n739), .A3(G50gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n735), .A2(new_n736), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n736), .B1(new_n735), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(G1331gat));
  NOR4_X1   g543(.A1(new_n539), .A2(new_n637), .A3(new_n672), .A4(new_n607), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n708), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n459), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(new_n521), .ZN(G1332gat));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n462), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(G1333gat));
  NOR3_X1   g552(.A1(new_n746), .A2(G71gat), .A3(new_n687), .ZN(new_n754));
  INV_X1    g553(.A(new_n746), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n724), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n754), .B1(G71gat), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g557(.A1(new_n746), .A2(new_n695), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(new_n515), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n701), .A2(new_n672), .ZN(new_n761));
  INV_X1    g560(.A(new_n460), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT90), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT35), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n482), .A2(new_n495), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n695), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n724), .B1(new_n768), .B2(new_n497), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n607), .B(new_n761), .C1(new_n766), .C2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n708), .A2(KEYINPUT51), .A3(new_n607), .A4(new_n761), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n637), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n459), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n565), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n761), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n637), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n712), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n775), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n776), .B1(new_n780), .B2(new_n565), .ZN(G1336gat));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n772), .A2(new_n773), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n462), .A2(new_n637), .A3(G92gat), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n351), .B(new_n778), .C1(new_n725), .C2(new_n727), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G92gat), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n784), .B(KEYINPUT110), .Z(new_n790));
  NAND2_X1  g589(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n782), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n785), .A2(new_n787), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n786), .A2(G92gat), .B1(new_n783), .B2(new_n790), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n794), .B(KEYINPUT111), .C1(new_n789), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(G1337gat));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n724), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G99gat), .ZN(new_n799));
  INV_X1    g598(.A(new_n774), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n687), .A2(G99gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(G1338gat));
  NOR2_X1   g601(.A1(new_n695), .A2(G106gat), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n774), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n712), .A2(new_n271), .A3(new_n778), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n807), .A2(G106gat), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT53), .B1(new_n813), .B2(new_n804), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1339gat));
  NAND3_X1  g614(.A1(new_n608), .A2(new_n673), .A3(new_n637), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n622), .A2(new_n817), .A3(new_n624), .ZN(new_n818));
  INV_X1    g617(.A(new_n620), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n627), .B(new_n819), .C1(new_n626), .C2(KEYINPUT10), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(KEYINPUT54), .A3(new_n621), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n634), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n818), .A2(KEYINPUT55), .A3(new_n634), .A4(new_n821), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n824), .A2(new_n607), .A3(new_n636), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n639), .B1(new_n657), .B2(new_n640), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n659), .A2(new_n660), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n667), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n671), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n702), .A2(new_n671), .A3(new_n829), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT114), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n825), .A2(new_n636), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n672), .A3(new_n824), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(KEYINPUT114), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n831), .B1(new_n837), .B2(new_n699), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n816), .B1(new_n838), .B2(new_n701), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(new_n695), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n840), .A2(new_n775), .A3(new_n462), .A4(new_n411), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT115), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(G113gat), .A3(new_n672), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n839), .A2(new_n775), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(new_n461), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n462), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n357), .B1(new_n846), .B2(new_n673), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n843), .A2(new_n847), .ZN(G1340gat));
  NAND3_X1  g647(.A1(new_n842), .A2(G120gat), .A3(new_n702), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n358), .B1(new_n846), .B2(new_n637), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(G1341gat));
  INV_X1    g650(.A(new_n842), .ZN(new_n852));
  OAI21_X1  g651(.A(G127gat), .B1(new_n852), .B2(new_n539), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n846), .A2(G127gat), .A3(new_n539), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1342gat));
  OAI21_X1  g654(.A(G134gat), .B1(new_n852), .B2(new_n699), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n351), .A2(new_n699), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT116), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n845), .A2(new_n370), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT56), .Z(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n860), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n724), .A2(new_n695), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n351), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n673), .A2(G141gat), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT118), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n228), .A2(new_n229), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n692), .A2(new_n775), .A3(new_n462), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n695), .A2(KEYINPUT57), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n839), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n822), .A2(new_n873), .A3(new_n823), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n822), .B2(new_n823), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n825), .A2(new_n672), .A3(new_n636), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n637), .A2(new_n830), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n699), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n539), .B1(new_n880), .B2(new_n831), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n695), .B1(new_n881), .B2(new_n816), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n871), .B1(new_n872), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n868), .B1(new_n883), .B2(new_n673), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT58), .ZN(G1344gat));
  NAND2_X1  g685(.A1(new_n225), .A2(new_n226), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n864), .A2(new_n888), .A3(new_n702), .ZN(new_n889));
  XOR2_X1   g688(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n890));
  NOR2_X1   g689(.A1(new_n695), .A2(new_n872), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n839), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n822), .A2(new_n873), .A3(new_n823), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(new_n672), .A3(new_n636), .A4(new_n825), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n832), .B1(new_n895), .B2(new_n875), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n830), .B1(new_n826), .B2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n834), .A2(KEYINPUT120), .A3(new_n607), .A4(new_n824), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n896), .A2(new_n699), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n816), .B1(new_n900), .B2(new_n701), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n893), .B(KEYINPUT57), .C1(new_n901), .C2(new_n271), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n899), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n701), .B1(new_n879), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n816), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n271), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT121), .B1(new_n906), .B2(new_n872), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n892), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n869), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n702), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n890), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n871), .B(new_n702), .C1(new_n872), .C2(new_n882), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n888), .A2(KEYINPUT59), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n889), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT122), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n917), .B(new_n889), .C1(new_n911), .C2(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1345gat));
  INV_X1    g718(.A(G155gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n864), .A2(new_n920), .A3(new_n701), .ZN(new_n921));
  OAI21_X1  g720(.A(G155gat), .B1(new_n883), .B2(new_n539), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n883), .B2(new_n699), .ZN(new_n924));
  INV_X1    g723(.A(G162gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n858), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n924), .B1(new_n863), .B2(new_n926), .ZN(G1347gat));
  AND2_X1   g726(.A1(new_n839), .A2(new_n459), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(new_n351), .A3(new_n461), .ZN(new_n929));
  AOI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n672), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n840), .A2(new_n459), .A3(new_n351), .A4(new_n411), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n665), .A3(new_n673), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT123), .ZN(G1348gat));
  INV_X1    g733(.A(G176gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n929), .A2(new_n935), .A3(new_n702), .ZN(new_n936));
  OAI21_X1  g735(.A(G176gat), .B1(new_n931), .B2(new_n637), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1349gat));
  NAND3_X1  g737(.A1(new_n929), .A2(new_n291), .A3(new_n701), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n931), .A2(new_n539), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n311), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n931), .B2(new_n699), .ZN(new_n943));
  NOR2_X1   g742(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n290), .A3(new_n607), .ZN(new_n946));
  XNOR2_X1  g745(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n945), .B(new_n946), .C1(new_n943), .C2(new_n947), .ZN(G1351gat));
  AND3_X1   g747(.A1(new_n928), .A2(new_n351), .A3(new_n862), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n672), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n692), .A2(new_n459), .A3(new_n351), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n908), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n672), .A2(G197gat), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(G1352gat));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  AOI21_X1  g756(.A(G204gat), .B1(new_n957), .B2(KEYINPUT62), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n949), .A2(new_n702), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n959), .B(new_n960), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n908), .A2(new_n702), .A3(new_n952), .ZN(new_n962));
  INV_X1    g761(.A(G204gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(G1353gat));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n210), .A3(new_n701), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n951), .A2(new_n539), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n908), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(G1354gat));
  AOI21_X1  g769(.A(G218gat), .B1(new_n949), .B2(new_n607), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n953), .B(KEYINPUT127), .Z(new_n972));
  NOR2_X1   g771(.A1(new_n699), .A2(new_n211), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G1355gat));
endmodule


