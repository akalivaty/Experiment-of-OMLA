//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G116), .ZN(new_n214));
  INV_X1    g0014(.A(G270), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT65), .B(G244), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n212), .B(new_n216), .C1(G77), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n219), .A2(new_n221), .B1(G1), .B2(G20), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G20), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n230), .B1(new_n231), .B2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G13), .ZN(new_n233));
  NAND4_X1  g0033(.A1(new_n233), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n235), .B(G250), .C1(G257), .C2(G264), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT0), .Z(new_n237));
  NOR4_X1   g0037(.A1(new_n224), .A2(new_n225), .A3(new_n229), .A4(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G58), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  AND2_X1   g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G226), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n259), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G223), .A3(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G77), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G222), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n267), .B1(new_n268), .B2(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT67), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n263), .B1(new_n272), .B2(new_n273), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n265), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT69), .ZN(new_n282));
  INV_X1    g0082(.A(G58), .ZN(new_n283));
  OR3_X1    g0083(.A1(new_n283), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n227), .A2(G33), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n280), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(new_n228), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n288), .B2(new_n228), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n233), .A2(new_n227), .A3(G1), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n287), .A2(new_n293), .B1(new_n202), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n292), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n294), .B1(new_n296), .B2(new_n290), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n258), .A2(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(G50), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n278), .B(new_n300), .C1(G169), .C2(new_n276), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G20), .A2(G77), .ZN(new_n302));
  INV_X1    g0102(.A(new_n279), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT15), .B(G87), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n302), .B1(new_n281), .B2(new_n303), .C1(new_n286), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n293), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n297), .A2(G77), .A3(new_n298), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n294), .A2(new_n268), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n266), .A2(G238), .A3(G1698), .ZN(new_n311));
  INV_X1    g0111(.A(G107), .ZN(new_n312));
  INV_X1    g0112(.A(G232), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n311), .B1(new_n312), .B2(new_n266), .C1(new_n270), .C2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n263), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n261), .B1(new_n217), .B2(new_n264), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n310), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n317), .B1(new_n314), .B2(new_n315), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n277), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n310), .A2(KEYINPUT70), .B1(new_n319), .B2(G200), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n309), .B1(new_n322), .B2(G190), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n300), .B(KEYINPUT9), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n276), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n276), .A2(G190), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n301), .B(new_n329), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n279), .A2(G50), .B1(G20), .B2(new_n208), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n268), .B2(new_n286), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n293), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT11), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  INV_X1    g0145(.A(new_n294), .ZN(new_n346));
  OR3_X1    g0146(.A1(new_n346), .A2(KEYINPUT12), .A3(G68), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT12), .B1(new_n346), .B2(G68), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n208), .B1(new_n258), .B2(G20), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n347), .A2(new_n348), .B1(new_n297), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n344), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT14), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT13), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n266), .A2(G232), .A3(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT71), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT71), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n266), .A2(new_n356), .A3(G232), .A4(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G97), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n270), .B2(new_n262), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n315), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n261), .ZN(new_n363));
  INV_X1    g0163(.A(new_n264), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(G238), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n353), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n361), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n263), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n365), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT13), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n352), .B(G169), .C1(new_n366), .C2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n362), .A2(new_n353), .A3(new_n365), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT13), .B1(new_n368), .B2(new_n369), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(G179), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n373), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n352), .B1(new_n376), .B2(G169), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n351), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n351), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(G200), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n379), .B(new_n380), .C1(new_n381), .C2(new_n376), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n262), .A2(G1698), .ZN(new_n385));
  AND2_X1   g0185(.A1(KEYINPUT3), .A2(G33), .ZN(new_n386));
  NOR2_X1   g0186(.A1(KEYINPUT3), .A2(G33), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n385), .B1(G223), .B2(G1698), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n388), .A2(KEYINPUT73), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT73), .B1(new_n388), .B2(new_n389), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n315), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OR3_X1    g0192(.A1(new_n264), .A2(KEYINPUT74), .A3(new_n313), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT74), .B1(new_n264), .B2(new_n313), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n363), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n392), .A2(G179), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n320), .B1(new_n392), .B2(new_n395), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n384), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n392), .A2(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G169), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n392), .A2(G179), .A3(new_n395), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(KEYINPUT75), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n266), .B2(G20), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n386), .A2(new_n387), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n208), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n283), .A2(new_n208), .ZN(new_n408));
  OAI21_X1  g0208(.A(G20), .B1(new_n408), .B2(new_n201), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n303), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT16), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n407), .A2(KEYINPUT16), .A3(new_n411), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n293), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n285), .B1(new_n258), .B2(G20), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(new_n297), .B1(new_n294), .B2(new_n285), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n398), .A2(new_n402), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n398), .A2(new_n402), .A3(new_n418), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n399), .A2(G200), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n392), .A2(G190), .A3(new_n395), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n415), .A2(new_n423), .A3(new_n417), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n417), .ZN(new_n428));
  INV_X1    g0228(.A(new_n414), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n412), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n428), .B1(new_n293), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n431), .A2(KEYINPUT17), .A3(new_n424), .A4(new_n423), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n420), .A2(new_n422), .A3(new_n427), .A4(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n338), .A2(new_n383), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n296), .A2(new_n290), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n227), .B(G87), .C1(new_n386), .C2(new_n387), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT22), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(KEYINPUT85), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n266), .A2(new_n227), .A3(G87), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G116), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G20), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT23), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n227), .B2(G107), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n312), .A2(KEYINPUT23), .A3(G20), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n438), .A2(new_n441), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT24), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT24), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n438), .A2(new_n441), .A3(new_n447), .A4(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n435), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n233), .A2(G1), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n227), .A2(G107), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT86), .A3(KEYINPUT25), .ZN(new_n456));
  OR2_X1    g0256(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n453), .A2(new_n454), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n258), .A2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n435), .A2(new_n346), .A3(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n456), .B(new_n459), .C1(new_n461), .C2(new_n312), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n452), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(G257), .B(G1698), .C1(new_n386), .C2(new_n387), .ZN(new_n464));
  OAI211_X1 g0264(.A(G250), .B(new_n269), .C1(new_n386), .C2(new_n387), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G294), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n315), .ZN(new_n468));
  INV_X1    g0268(.A(G41), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n258), .B(G45), .C1(new_n469), .C2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G41), .ZN(new_n472));
  OAI211_X1 g0272(.A(G264), .B(new_n263), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(G41), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n258), .A4(G45), .ZN(new_n477));
  INV_X1    g0277(.A(new_n472), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n474), .A2(new_n477), .A3(new_n257), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n468), .A2(new_n473), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n331), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n468), .A2(new_n381), .A3(new_n473), .A4(new_n479), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(KEYINPUT87), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT87), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n484), .A3(new_n331), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n463), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n480), .A2(new_n320), .ZN(new_n487));
  OAI221_X1 g0287(.A(new_n487), .B1(G179), .B2(new_n480), .C1(new_n452), .C2(new_n462), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(G238), .B(new_n269), .C1(new_n386), .C2(new_n387), .ZN(new_n490));
  OAI211_X1 g0290(.A(G244), .B(G1698), .C1(new_n386), .C2(new_n387), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(new_n491), .A3(new_n442), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n315), .ZN(new_n493));
  INV_X1    g0293(.A(G45), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n211), .B1(new_n494), .B2(G1), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n258), .A2(new_n254), .A3(G45), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n263), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT79), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n493), .A2(KEYINPUT79), .A3(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(G190), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT79), .B1(new_n493), .B2(new_n498), .ZN(new_n506));
  AOI211_X1 g0306(.A(new_n500), .B(new_n497), .C1(new_n492), .C2(new_n315), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(KEYINPUT80), .A3(G190), .ZN(new_n509));
  OAI21_X1  g0309(.A(G200), .B1(new_n506), .B2(new_n507), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n297), .A2(G87), .A3(new_n460), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n266), .A2(new_n227), .A3(G68), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT19), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n227), .B1(new_n360), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(G87), .B2(new_n206), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n513), .B1(new_n286), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n293), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n304), .A2(new_n294), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n511), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n505), .A2(new_n509), .A3(new_n510), .A4(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n501), .A2(new_n277), .A3(new_n502), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n519), .B(new_n520), .C1(new_n304), .C2(new_n461), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n524), .C1(G169), .C2(new_n508), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(G244), .B(new_n269), .C1(new_n386), .C2(new_n387), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(KEYINPUT77), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(KEYINPUT77), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n266), .A2(G244), .A3(new_n530), .A4(new_n269), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n529), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n315), .ZN(new_n535));
  OAI211_X1 g0335(.A(G257), .B(new_n263), .C1(new_n470), .C2(new_n472), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n479), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n535), .A2(new_n277), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n320), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n312), .A2(KEYINPUT6), .A3(G97), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT6), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n545), .A2(new_n227), .B1(new_n268), .B2(new_n303), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n312), .B1(new_n404), .B2(new_n406), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(KEYINPUT76), .B2(new_n547), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n266), .A2(new_n403), .A3(G20), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT7), .B1(new_n405), .B2(new_n227), .ZN(new_n550));
  OAI21_X1  g0350(.A(G107), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT76), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n435), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n294), .A2(new_n516), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n461), .B2(new_n516), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n539), .B(new_n541), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n516), .A2(new_n312), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n544), .B1(new_n558), .B2(new_n205), .ZN(new_n559));
  INV_X1    g0359(.A(new_n542), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n551), .B2(new_n552), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n547), .A2(KEYINPUT76), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n293), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n556), .ZN(new_n566));
  AOI211_X1 g0366(.A(G190), .B(new_n537), .C1(new_n315), .C2(new_n534), .ZN(new_n567));
  AOI21_X1  g0367(.A(G200), .B1(new_n535), .B2(new_n538), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n565), .B(new_n566), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n557), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n526), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n489), .B1(new_n571), .B2(KEYINPUT81), .ZN(new_n572));
  OAI211_X1 g0372(.A(G264), .B(G1698), .C1(new_n386), .C2(new_n387), .ZN(new_n573));
  OAI211_X1 g0373(.A(G257), .B(new_n269), .C1(new_n386), .C2(new_n387), .ZN(new_n574));
  INV_X1    g0374(.A(G303), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(new_n266), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n315), .ZN(new_n577));
  OAI211_X1 g0377(.A(G270), .B(new_n263), .C1(new_n470), .C2(new_n472), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n479), .A2(KEYINPUT82), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT82), .B1(new_n479), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT83), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n288), .A2(new_n228), .B1(G20), .B2(new_n214), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n533), .B(new_n227), .C1(G33), .C2(new_n516), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(KEYINPUT83), .A3(new_n584), .A4(KEYINPUT20), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n586), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n214), .B1(new_n297), .B2(new_n460), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n294), .A2(G116), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n581), .A2(new_n593), .A3(KEYINPUT21), .A4(G169), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n479), .A2(new_n578), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n479), .A2(KEYINPUT82), .A3(new_n578), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n315), .B2(new_n576), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G179), .A3(new_n593), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n581), .A2(new_n593), .A3(G169), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n593), .ZN(new_n606));
  OAI211_X1 g0406(.A(G190), .B(new_n577), .C1(new_n579), .C2(new_n580), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n599), .C2(new_n331), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n601), .A2(new_n602), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(new_n605), .A3(new_n600), .A4(new_n594), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT84), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n522), .A2(new_n557), .A3(new_n569), .A4(new_n525), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT81), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n609), .A2(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n434), .A2(new_n572), .A3(new_n614), .ZN(G372));
  INV_X1    g0415(.A(new_n337), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n335), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n432), .A2(new_n427), .ZN(new_n618));
  INV_X1    g0418(.A(new_n324), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n382), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n618), .B1(new_n620), .B2(new_n378), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n400), .A2(new_n401), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n418), .A2(new_n421), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n421), .B1(new_n418), .B2(new_n622), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n617), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n301), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n434), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n499), .A2(new_n320), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n523), .A2(new_n524), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n499), .A2(G200), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n503), .A2(new_n521), .A3(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n486), .A2(new_n557), .A3(new_n569), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n601), .A2(new_n488), .A3(new_n605), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n547), .A2(KEYINPUT76), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n553), .A2(new_n638), .A3(new_n562), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n556), .B1(new_n639), .B2(new_n293), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n537), .B1(new_n534), .B2(new_n315), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n539), .B1(G169), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n522), .A2(KEYINPUT26), .A3(new_n643), .A4(new_n525), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n631), .A2(new_n634), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n557), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n637), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n628), .B1(new_n629), .B2(new_n650), .ZN(G369));
  NAND2_X1  g0451(.A1(new_n453), .A2(new_n227), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n611), .A2(new_n609), .B1(new_n593), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n601), .A2(new_n605), .ZN(new_n659));
  INV_X1    g0459(.A(new_n657), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n659), .A2(new_n606), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G330), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n489), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n463), .B2(new_n660), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n488), .B2(new_n660), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n657), .B(KEYINPUT88), .Z(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n488), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n659), .A2(new_n657), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n671), .B1(new_n672), .B2(new_n665), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0475(.A(new_n235), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n677), .A2(new_n258), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n226), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n677), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT28), .Z(new_n683));
  NAND3_X1  g0483(.A1(new_n572), .A2(new_n614), .A3(new_n669), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT31), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n540), .A2(new_n480), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT90), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n493), .A2(new_n687), .A3(new_n498), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n499), .A2(KEYINPUT90), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n581), .A2(new_n277), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n686), .B1(new_n690), .B2(KEYINPUT91), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n689), .A2(new_n688), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT91), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(new_n277), .A4(new_n581), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n691), .A2(KEYINPUT93), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT93), .B1(new_n691), .B2(new_n694), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT92), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n468), .A2(new_n473), .A3(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n641), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g0500(.A(G179), .B(new_n577), .C1(new_n579), .C2(new_n580), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n697), .A2(KEYINPUT92), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n700), .A2(new_n702), .A3(new_n508), .A4(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n501), .A2(new_n641), .A3(new_n699), .A4(new_n502), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n706), .B2(new_n701), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n695), .A2(new_n696), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n685), .B1(new_n709), .B2(new_n660), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n691), .A2(new_n694), .ZN(new_n711));
  OAI211_X1 g0511(.A(KEYINPUT31), .B(new_n670), .C1(new_n711), .C2(new_n708), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n684), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT26), .B1(new_n646), .B2(new_n557), .ZN(new_n715));
  AND4_X1   g0515(.A1(new_n488), .A2(new_n605), .A3(new_n600), .A4(new_n594), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n557), .A2(new_n569), .A3(new_n486), .A4(new_n634), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n715), .B(new_n631), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n526), .A2(KEYINPUT26), .A3(new_n557), .ZN(new_n719));
  OAI211_X1 g0519(.A(KEYINPUT29), .B(new_n660), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT94), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n670), .B1(new_n637), .B2(new_n648), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(KEYINPUT29), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n714), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n683), .B1(new_n726), .B2(G1), .ZN(G364));
  INV_X1    g0527(.A(new_n664), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n233), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n258), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n677), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n662), .A2(new_n663), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n728), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n662), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n235), .A2(G355), .A3(new_n266), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n252), .A2(new_n494), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n676), .A2(new_n266), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G45), .B2(new_n226), .ZN(new_n743));
  OAI221_X1 g0543(.A(new_n740), .B1(G116), .B2(new_n235), .C1(new_n741), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n228), .B1(G20), .B2(new_n320), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n738), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT95), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n733), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n745), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n227), .A2(G179), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G190), .A2(G200), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT96), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT96), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n410), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT32), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n227), .A2(new_n277), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n752), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n268), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n751), .A2(G190), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n210), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n759), .A2(new_n381), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n761), .B(new_n763), .C1(G68), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n751), .A2(new_n381), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n312), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n759), .A2(G190), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n331), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n405), .B(new_n768), .C1(G50), .C2(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n381), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n227), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n516), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n769), .A2(G200), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G58), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n758), .A2(new_n766), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT97), .Z(new_n778));
  NAND2_X1  g0578(.A1(new_n770), .A2(G326), .ZN(new_n779));
  INV_X1    g0579(.A(G294), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n780), .B2(new_n773), .ZN(new_n781));
  INV_X1    g0581(.A(new_n760), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n781), .A2(KEYINPUT98), .B1(G311), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(KEYINPUT98), .B2(new_n781), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT99), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  INV_X1    g0586(.A(new_n762), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n765), .A2(new_n786), .B1(new_n787), .B2(G303), .ZN(new_n788));
  INV_X1    g0588(.A(new_n767), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n266), .B1(new_n789), .B2(G283), .ZN(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  INV_X1    g0591(.A(new_n775), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n788), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n756), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(G329), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n778), .B1(new_n785), .B2(new_n795), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n739), .B(new_n749), .C1(new_n750), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n735), .A2(new_n797), .ZN(G396));
  NAND3_X1  g0598(.A1(new_n321), .A2(new_n323), .A3(new_n660), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n325), .A2(new_n327), .B1(new_n309), .B2(new_n657), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n669), .B(new_n799), .C1(new_n619), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n644), .A2(new_n647), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n631), .B1(new_n716), .B2(new_n717), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n309), .A2(new_n657), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n328), .A2(new_n806), .B1(new_n323), .B2(new_n321), .ZN(new_n807));
  INV_X1    g0607(.A(new_n799), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n805), .B1(new_n722), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n732), .B1(new_n714), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n714), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n745), .A2(new_n736), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n733), .B1(new_n268), .B2(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n789), .A2(G87), .B1(new_n782), .B2(G116), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(new_n764), .C1(new_n756), .C2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n405), .B1(new_n762), .B2(new_n312), .ZN(new_n819));
  INV_X1    g0619(.A(new_n770), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n792), .A2(new_n780), .B1(new_n820), .B2(new_n575), .ZN(new_n821));
  NOR4_X1   g0621(.A1(new_n818), .A2(new_n774), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n789), .A2(G68), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n202), .B2(new_n762), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT100), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n765), .A2(G150), .B1(new_n782), .B2(G159), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n775), .A2(G143), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n820), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT34), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n266), .B1(new_n283), .B2(new_n773), .C1(new_n756), .C2(new_n832), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n825), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n829), .A2(new_n830), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n822), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n814), .B1(new_n750), .B2(new_n836), .C1(new_n809), .C2(new_n737), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n812), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  INV_X1    g0639(.A(KEYINPUT104), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n378), .A2(new_n382), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n351), .A2(new_n657), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT104), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n375), .A2(new_n842), .A3(new_n377), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n843), .A2(new_n846), .A3(new_n809), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n696), .A2(new_n708), .ZN(new_n848));
  OAI211_X1 g0648(.A(KEYINPUT31), .B(new_n657), .C1(new_n848), .C2(new_n695), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n684), .A2(new_n710), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  INV_X1    g0653(.A(new_n655), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n418), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n618), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n623), .A2(new_n624), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n419), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n855), .A2(new_n425), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n418), .A2(new_n622), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n855), .A3(new_n425), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n860), .A2(new_n861), .B1(new_n863), .B2(KEYINPUT37), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n853), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n855), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n433), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n419), .A2(new_n859), .A3(new_n425), .A4(new_n855), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n852), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n851), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n867), .A2(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n853), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n871), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n850), .A3(new_n847), .ZN(new_n877));
  XOR2_X1   g0677(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n434), .A2(new_n850), .ZN(new_n881));
  OAI21_X1  g0681(.A(G330), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n801), .B1(new_n637), .B2(new_n648), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT103), .B1(new_n884), .B2(new_n808), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT103), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n805), .A2(new_n886), .A3(new_n799), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n843), .A2(new_n846), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n876), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n870), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n866), .B1(new_n625), .B2(new_n618), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n893), .B2(new_n870), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n891), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n875), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n378), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n660), .ZN(new_n899));
  OAI221_X1 g0699(.A(new_n890), .B1(new_n857), .B2(new_n854), .C1(new_n897), .C2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n629), .B1(new_n723), .B2(new_n724), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(new_n627), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n900), .B(new_n902), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n883), .A2(new_n903), .B1(new_n258), .B2(new_n729), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n903), .B2(new_n883), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n561), .A2(KEYINPUT35), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n228), .A2(new_n227), .A3(new_n214), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n561), .B2(KEYINPUT35), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT101), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n909), .B2(new_n908), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT36), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n408), .A2(new_n226), .A3(new_n268), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT102), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n913), .A2(new_n914), .B1(new_n202), .B2(G68), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n258), .B(G13), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  OR3_X1    g0717(.A1(new_n905), .A2(new_n912), .A3(new_n917), .ZN(G367));
  NOR3_X1   g0718(.A1(new_n245), .A2(new_n676), .A3(new_n266), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n746), .B1(new_n235), .B2(new_n304), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n732), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n266), .B1(new_n762), .B2(new_n283), .C1(new_n268), .C2(new_n767), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n794), .B2(G137), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n764), .A2(new_n410), .B1(new_n760), .B2(new_n202), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT107), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n775), .A2(G150), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n773), .A2(new_n208), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(G143), .B2(new_n770), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n923), .A2(new_n925), .A3(new_n926), .A4(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT108), .Z(new_n930));
  NOR2_X1   g0730(.A1(new_n762), .A2(new_n214), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n820), .A2(new_n817), .B1(KEYINPUT46), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(KEYINPUT46), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n794), .A2(G317), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n764), .A2(new_n780), .B1(new_n760), .B2(new_n816), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n266), .B(new_n935), .C1(G97), .C2(new_n789), .ZN(new_n936));
  INV_X1    g0736(.A(new_n773), .ZN(new_n937));
  AOI22_X1  g0737(.A1(G107), .A2(new_n937), .B1(new_n775), .B2(G303), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n933), .A2(new_n934), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n930), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT47), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n921), .B1(new_n941), .B2(new_n745), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n521), .A2(new_n660), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n632), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT106), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n646), .A2(new_n943), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n945), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n738), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n942), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n557), .B(new_n569), .C1(new_n640), .C2(new_n669), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n643), .A2(new_n670), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n673), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT45), .Z(new_n958));
  NOR2_X1   g0758(.A1(new_n673), .A2(new_n956), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n668), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n672), .A2(new_n665), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n667), .B2(new_n672), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n664), .B(new_n965), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n726), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n677), .B(KEYINPUT41), .Z(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n731), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n954), .A2(new_n488), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n670), .B1(new_n971), .B2(new_n557), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n672), .A2(new_n665), .A3(new_n956), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n972), .B1(new_n973), .B2(KEYINPUT42), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(KEYINPUT42), .B2(new_n973), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT43), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n976), .B2(new_n950), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n950), .A2(new_n976), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n956), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n668), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n953), .B1(new_n970), .B2(new_n982), .ZN(G387));
  INV_X1    g0783(.A(new_n966), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n667), .A2(new_n952), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n742), .B1(new_n242), .B2(new_n494), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n679), .A2(new_n235), .A3(new_n266), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n281), .A2(KEYINPUT50), .A3(G50), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT50), .B1(new_n281), .B2(G50), .ZN(new_n990));
  AOI21_X1  g0790(.A(G45), .B1(G68), .B2(G77), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n989), .A2(new_n678), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n988), .A2(new_n992), .B1(new_n312), .B2(new_n676), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n732), .B1(new_n993), .B2(new_n747), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n765), .A2(G311), .B1(new_n782), .B2(G303), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n775), .A2(G317), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(new_n791), .C2(new_n820), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT48), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n816), .B2(new_n773), .C1(new_n780), .C2(new_n762), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n997), .A2(new_n998), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT49), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n794), .A2(G326), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n266), .B1(new_n789), .B2(G116), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1002), .A2(KEYINPUT49), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n773), .A2(new_n304), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G159), .B2(new_n770), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n202), .B2(new_n792), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n794), .A2(G150), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n268), .A2(new_n762), .B1(new_n760), .B2(new_n208), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n405), .B(new_n1012), .C1(G97), .C2(new_n789), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n765), .A2(new_n284), .A3(new_n282), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1006), .A2(new_n1007), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n994), .B1(new_n1016), .B2(new_n745), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n984), .A2(new_n731), .B1(new_n985), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n984), .A2(new_n726), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n677), .B1(new_n966), .B2(new_n725), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(G393));
  AND2_X1   g0821(.A1(new_n249), .A2(new_n742), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n746), .B1(new_n516), .B2(new_n235), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n732), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n266), .B1(new_n767), .B2(new_n210), .C1(new_n773), .C2(new_n268), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n762), .A2(new_n208), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n764), .A2(new_n202), .B1(new_n760), .B2(new_n281), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(G143), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n756), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G150), .A2(new_n770), .B1(new_n775), .B2(G159), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n1032));
  XNOR2_X1  g0832(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n266), .B(new_n768), .C1(G116), .C2(new_n937), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n764), .A2(new_n575), .B1(new_n760), .B2(new_n780), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G283), .B2(new_n787), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(new_n791), .C2(new_n756), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G311), .A2(new_n775), .B1(new_n770), .B2(G317), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1030), .A2(new_n1033), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1024), .B1(new_n1040), .B2(new_n745), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n956), .B2(new_n952), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n963), .B2(new_n730), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n677), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n961), .B(new_n668), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n966), .A2(new_n725), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n963), .B1(new_n725), .B2(new_n966), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1043), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(G390));
  AOI21_X1  g0850(.A(KEYINPUT39), .B1(new_n865), .B2(new_n871), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT38), .B1(new_n867), .B2(new_n870), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n892), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1051), .B1(new_n1053), .B2(KEYINPUT39), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(new_n737), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n823), .B1(new_n312), .B2(new_n764), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G97), .B2(new_n782), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n266), .B(new_n763), .C1(G283), .C2(new_n770), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n780), .C2(new_n756), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n792), .A2(new_n214), .B1(new_n268), .B2(new_n773), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT115), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n794), .A2(G125), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n266), .B1(new_n767), .B2(new_n202), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT114), .Z(new_n1064));
  INV_X1    g0864(.A(G150), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n762), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT53), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1062), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G128), .A2(new_n770), .B1(new_n775), .B2(G132), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT54), .B(G143), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n765), .A2(G137), .B1(new_n782), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1069), .B(new_n1072), .C1(new_n410), .C2(new_n773), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1059), .A2(new_n1061), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n745), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n285), .A2(new_n813), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n732), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1055), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n847), .A2(G330), .A3(new_n850), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n884), .A2(KEYINPUT103), .A3(new_n808), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n886), .B1(new_n805), .B2(new_n799), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n889), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1083), .A2(new_n899), .B1(new_n895), .B2(new_n896), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n807), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n660), .B(new_n1085), .C1(new_n718), .C2(new_n719), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1086), .A2(new_n799), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n843), .A2(new_n846), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n899), .B1(new_n892), .B2(new_n894), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1080), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n899), .B1(new_n892), .B2(new_n894), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n889), .A2(new_n713), .A3(G330), .A4(new_n809), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n888), .A2(new_n889), .B1(new_n898), .B2(new_n660), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1094), .C1(new_n1054), .C2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(KEYINPUT113), .B1(new_n1097), .B2(new_n730), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT113), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1092), .A2(new_n1096), .A3(new_n1099), .A4(new_n731), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1078), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT112), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n850), .A2(G330), .A3(new_n809), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1088), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n1087), .A3(new_n1094), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n850), .A2(G330), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n713), .A2(G330), .A3(new_n809), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1106), .A2(new_n847), .B1(new_n1107), .B2(new_n1088), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n888), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n434), .A2(new_n850), .A3(G330), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n901), .A2(new_n1111), .A3(new_n627), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1110), .A2(new_n1092), .A3(new_n1096), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n677), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT110), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT110), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1116), .A3(new_n677), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT111), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1097), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1092), .A2(new_n1096), .A3(KEYINPUT111), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1105), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1107), .A2(new_n1088), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1109), .B1(new_n1123), .B2(new_n1079), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1112), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1120), .A2(new_n1121), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1102), .B1(new_n1118), .B2(new_n1126), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1113), .A2(new_n1116), .A3(new_n677), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1116), .B1(new_n1113), .B2(new_n677), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1102), .B(new_n1126), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1101), .B1(new_n1127), .B2(new_n1131), .ZN(G378));
  XOR2_X1   g0932(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n300), .A2(new_n854), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT55), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n617), .A2(new_n301), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n617), .B2(new_n301), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1134), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n617), .A2(new_n301), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1136), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n617), .A2(new_n301), .A3(new_n1136), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1133), .A3(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(new_n737), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n266), .A2(G41), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1147), .B1(new_n767), .B2(new_n283), .C1(new_n268), .C2(new_n762), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n794), .B2(G283), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n764), .A2(new_n516), .B1(new_n760), .B2(new_n304), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT116), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n775), .A2(G107), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n927), .B1(G116), .B2(new_n770), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT58), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1149), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n775), .A2(G128), .B1(new_n787), .B2(new_n1071), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT117), .Z(new_n1160));
  NOR2_X1   g0960(.A1(new_n773), .A2(new_n1065), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n764), .A2(new_n832), .B1(new_n760), .B2(new_n828), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1161), .B(new_n1162), .C1(G125), .C2(new_n770), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n794), .A2(G124), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G33), .B(G41), .C1(new_n789), .C2(G159), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1158), .B1(new_n1157), .B2(new_n1156), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n745), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n813), .A2(new_n202), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n732), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1146), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT119), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n851), .A2(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1145), .B1(new_n1176), .B2(G330), .ZN(new_n1177));
  AND4_X1   g0977(.A1(G330), .A2(new_n873), .A3(new_n879), .A4(new_n1145), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1175), .B(new_n900), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1145), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n880), .B2(new_n663), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1176), .A2(G330), .A3(new_n1145), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n900), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(new_n1182), .C1(KEYINPUT119), .C2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1174), .B1(new_n1185), .B2(new_n731), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1183), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1181), .A2(new_n900), .A3(new_n1182), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(KEYINPUT57), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1113), .A2(new_n1112), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n677), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1186), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT120), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1194), .B(new_n1195), .ZN(G375));
  NAND2_X1  g0996(.A1(new_n1110), .A2(new_n731), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n733), .B1(new_n208), .B2(new_n813), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G97), .A2(new_n787), .B1(new_n782), .B2(G107), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n214), .B2(new_n764), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n405), .B1(new_n268), .B2(new_n767), .C1(new_n820), .C2(new_n780), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(G303), .C2(new_n794), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1008), .B1(G283), .B2(new_n775), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT121), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n266), .B1(new_n767), .B2(new_n283), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n792), .A2(new_n828), .B1(new_n820), .B2(new_n832), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(G50), .C2(new_n937), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G159), .A2(new_n787), .B1(new_n782), .B2(G150), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n764), .B2(new_n1070), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G128), .B2(new_n794), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1202), .A2(new_n1204), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1198), .B1(new_n750), .B2(new_n1211), .C1(new_n889), .C2(new_n737), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1197), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1124), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1111), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n724), .A2(new_n723), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n434), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1218), .A3(new_n628), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1215), .A2(new_n1219), .A3(new_n1105), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1125), .A2(new_n1220), .A3(new_n969), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1214), .A2(new_n1221), .ZN(G381));
  XNOR2_X1  g1022(.A(new_n1194), .B(KEYINPUT120), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1101), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1049), .A2(new_n838), .ZN(new_n1226));
  OR2_X1    g1026(.A1(G393), .A2(G396), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(G387), .A2(new_n1226), .A3(G381), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT122), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1225), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1223), .B(new_n1230), .C1(new_n1229), .C2(new_n1228), .ZN(G407));
  INV_X1    g1031(.A(new_n1225), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n656), .A2(G213), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1223), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(G213), .A3(new_n1235), .ZN(G409));
  OAI211_X1 g1036(.A(G390), .B(new_n953), .C1(new_n970), .C2(new_n982), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(new_n1049), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(G393), .A2(G396), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1227), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT125), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1243), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1237), .B(new_n1238), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1185), .A2(new_n969), .A3(new_n1190), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1174), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1187), .A2(new_n1188), .A3(new_n731), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n1101), .A3(new_n1224), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1101), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1224), .A2(KEYINPUT112), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n1130), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1254), .B1(new_n1257), .B2(new_n1194), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1233), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1125), .A2(KEYINPUT60), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1220), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1215), .A2(KEYINPUT60), .A3(new_n1219), .A4(new_n1105), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1262), .A2(new_n677), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1214), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n838), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(G384), .A3(new_n1214), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1234), .A2(G2897), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT123), .Z(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1269), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G384), .B1(new_n1264), .B2(new_n1214), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n838), .B(new_n1213), .C1(new_n1261), .C2(new_n1263), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1271), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1270), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT61), .B1(new_n1259), .B2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1258), .A2(new_n1233), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1279), .A2(KEYINPUT62), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1249), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT63), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1279), .A2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1233), .A4(new_n1278), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT61), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1259), .B2(new_n1276), .ZN(new_n1291));
  AOI211_X1 g1091(.A(KEYINPUT124), .B(new_n1275), .C1(new_n1258), .C2(new_n1233), .ZN(new_n1292));
  NOR4_X1   g1092(.A1(new_n1288), .A2(new_n1289), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1185), .A2(new_n731), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1251), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1192), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1193), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G378), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1234), .B1(new_n1299), .B2(new_n1254), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT63), .B1(new_n1300), .B2(new_n1278), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT126), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1283), .B1(new_n1293), .B2(new_n1305), .ZN(G405));
  NOR2_X1   g1106(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1299), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1278), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G375), .A2(new_n1232), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1278), .B1(new_n1311), .B2(new_n1299), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT127), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1309), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1311), .A2(new_n1299), .A3(new_n1278), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1313), .A2(new_n1249), .A3(new_n1317), .ZN(new_n1318));
  OAI211_X1 g1118(.A(KEYINPUT127), .B(new_n1248), .C1(new_n1310), .C2(new_n1312), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(G402));
endmodule


