//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT66), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT67), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(KEYINPUT68), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n460), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n462), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(G137), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n470), .A2(new_n472), .A3(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n473), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(G136), .B2(new_n483), .ZN(G162));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  AND2_X1   g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n458), .B2(new_n459), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT69), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(new_n488), .C1(new_n458), .C2(new_n459), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n460), .A2(new_n466), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n474), .C1(new_n458), .C2(new_n459), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n507), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n509), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(new_n505), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n516), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n508), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n506), .B2(new_n507), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n505), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT72), .B(G52), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n529), .A2(G90), .B1(new_n508), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n533), .A2(new_n534), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n505), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n529), .A2(G81), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n508), .A2(G43), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(KEYINPUT73), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(KEYINPUT73), .B1(new_n543), .B2(new_n544), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  XNOR2_X1  g129(.A(new_n528), .B(KEYINPUT74), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g132(.A1(G78), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n508), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n508), .A2(new_n563), .A3(G53), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n562), .A2(new_n564), .B1(G91), .B2(new_n529), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n559), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  NAND2_X1  g143(.A1(new_n529), .A2(G87), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n508), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n508), .A2(G48), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n512), .B2(new_n513), .ZN(new_n575));
  INV_X1    g150(.A(G73), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n502), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n511), .A2(G86), .A3(new_n514), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(new_n529), .A2(G85), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n508), .A2(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n581), .B(new_n582), .C1(new_n505), .C2(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT75), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT75), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G290));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n555), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g164(.A1(G79), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n515), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n594), .A2(new_n595), .B1(G54), .B2(new_n508), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(G171), .ZN(G284));
  OAI21_X1  g175(.A(new_n599), .B1(new_n598), .B2(G171), .ZN(G321));
  NOR2_X1   g176(.A1(G286), .A2(new_n598), .ZN(new_n602));
  XNOR2_X1  g177(.A(G299), .B(KEYINPUT76), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n598), .ZN(G297));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n598), .ZN(G280));
  INV_X1    g180(.A(new_n597), .ZN(new_n606));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g187(.A1(new_n460), .A2(new_n466), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n613), .A2(new_n471), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT12), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT77), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n483), .A2(G135), .ZN(new_n623));
  INV_X1    g198(.A(new_n479), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G123), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n474), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n623), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2096), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n620), .B2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT79), .Z(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT80), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n646), .A2(G14), .A3(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT82), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  OAI21_X1  g233(.A(KEYINPUT17), .B1(new_n650), .B2(new_n651), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(new_n653), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n653), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n652), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT83), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT20), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n667), .A2(new_n669), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n676), .A2(new_n672), .A3(new_n670), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n674), .B(new_n677), .C1(new_n672), .C2(new_n676), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT84), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n683), .A2(new_n686), .A3(new_n684), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(G229));
  XOR2_X1   g265(.A(KEYINPUT31), .B(G11), .Z(new_n691));
  INV_X1    g266(.A(G28), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(KEYINPUT30), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT95), .ZN(new_n694));
  AOI21_X1  g269(.A(G29), .B1(new_n692), .B2(KEYINPUT30), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n691), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NOR2_X1   g273(.A1(G168), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n698), .B2(G21), .ZN(new_n700));
  INV_X1    g275(.A(G1966), .ZN(new_n701));
  OAI221_X1 g276(.A(new_n696), .B1(new_n697), .B2(new_n628), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G1961), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n698), .A2(G5), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G171), .B2(new_n698), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n704), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NOR2_X1   g287(.A1(G29), .A2(G35), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G162), .B2(G29), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2090), .ZN(new_n717));
  NOR2_X1   g292(.A1(G27), .A2(G29), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G164), .B2(G29), .ZN(new_n719));
  INV_X1    g294(.A(G2078), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n722));
  INV_X1    g297(.A(G34), .ZN(new_n723));
  AOI21_X1  g298(.A(G29), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G160), .B2(new_n697), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n721), .B1(G2084), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n717), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G4), .A2(G16), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n606), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G1348), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n711), .A2(new_n712), .A3(new_n728), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n697), .A2(G32), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n624), .A2(G129), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT26), .Z(new_n738));
  NAND3_X1  g313(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n697), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT27), .ZN(new_n743));
  INV_X1    g318(.A(G1996), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n613), .A2(G127), .ZN(new_n746));
  INV_X1    g321(.A(G115), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n462), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n474), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n483), .A2(G139), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(G29), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G33), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(G29), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G2072), .Z(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G19), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n549), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT90), .B(G1341), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n698), .A2(G20), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT23), .Z(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G299), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1956), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n708), .A2(new_n705), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n697), .A2(G26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G128), .ZN(new_n777));
  OR3_X1    g352(.A1(new_n479), .A2(KEYINPUT91), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT91), .B1(new_n479), .B2(new_n777), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n781));
  INV_X1    g356(.A(G116), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(G2105), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n483), .B2(G140), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n776), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2067), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n726), .A2(G2084), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n772), .A2(new_n773), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n733), .A2(new_n745), .A3(new_n768), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G24), .B(G290), .S(G16), .Z(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT87), .Z(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(G1986), .ZN(new_n794));
  NOR2_X1   g369(.A1(G25), .A2(G29), .ZN(new_n795));
  OR2_X1    g370(.A1(G95), .A2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT85), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n483), .A2(G131), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n624), .A2(G119), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n795), .B1(new_n802), .B2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT86), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n793), .A2(G1986), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n698), .A2(G22), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G166), .B2(new_n698), .ZN(new_n809));
  INV_X1    g384(.A(G1971), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n698), .A2(G23), .ZN(new_n812));
  INV_X1    g387(.A(G288), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n698), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT33), .B(G1976), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G6), .B(G305), .S(G16), .Z(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n811), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT34), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n794), .A2(new_n806), .A3(new_n807), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(KEYINPUT34), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT88), .Z(new_n824));
  NOR2_X1   g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g402(.A(KEYINPUT89), .B(KEYINPUT36), .C1(new_n822), .C2(new_n824), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n791), .B1(new_n827), .B2(new_n828), .ZN(G311));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(new_n790), .ZN(G150));
  NOR2_X1   g406(.A1(new_n597), .A2(new_n607), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n505), .A2(new_n835), .B1(new_n515), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n508), .A2(G55), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n548), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n839), .B(new_n542), .C1(new_n546), .C2(new_n547), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n834), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT100), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT99), .B(G860), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n844), .B2(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n840), .A2(new_n848), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  XNOR2_X1  g428(.A(G160), .B(new_n628), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n618), .A2(KEYINPUT102), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n618), .A2(KEYINPUT102), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  INV_X1    g434(.A(G118), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n860), .B2(G2105), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n624), .B2(G130), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n483), .A2(G142), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n856), .A2(new_n868), .A3(new_n857), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n867), .A2(new_n869), .A3(new_n801), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n801), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n740), .B(G164), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n875));
  INV_X1    g450(.A(new_n785), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n752), .A2(new_n758), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n752), .B2(new_n758), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  INV_X1    g456(.A(new_n875), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n874), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n873), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n872), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n872), .B1(new_n886), .B2(new_n884), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n855), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n884), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n871), .B2(new_n870), .ZN(new_n893));
  INV_X1    g468(.A(new_n855), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n893), .A2(new_n888), .A3(new_n894), .A4(new_n887), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g473(.A1(G303), .A2(G305), .ZN(new_n899));
  NAND2_X1  g474(.A1(G303), .A2(G305), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(G288), .B1(new_n585), .B2(new_n586), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n585), .A2(G288), .A3(new_n586), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n899), .A2(KEYINPUT106), .A3(new_n900), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n903), .A2(new_n905), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n906), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n902), .B(new_n901), .C1(new_n909), .C2(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT42), .Z(new_n912));
  NAND2_X1  g487(.A1(new_n597), .A2(G299), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n559), .A2(new_n591), .A3(new_n565), .A4(new_n596), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n915), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n843), .B(new_n609), .ZN(new_n921));
  MUX2_X1   g496(.A(new_n919), .B(new_n920), .S(new_n921), .Z(new_n922));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n912), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n912), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(G868), .B2(new_n839), .ZN(G295));
  OAI21_X1  g504(.A(new_n928), .B1(G868), .B2(new_n839), .ZN(G331));
  AND3_X1   g505(.A1(new_n841), .A2(new_n842), .A3(G286), .ZN(new_n931));
  AOI21_X1  g506(.A(G286), .B1(new_n841), .B2(new_n842), .ZN(new_n932));
  OAI21_X1  g507(.A(G301), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n843), .A2(G168), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n841), .A2(new_n842), .A3(G286), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(G171), .A3(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n933), .A2(new_n936), .A3(new_n919), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n915), .B1(new_n933), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n911), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n931), .A2(new_n932), .A3(G301), .ZN(new_n940));
  AOI21_X1  g515(.A(G171), .B1(new_n934), .B2(new_n935), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n920), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n911), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n933), .A2(new_n936), .A3(new_n919), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n939), .A2(new_n945), .A3(new_n946), .A4(new_n896), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT110), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n896), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n916), .A2(KEYINPUT109), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n916), .A2(KEYINPUT109), .A3(new_n918), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n936), .A3(new_n933), .A4(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n943), .B1(new_n952), .B2(new_n942), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n947), .A2(KEYINPUT110), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n939), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n949), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT108), .ZN(new_n960));
  OR3_X1    g535(.A1(new_n949), .A2(new_n953), .A3(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n963), .B(KEYINPUT43), .C1(new_n949), .C2(new_n958), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n961), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n957), .A2(new_n965), .ZN(G397));
  INV_X1    g541(.A(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n785), .A2(G2067), .ZN(new_n968));
  INV_X1    g543(.A(G2067), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n780), .A2(new_n969), .A3(new_n784), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n968), .A2(KEYINPUT113), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT113), .B1(new_n968), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n741), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n493), .B2(new_n499), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n974), .A2(KEYINPUT111), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n974), .B2(KEYINPUT111), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n475), .A2(G40), .A3(new_n472), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n469), .B2(G2105), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n973), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n744), .B1(new_n971), .B2(new_n972), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n744), .A3(new_n980), .ZN(new_n985));
  OR3_X1    g560(.A1(new_n985), .A2(KEYINPUT112), .A3(new_n740), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT112), .B1(new_n985), .B2(new_n740), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n983), .A2(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n801), .B(new_n805), .Z(new_n989));
  NAND2_X1  g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(G290), .B(G1986), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n982), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n974), .A2(new_n980), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT115), .B1(new_n995), .B2(G8), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n997));
  INV_X1    g572(.A(G8), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n997), .B(new_n998), .C1(new_n974), .C2(new_n980), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n528), .A2(new_n574), .B1(new_n576), .B2(new_n502), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n1001), .A2(G651), .B1(new_n508), .B2(G48), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n579), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G305), .A2(G1981), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1002), .B2(new_n579), .ZN(new_n1007));
  AND4_X1   g582(.A1(new_n1003), .A2(new_n573), .A3(new_n578), .A4(new_n579), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT49), .ZN(new_n1009));
  OAI22_X1  g584(.A1(new_n996), .A2(new_n999), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n813), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n995), .A2(KEYINPUT115), .A3(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n995), .A2(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n997), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1012), .A2(new_n1004), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1013), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n813), .A2(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT116), .B(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1020), .B(new_n1023), .C1(new_n996), .C2(new_n999), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1010), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1017), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1020), .B1(new_n996), .B2(new_n999), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT52), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(KEYINPUT117), .A3(new_n1024), .A4(new_n1010), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n976), .A2(G1384), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n500), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1032), .B(new_n980), .C1(KEYINPUT45), .C2(new_n974), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n810), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n496), .A2(new_n498), .ZN(new_n1036));
  INV_X1    g611(.A(new_n487), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n491), .B1(new_n473), .B2(new_n488), .ZN(new_n1038));
  INV_X1    g613(.A(new_n492), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT50), .ZN(new_n1042));
  INV_X1    g617(.A(G2090), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n974), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n980), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1034), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G303), .A2(G8), .ZN(new_n1050));
  XOR2_X1   g625(.A(new_n1050), .B(KEYINPUT55), .Z(new_n1051));
  NAND3_X1  g626(.A1(new_n1034), .A2(new_n1046), .A3(KEYINPUT114), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1049), .A2(new_n1051), .A3(G8), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1016), .B1(new_n1030), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1032), .A2(new_n980), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n701), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(G2084), .B1(new_n974), .B2(new_n1044), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(new_n1042), .A3(new_n980), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n998), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G168), .A2(new_n998), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(KEYINPUT122), .B2(KEYINPUT51), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1056), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1056), .ZN(new_n1067));
  INV_X1    g642(.A(new_n979), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n470), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n1041), .B2(KEYINPUT50), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n701), .A2(new_n1033), .B1(new_n1070), .B2(new_n1060), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1064), .B(new_n1067), .C1(new_n1071), .C2(new_n998), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1063), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1066), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT62), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1066), .A2(new_n1072), .A3(new_n1077), .A4(new_n1074), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1961), .B1(new_n1070), .B2(new_n1045), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1033), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n720), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(KEYINPUT53), .A3(new_n720), .ZN(new_n1084));
  AOI21_X1  g659(.A(G301), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1076), .A2(new_n1078), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n980), .B1(new_n974), .B2(new_n1044), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT118), .B(new_n980), .C1(new_n974), .C2(new_n1044), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1045), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1034), .B1(new_n1091), .B2(G2090), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G8), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1050), .B(KEYINPUT55), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1053), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1055), .B1(new_n1086), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1071), .A2(new_n998), .A3(G286), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1095), .A2(new_n1053), .A3(new_n1096), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1052), .A2(G8), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT114), .B1(new_n1034), .B2(new_n1046), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1094), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR4_X1   g679(.A1(new_n1071), .A2(new_n1099), .A3(new_n998), .A4(G286), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n1053), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1099), .A2(new_n1101), .B1(new_n1106), .B2(new_n1030), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1098), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  XNOR2_X1  g684(.A(G299), .B(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT120), .Z(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1091), .A2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT56), .B(G2072), .Z(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(new_n1033), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1032), .A2(new_n980), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1041), .A2(new_n976), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1114), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1113), .A2(new_n1121), .A3(new_n1110), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1041), .A2(KEYINPUT50), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n731), .B1(new_n1125), .B2(new_n1087), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n974), .A2(new_n980), .A3(new_n969), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n597), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1111), .A2(new_n1123), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT121), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n606), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(KEYINPUT121), .A3(new_n597), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1130), .A2(KEYINPUT121), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1134), .A2(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1110), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1124), .B1(new_n1139), .B2(KEYINPUT61), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1122), .A2(new_n1141), .A3(new_n1110), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1033), .A2(G1996), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT58), .B(G1341), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n974), .B2(new_n980), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n549), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT59), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1140), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1129), .B1(new_n1138), .B2(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1095), .A2(new_n1053), .A3(new_n1096), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n1152));
  XNOR2_X1  g727(.A(G171), .B(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n978), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1057), .A2(new_n1082), .A3(G2078), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1151), .A2(new_n1153), .B1(new_n1156), .B2(new_n1083), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1157), .A2(new_n1075), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1149), .A2(new_n1150), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n994), .B1(new_n1108), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT46), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n985), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT125), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT47), .ZN(new_n1164));
  INV_X1    g739(.A(new_n985), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n982), .A2(new_n973), .B1(new_n1165), .B2(KEYINPUT46), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n983), .A2(new_n984), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n986), .A2(new_n987), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n990), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n981), .A2(G1986), .A3(G290), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT48), .Z(new_n1177));
  NAND3_X1  g752(.A1(new_n1171), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n802), .A2(new_n805), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT123), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n988), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n1182), .A3(new_n970), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n982), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n988), .A2(new_n1180), .B1(new_n969), .B2(new_n876), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1185), .A2(new_n1182), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1170), .B(new_n1178), .C1(new_n1184), .C2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n967), .B1(new_n1160), .B2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1150), .A2(new_n1076), .A3(new_n1078), .A4(new_n1085), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1101), .A2(new_n1099), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1106), .A2(new_n1030), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1189), .B(new_n1055), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1150), .A2(new_n1075), .A3(new_n1157), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1133), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n597), .B1(new_n1130), .B2(KEYINPUT121), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1135), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1137), .A2(new_n1136), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1198), .A2(new_n1142), .A3(new_n1140), .A4(new_n1147), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1193), .B1(new_n1199), .B2(new_n1129), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n993), .B1(new_n1192), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1174), .B1(new_n988), .B2(new_n990), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1202), .A2(new_n1203), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1186), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n981), .B1(new_n1185), .B2(new_n1182), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1201), .A2(KEYINPUT127), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1188), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g784(.A1(new_n960), .A2(new_n964), .A3(new_n961), .ZN(new_n1211));
  INV_X1    g785(.A(new_n456), .ZN(new_n1212));
  OR2_X1    g786(.A1(G227), .A2(new_n1212), .ZN(new_n1213));
  NOR3_X1   g787(.A1(G229), .A2(G401), .A3(new_n1213), .ZN(new_n1214));
  AND3_X1   g788(.A1(new_n1211), .A2(new_n1214), .A3(new_n897), .ZN(G308));
  NAND3_X1  g789(.A1(new_n1211), .A2(new_n1214), .A3(new_n897), .ZN(G225));
endmodule


