//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(new_n203), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n211), .B1(new_n215), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(KEYINPUT67), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT67), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G1), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n248), .A2(new_n250), .A3(G13), .A4(G20), .ZN(new_n251));
  AND2_X1   g0051(.A1(new_n248), .A2(new_n250), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n212), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  MUX2_X1   g0057(.A(new_n251), .B(new_n257), .S(G50), .Z(new_n258));
  NOR3_X1   g0058(.A1(new_n202), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(KEYINPUT69), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n213), .A3(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n255), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  OR2_X1    g0068(.A1(G41), .A2(G45), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(new_n248), .A3(new_n250), .ZN(new_n270));
  INV_X1    g0070(.A(new_n212), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT68), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT68), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n270), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT66), .B(G226), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n271), .B2(new_n272), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n247), .A3(new_n269), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(G222), .A2(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(G223), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n273), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT3), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n219), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n285), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n281), .A2(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n267), .A2(new_n268), .B1(new_n298), .B2(G200), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n299), .B1(new_n268), .B2(new_n267), .C1(new_n300), .C2(new_n298), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n267), .C1(G179), .C2(new_n298), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n251), .A2(new_n256), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT70), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT70), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n251), .A2(new_n256), .A3(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n311), .A2(new_n253), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G77), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G20), .A2(G77), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n213), .A2(new_n291), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n213), .A2(G33), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n316), .B1(new_n260), .B2(new_n317), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n251), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n320), .A2(new_n255), .B1(new_n219), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n278), .A2(G244), .ZN(new_n325));
  NOR2_X1   g0125(.A1(G232), .A2(G1698), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n287), .A2(G238), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n289), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n273), .B1(new_n295), .B2(new_n221), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n285), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT71), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n324), .A2(KEYINPUT71), .A3(new_n332), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n335), .B(new_n336), .C1(new_n300), .C2(new_n331), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n331), .A2(new_n305), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n325), .A2(new_n339), .A3(new_n330), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n323), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n309), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n314), .A2(G68), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n321), .A2(new_n203), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT12), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT75), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n263), .A2(G50), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT74), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n348), .B(new_n349), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n318), .A2(new_n219), .B1(new_n213), .B2(G68), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n255), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT11), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n352), .B(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n346), .B2(KEYINPUT75), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n347), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT14), .ZN(new_n358));
  AND3_X1   g0158(.A1(new_n270), .A2(new_n276), .A3(new_n273), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n276), .B1(new_n270), .B2(new_n273), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT73), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT73), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n275), .A2(new_n362), .A3(new_n277), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n363), .A3(G238), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n287), .A2(G226), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT72), .B1(new_n295), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT72), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n289), .A2(new_n368), .A3(G226), .A4(new_n287), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G97), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n289), .A2(G232), .A3(G1698), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n367), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n273), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n285), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n364), .A2(new_n365), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n365), .B1(new_n364), .B2(new_n374), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n358), .B(G169), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT77), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n364), .A2(new_n374), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT13), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n364), .A2(new_n365), .A3(new_n374), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n383), .A2(KEYINPUT77), .A3(new_n358), .A4(G169), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n375), .A2(new_n376), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G179), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n305), .B1(new_n381), .B2(new_n382), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n389), .A2(KEYINPUT76), .A3(new_n358), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT76), .ZN(new_n391));
  OAI21_X1  g0191(.A(G169), .B1(new_n375), .B2(new_n376), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(KEYINPUT14), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n357), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n383), .A2(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n386), .A2(G190), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n356), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G58), .A2(G68), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n213), .B1(new_n216), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G159), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n317), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT80), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT80), .B1(new_n401), .B2(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n293), .A2(KEYINPUT79), .A3(G33), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT79), .B1(new_n293), .B2(G33), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT78), .B1(new_n293), .B2(G33), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT78), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(new_n291), .A3(KEYINPUT3), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n409), .B(new_n213), .C1(new_n412), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G68), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n413), .B(new_n415), .C1(new_n410), .C2(new_n411), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n409), .B1(new_n419), .B2(new_n213), .ZN(new_n420));
  OAI211_X1 g0220(.A(KEYINPUT16), .B(new_n408), .C1(new_n418), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT16), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n409), .B1(new_n289), .B2(G20), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n295), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n203), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n404), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n421), .A2(new_n255), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n257), .A2(new_n261), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n321), .B2(new_n261), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n413), .A2(new_n415), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT79), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n291), .B2(KEYINPUT3), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n293), .A2(KEYINPUT79), .A3(G33), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  MUX2_X1   g0235(.A(G223), .B(G226), .S(G1698), .Z(new_n436));
  NAND3_X1  g0236(.A1(new_n431), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G87), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n373), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n284), .B1(new_n274), .B2(new_n231), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n442), .A3(new_n300), .ZN(new_n443));
  INV_X1    g0243(.A(G200), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n273), .B1(new_n437), .B2(new_n438), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n441), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n428), .A2(new_n430), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n428), .A2(new_n447), .A3(KEYINPUT17), .A4(new_n430), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT82), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n440), .A2(new_n442), .A3(G179), .ZN(new_n454));
  OAI21_X1  g0254(.A(G169), .B1(new_n445), .B2(new_n441), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT81), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n454), .B2(new_n455), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n428), .A2(new_n430), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT18), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n452), .B1(new_n453), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT18), .ZN(new_n463));
  INV_X1    g0263(.A(new_n460), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n305), .B1(new_n440), .B2(new_n442), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n445), .A2(new_n339), .A3(new_n441), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT81), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n454), .A2(new_n456), .A3(new_n455), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n463), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n459), .A2(KEYINPUT18), .A3(new_n460), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT82), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n462), .A2(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n342), .A2(new_n399), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT19), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n213), .B1(new_n370), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G87), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n221), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n476), .A2(new_n479), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n435), .A2(new_n213), .A3(new_n413), .A4(new_n415), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n203), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n255), .ZN(new_n484));
  INV_X1    g0284(.A(new_n319), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(new_n251), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n248), .A2(new_n250), .A3(G33), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n310), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n485), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n484), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G238), .A2(G1698), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n220), .B2(G1698), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n435), .A2(new_n493), .A3(new_n413), .A4(new_n415), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G116), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n273), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n248), .A2(new_n250), .A3(G45), .ZN(new_n497));
  INV_X1    g0297(.A(G250), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n248), .A2(new_n250), .A3(G45), .A4(new_n282), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n273), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n305), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n494), .A2(new_n495), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n373), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n339), .A3(new_n501), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n491), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(G190), .A3(new_n501), .ZN(new_n508));
  OAI21_X1  g0308(.A(G200), .B1(new_n496), .B2(new_n502), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n486), .B1(new_n483), .B2(new_n255), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n310), .A2(new_n488), .A3(new_n477), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n508), .A2(new_n509), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n507), .A2(new_n513), .A3(KEYINPUT86), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT86), .B1(new_n507), .B2(new_n513), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(KEYINPUT5), .A2(G41), .ZN(new_n518));
  NOR2_X1   g0318(.A1(KEYINPUT5), .A2(G41), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n252), .A2(new_n520), .A3(new_n283), .A4(G45), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  OAI211_X1 g0322(.A(G257), .B(new_n273), .C1(new_n497), .C2(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G283), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G250), .A2(G1698), .ZN(new_n526));
  NAND2_X1  g0326(.A1(KEYINPUT4), .A2(G244), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(G1698), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n525), .B1(new_n529), .B2(new_n295), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n431), .A2(G244), .A3(new_n287), .A4(new_n435), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n524), .B1(new_n533), .B2(new_n273), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n535), .A2(new_n478), .A3(G107), .ZN(new_n536));
  XNOR2_X1  g0336(.A(G97), .B(G107), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n538), .A2(new_n213), .B1(new_n219), .B2(new_n317), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n221), .B1(new_n423), .B2(new_n424), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n255), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n251), .A2(G97), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n489), .B2(G97), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n534), .A2(new_n305), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n339), .B(new_n524), .C1(new_n533), .C2(new_n273), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n545), .A2(KEYINPUT83), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(KEYINPUT83), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT84), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n435), .A2(new_n287), .A3(new_n413), .A4(new_n415), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n532), .B1(new_n551), .B2(new_n220), .ZN(new_n552));
  INV_X1    g0352(.A(new_n530), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n373), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT83), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n339), .A4(new_n524), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n545), .A2(KEYINPUT83), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(KEYINPUT84), .A3(new_n544), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n534), .A2(G200), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n541), .A2(new_n543), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n300), .C2(new_n534), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n550), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT85), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n550), .A2(KEYINPUT85), .A3(new_n560), .A4(new_n563), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n517), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G264), .B(new_n273), .C1(new_n497), .C2(new_n522), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G294), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G250), .A2(G1698), .ZN(new_n572));
  INV_X1    g0372(.A(G257), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(G1698), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n571), .B1(new_n419), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n570), .B1(new_n576), .B2(new_n373), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n521), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n305), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n431), .A2(new_n435), .A3(new_n574), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n273), .B1(new_n580), .B2(new_n571), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n273), .A2(G274), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n582), .A2(new_n497), .A3(new_n522), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n581), .A2(new_n583), .A3(new_n570), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n339), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n477), .A2(G20), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT22), .B1(new_n289), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n221), .A2(KEYINPUT23), .A3(G20), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT23), .B1(new_n221), .B2(G20), .ZN(new_n590));
  INV_X1    g0390(.A(G116), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n589), .A2(new_n590), .B1(new_n591), .B2(new_n318), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(KEYINPUT22), .A2(G87), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n431), .A2(new_n213), .A3(new_n435), .A4(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n586), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(new_n586), .A3(new_n595), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n256), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n321), .A2(KEYINPUT25), .A3(new_n221), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT25), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n251), .B2(G107), .ZN(new_n602));
  AOI22_X1  g0402(.A1(G107), .A2(new_n489), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n579), .B(new_n585), .C1(new_n599), .C2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n593), .A2(new_n586), .A3(new_n595), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n255), .B1(new_n606), .B2(new_n596), .ZN(new_n607));
  AOI21_X1  g0407(.A(G200), .B1(new_n577), .B2(new_n521), .ZN(new_n608));
  NOR4_X1   g0408(.A1(new_n581), .A2(G190), .A3(new_n570), .A4(new_n583), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n607), .B(new_n603), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT87), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n222), .A2(new_n287), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n419), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n295), .A2(G303), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n431), .A2(G257), .A3(new_n287), .A4(new_n435), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n431), .A2(KEYINPUT87), .A3(new_n435), .A4(new_n614), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n373), .ZN(new_n621));
  OAI211_X1 g0421(.A(G270), .B(new_n273), .C1(new_n497), .C2(new_n522), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n521), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n254), .A2(new_n212), .B1(G20), .B2(new_n591), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n525), .B(new_n213), .C1(G33), .C2(new_n478), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(KEYINPUT20), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT20), .B1(new_n626), .B2(new_n627), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n629), .A2(new_n630), .B1(G116), .B2(new_n251), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n488), .A2(new_n591), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n311), .A2(new_n313), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n305), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n625), .A2(KEYINPUT21), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n623), .B1(new_n620), .B2(new_n373), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n311), .A2(new_n313), .A3(new_n633), .ZN(new_n639));
  OAI21_X1  g0439(.A(G169), .B1(new_n639), .B2(new_n631), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n632), .A2(new_n634), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n638), .A2(G179), .A3(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n636), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n642), .B1(new_n625), .B2(G200), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n300), .B2(new_n625), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n474), .A2(new_n568), .A3(new_n612), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n379), .A2(new_n384), .B1(G179), .B2(new_n386), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT76), .B1(new_n389), .B2(new_n358), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n392), .A2(new_n391), .A3(KEYINPUT14), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n356), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n341), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n398), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n649), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n395), .A2(KEYINPUT89), .A3(new_n656), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n450), .A2(new_n451), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n454), .A2(new_n455), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n460), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(new_n463), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n304), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n308), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n507), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n550), .A2(new_n560), .A3(new_n563), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n509), .A2(KEYINPUT88), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n431), .A2(new_n213), .A3(G68), .A4(new_n435), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n256), .B1(new_n671), .B2(new_n481), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n672), .A2(new_n486), .A3(new_n511), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT88), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n674), .B(G200), .C1(new_n496), .C2(new_n502), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n670), .A2(new_n508), .A3(new_n673), .A4(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n610), .A2(new_n507), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n644), .B2(new_n605), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n668), .B1(new_n669), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n507), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n548), .A2(new_n680), .A3(KEYINPUT26), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n559), .A2(KEYINPUT84), .A3(new_n544), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT84), .B1(new_n559), .B2(new_n544), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n516), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n681), .B1(new_n684), .B2(KEYINPUT26), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n474), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n667), .A2(new_n687), .ZN(G369));
  AND2_X1   g0488(.A1(new_n213), .A2(G13), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n252), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n642), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n647), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n636), .A2(new_n641), .A3(new_n643), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(new_n642), .A3(new_n695), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT90), .A3(G330), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT90), .B1(new_n700), .B2(G330), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n695), .B1(new_n599), .B2(new_n604), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n612), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n605), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n695), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n704), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n695), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n698), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n611), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n707), .B2(new_n711), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(G399));
  AOI21_X1  g0515(.A(new_n695), .B1(new_n679), .B2(new_n685), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT26), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n548), .A2(new_n680), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n684), .B2(new_n718), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n605), .A2(new_n641), .A3(new_n643), .A4(new_n636), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n610), .A2(new_n507), .A3(new_n676), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n507), .B1(new_n564), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n711), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT91), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT91), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n727), .B(new_n711), .C1(new_n720), .C2(new_n724), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n717), .B1(new_n729), .B2(KEYINPUT29), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n612), .A2(new_n644), .A3(new_n646), .A4(new_n711), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n682), .A2(new_n683), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT85), .B1(new_n733), .B2(new_n563), .ZN(new_n734));
  INV_X1    g0534(.A(new_n567), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n516), .B(new_n732), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n638), .A2(G179), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n496), .A2(new_n502), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n555), .A2(new_n738), .A3(new_n524), .A4(new_n577), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  OR3_X1    g0540(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n584), .A2(G179), .A3(new_n738), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n534), .A3(new_n625), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n740), .B1(new_n737), .B2(new_n739), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT31), .B1(new_n745), .B2(new_n695), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n736), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n730), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT92), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(new_n247), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n209), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G41), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n479), .A2(G116), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n760), .A2(G1), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(new_n217), .B2(new_n760), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n764), .ZN(G364));
  AOI21_X1  g0565(.A(new_n247), .B1(new_n689), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n759), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n704), .B(new_n769), .C1(G330), .C2(new_n700), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n212), .B1(G20), .B2(new_n305), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n245), .A2(G45), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT93), .Z(new_n778));
  INV_X1    g0578(.A(new_n419), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n758), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n778), .B(new_n780), .C1(G45), .C2(new_n217), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n758), .A2(new_n295), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n782), .A2(G355), .B1(new_n591), .B2(new_n758), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n776), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n774), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n213), .A2(new_n339), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(new_n444), .A3(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n787), .A2(new_n300), .A3(new_n444), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n789), .A2(new_n203), .B1(new_n791), .B2(new_n201), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n792), .B1(G77), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n213), .A2(G179), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(new_n300), .A3(G200), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT94), .Z(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G107), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n797), .A2(new_n793), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n801), .A2(KEYINPUT32), .A3(new_n402), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n300), .A2(G179), .A3(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n213), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n478), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n802), .B(new_n805), .C1(G87), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT32), .ZN(new_n809));
  INV_X1    g0609(.A(new_n801), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(G159), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n787), .A2(new_n300), .A3(G200), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n295), .B(new_n811), .C1(G58), .C2(new_n812), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n796), .A2(new_n800), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n812), .A2(G322), .B1(G329), .B2(new_n810), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT95), .B(G326), .Z(new_n816));
  NAND2_X1  g0616(.A1(new_n790), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(KEYINPUT33), .A2(G317), .ZN(new_n818));
  AND2_X1   g0618(.A1(KEYINPUT33), .A2(G317), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n788), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n815), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  INV_X1    g0622(.A(G294), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n295), .B1(new_n794), .B2(new_n822), .C1(new_n804), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G303), .B2(new_n807), .ZN(new_n825));
  INV_X1    g0625(.A(G283), .ZN(new_n826));
  INV_X1    g0626(.A(new_n799), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n821), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n785), .B1(new_n814), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n784), .A2(new_n829), .A3(new_n769), .ZN(new_n830));
  INV_X1    g0630(.A(new_n773), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n700), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n770), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NOR2_X1   g0634(.A1(new_n341), .A2(new_n695), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n323), .A2(new_n695), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n337), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n835), .B1(new_n837), .B2(new_n341), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n716), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n686), .A2(new_n711), .A3(new_n838), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n768), .B1(new_n841), .B2(new_n750), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n750), .B2(new_n841), .ZN(new_n843));
  INV_X1    g0643(.A(new_n812), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n826), .A2(new_n789), .B1(new_n844), .B2(new_n823), .ZN(new_n845));
  INV_X1    g0645(.A(G303), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n791), .A2(new_n846), .B1(new_n801), .B2(new_n822), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n289), .B(new_n805), .C1(G116), .C2(new_n795), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n799), .A2(G87), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n807), .A2(G107), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n788), .A2(G150), .B1(G159), .B2(new_n795), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  INV_X1    g0654(.A(G143), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n854), .B2(new_n791), .C1(new_n855), .C2(new_n844), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT34), .Z(new_n857));
  NAND2_X1  g0657(.A1(new_n799), .A2(G68), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n419), .B1(G132), .B2(new_n810), .ZN(new_n859));
  INV_X1    g0659(.A(new_n804), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n860), .A2(G58), .B1(new_n807), .B2(G50), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n852), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n774), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n774), .A2(new_n771), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n769), .B1(new_n219), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n864), .B(new_n866), .C1(new_n838), .C2(new_n772), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n843), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(G384));
  INV_X1    g0669(.A(new_n538), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n591), .B(new_n215), .C1(new_n870), .C2(KEYINPUT35), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(KEYINPUT35), .B2(new_n870), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT36), .Z(new_n873));
  NAND2_X1  g0673(.A1(new_n400), .A2(G77), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n217), .A2(new_n874), .B1(G50), .B2(new_n203), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n252), .A2(G13), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n421), .A2(new_n255), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n419), .A2(new_n213), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT7), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(G68), .A3(new_n417), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT16), .B1(new_n881), .B2(new_n408), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n430), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n693), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT82), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n453), .B(new_n463), .C1(new_n464), .C2(new_n469), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n660), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n886), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n883), .A2(new_n662), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n885), .A3(new_n448), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n460), .A2(new_n884), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(new_n448), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT37), .B1(new_n459), .B2(new_n460), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n890), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n894), .B1(new_n664), .B2(new_n660), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n663), .A2(new_n894), .A3(new_n448), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n895), .A2(new_n896), .B1(new_n903), .B2(KEYINPUT37), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n901), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n899), .A2(new_n900), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT99), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n885), .B1(new_n462), .B2(new_n472), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n893), .A2(new_n897), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n908), .A2(new_n909), .A3(new_n901), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n890), .B2(new_n898), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT39), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT99), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n899), .A2(new_n905), .A3(new_n913), .A4(new_n900), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT98), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n395), .B2(new_n695), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n654), .A2(KEYINPUT98), .A3(new_n711), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n835), .B(KEYINPUT96), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n840), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n901), .B1(new_n908), .B2(new_n909), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n899), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n650), .A2(new_n653), .A3(new_n398), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n356), .A2(new_n711), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT97), .ZN(new_n929));
  INV_X1    g0729(.A(new_n927), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n395), .A2(new_n398), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT97), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(new_n932), .A3(new_n927), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n929), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n923), .A2(new_n925), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n664), .A2(new_n884), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n920), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n729), .A2(KEYINPUT29), .ZN(new_n938));
  INV_X1    g0738(.A(new_n717), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n474), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n667), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n937), .B(new_n941), .Z(new_n942));
  NAND2_X1  g0742(.A1(new_n837), .A2(new_n341), .ZN(new_n943));
  INV_X1    g0743(.A(new_n835), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n736), .B2(new_n748), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n934), .A2(new_n925), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n899), .A2(new_n905), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n934), .A2(new_n946), .A3(new_n950), .A4(KEYINPUT40), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n474), .A2(new_n749), .ZN(new_n953));
  OAI21_X1  g0753(.A(G330), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n942), .A2(new_n955), .B1(new_n252), .B2(new_n689), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n942), .A2(new_n955), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n877), .B1(new_n956), .B2(new_n957), .ZN(G367));
  INV_X1    g0758(.A(new_n780), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n775), .B1(new_n209), .B2(new_n319), .C1(new_n959), .C2(new_n237), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n768), .ZN(new_n961));
  INV_X1    g0761(.A(G150), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n844), .A2(new_n962), .B1(new_n791), .B2(new_n855), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n804), .A2(new_n203), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(KEYINPUT106), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT107), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n289), .B1(new_n798), .B2(new_n219), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n967), .B2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n965), .A2(KEYINPUT106), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n789), .A2(new_n402), .B1(new_n801), .B2(new_n854), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G50), .B2(new_n795), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n971), .B(new_n973), .C1(new_n202), .C2(new_n806), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n806), .A2(new_n591), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT46), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G294), .A2(new_n788), .B1(new_n812), .B2(G303), .ZN(new_n977));
  INV_X1    g0777(.A(new_n798), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n860), .A2(G107), .B1(new_n978), .B2(G97), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n977), .A2(new_n419), .A3(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n790), .A2(G311), .B1(G317), .B2(new_n810), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(new_n826), .C2(new_n794), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n970), .A2(new_n974), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n961), .B1(new_n984), .B2(new_n774), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n711), .A2(new_n673), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n680), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n668), .B2(new_n986), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT100), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n773), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n548), .A2(new_n711), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT101), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n711), .A2(new_n562), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n564), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n709), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n550), .A2(new_n560), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n995), .B2(new_n707), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n695), .B1(new_n999), .B2(KEYINPUT102), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT102), .B2(new_n999), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n995), .A2(new_n713), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT42), .Z(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT103), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n989), .B(KEYINPUT43), .Z(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(new_n989), .C2(new_n1004), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1006), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(KEYINPUT103), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n997), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1007), .A2(new_n997), .A3(new_n1009), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n995), .A2(new_n714), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n1015));
  XOR2_X1   g0815(.A(new_n1014), .B(new_n1015), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n995), .A2(new_n714), .ZN(new_n1017));
  XOR2_X1   g0817(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(new_n709), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n706), .A2(new_n708), .A3(new_n712), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n611), .B2(new_n712), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n704), .B(new_n1023), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n756), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1021), .A2(new_n1025), .B1(new_n1026), .B2(new_n754), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n759), .B(KEYINPUT41), .Z(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n767), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n991), .B1(new_n1013), .B2(new_n1030), .ZN(G387));
  NAND3_X1  g0831(.A1(new_n755), .A2(new_n1025), .A3(new_n756), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT110), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1024), .B1(new_n1026), .B2(new_n754), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n755), .A2(new_n1025), .A3(KEYINPUT110), .A4(new_n756), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1034), .A2(new_n759), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n1025), .A2(KEYINPUT108), .A3(new_n766), .ZN(new_n1038));
  OAI21_X1  g0838(.A(KEYINPUT108), .B1(new_n1025), .B2(new_n766), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n706), .A2(new_n708), .A3(new_n773), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n812), .A2(G317), .B1(new_n790), .B2(G322), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n788), .A2(G311), .B1(G303), .B2(new_n795), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1043), .A2(KEYINPUT48), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(KEYINPUT48), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n804), .A2(new_n826), .B1(new_n806), .B2(new_n823), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1047), .A2(KEYINPUT49), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(KEYINPUT49), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n798), .A2(new_n591), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1050), .B(new_n779), .C1(new_n816), .C2(new_n810), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G68), .A2(new_n795), .B1(new_n810), .B2(G150), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n791), .B2(new_n402), .C1(new_n201), .C2(new_n844), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n261), .B2(new_n788), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n804), .A2(new_n319), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n806), .A2(new_n219), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1056), .A2(new_n1057), .A3(new_n419), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1055), .B(new_n1058), .C1(new_n478), .C2(new_n827), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n785), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n234), .A2(G45), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT109), .Z(new_n1062));
  NOR2_X1   g0862(.A1(new_n260), .A2(G50), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT50), .Z(new_n1064));
  AOI21_X1  g0864(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n761), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1062), .B(new_n780), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n761), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n782), .A2(new_n1068), .B1(new_n221), .B2(new_n758), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n776), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1060), .A2(new_n769), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1038), .A2(new_n1039), .B1(new_n1040), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1037), .A2(new_n1072), .ZN(G393));
  XNOR2_X1  g0873(.A(new_n1020), .B(new_n710), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n767), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n775), .B1(new_n478), .B2(new_n209), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n242), .B2(new_n780), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n812), .A2(G159), .B1(new_n790), .B2(G150), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT51), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n794), .A2(new_n260), .B1(new_n801), .B2(new_n855), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G50), .B2(new_n788), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n779), .B1(new_n203), .B2(new_n806), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G77), .B2(new_n860), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1079), .A2(new_n850), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n289), .B1(new_n810), .B2(G322), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n800), .B(new_n1085), .C1(new_n826), .C2(new_n806), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT112), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n812), .A2(G311), .B1(new_n790), .B2(G317), .ZN(new_n1088));
  XOR2_X1   g0888(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n1089));
  AND2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n788), .A2(G303), .B1(G294), .B2(new_n795), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n591), .B2(new_n804), .ZN(new_n1093));
  OR3_X1    g0893(.A1(new_n1090), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1084), .B1(new_n1087), .B2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n769), .B(new_n1077), .C1(new_n1095), .C2(new_n774), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n995), .B2(new_n831), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1074), .B(new_n1024), .C1(new_n1026), .C2(new_n754), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n759), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1035), .A2(new_n1021), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1075), .B(new_n1097), .C1(new_n1099), .C2(new_n1101), .ZN(G390));
  NAND3_X1  g0902(.A1(new_n934), .A2(new_n946), .A3(G330), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n919), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n950), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n678), .A2(new_n733), .A3(new_n563), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT26), .B1(new_n998), .B2(new_n516), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n507), .C1(new_n1108), .C2(new_n719), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n727), .B1(new_n1109), .B2(new_n711), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n728), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n838), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n922), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1106), .B1(new_n1113), .B2(new_n934), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n919), .B1(new_n923), .B2(new_n934), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n915), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1104), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n921), .B1(new_n729), .B2(new_n838), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n929), .A2(new_n931), .A3(new_n933), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1105), .B(new_n950), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n921), .B1(new_n716), .B2(new_n838), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1105), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1122), .A2(new_n907), .A3(new_n912), .A4(new_n914), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1120), .A2(new_n1123), .A3(new_n1103), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1117), .A2(new_n767), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n865), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n768), .B1(new_n261), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n794), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G132), .ZN(new_n1130));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n844), .A2(new_n1130), .B1(new_n791), .B2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1129), .B(new_n1132), .C1(G125), .C2(new_n810), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n806), .A2(new_n962), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n978), .A2(G50), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n289), .B1(new_n789), .B2(new_n854), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G159), .B2(new_n860), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n844), .A2(new_n591), .B1(new_n791), .B2(new_n826), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G77), .B2(new_n860), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n794), .A2(new_n478), .B1(new_n801), .B2(new_n823), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G107), .B2(new_n788), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n858), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n295), .B1(new_n806), .B2(new_n477), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT114), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1139), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1127), .B1(new_n1147), .B2(new_n774), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n915), .B2(new_n772), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1125), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n751), .A2(new_n474), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n940), .A2(new_n667), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n517), .B(new_n731), .C1(new_n566), .C2(new_n567), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n746), .A2(new_n747), .ZN(new_n1156));
  OAI211_X1 g0956(.A(G330), .B(new_n838), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1119), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1103), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n923), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1118), .A2(new_n1103), .A3(new_n1158), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1117), .A2(new_n1124), .A3(new_n1154), .A4(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1163), .A2(KEYINPUT113), .A3(new_n759), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1154), .A2(new_n1162), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT113), .B1(new_n1163), .B2(new_n759), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1151), .B1(new_n1168), .B2(new_n1169), .ZN(G378));
  NAND2_X1  g0970(.A1(new_n1163), .A2(new_n1154), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT115), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n947), .A2(new_n948), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n951), .A2(G330), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n949), .A2(KEYINPUT115), .A3(G330), .A4(new_n951), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n267), .A2(new_n884), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n309), .A2(new_n1177), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n309), .A2(new_n1177), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1179), .B2(new_n1178), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1175), .A2(new_n1176), .A3(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1172), .B1(new_n1181), .B2(new_n1182), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n937), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n937), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1184), .A2(new_n1188), .A3(new_n1185), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1171), .A2(new_n1187), .A3(KEYINPUT57), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n759), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1184), .A2(new_n1188), .A3(new_n1185), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1188), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1171), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1187), .A2(new_n767), .A3(new_n1189), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1183), .A2(new_n771), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n769), .B1(new_n201), .B2(new_n865), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n788), .A2(G132), .B1(new_n790), .B2(G125), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n1131), .B2(new_n844), .C1(new_n854), .C2(new_n794), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n804), .A2(new_n962), .B1(new_n806), .B2(new_n1128), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n978), .A2(G159), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n810), .C2(G124), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n779), .A2(G41), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n790), .A2(G116), .B1(new_n485), .B2(new_n795), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(new_n478), .C2(new_n789), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n844), .A2(new_n221), .B1(new_n801), .B2(new_n826), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n798), .A2(new_n202), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1057), .A2(new_n1214), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n1212), .A2(new_n964), .A3(new_n1213), .A4(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1210), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1220));
  AND4_X1   g1020(.A1(new_n1209), .A2(new_n1217), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1198), .B(new_n1199), .C1(new_n785), .C2(new_n1221), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1197), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1196), .A2(new_n1223), .ZN(G375));
  NAND3_X1  g1024(.A1(new_n1153), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1166), .A2(new_n1029), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1119), .A2(new_n771), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT116), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n790), .A2(G294), .B1(G107), .B2(new_n795), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n591), .B2(new_n789), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT117), .Z(new_n1231));
  OAI22_X1  g1031(.A1(new_n806), .A2(new_n478), .B1(new_n801), .B2(new_n846), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT118), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n289), .B(new_n1056), .C1(G283), .C2(new_n812), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n219), .B2(new_n827), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1231), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n806), .A2(new_n402), .B1(new_n801), .B2(new_n1131), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT120), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n419), .B1(G150), .B2(new_n795), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1214), .B1(G50), .B2(new_n860), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT121), .Z(new_n1242));
  OAI22_X1  g1042(.A1(new_n854), .A2(new_n844), .B1(new_n789), .B2(new_n1128), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT119), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n791), .B2(new_n1130), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n790), .A2(KEYINPUT119), .A3(G132), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1243), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1236), .B1(new_n1242), .B2(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n768), .B1(G68), .B2(new_n1126), .C1(new_n1248), .C2(new_n785), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1162), .A2(new_n767), .B1(new_n1228), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1226), .A2(new_n1251), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT122), .Z(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(G381));
  NAND3_X1  g1054(.A1(new_n1037), .A2(new_n833), .A3(new_n1072), .ZN(new_n1255));
  NOR4_X1   g1055(.A1(G381), .A2(G384), .A3(G390), .A4(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(G375), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1012), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1258), .A2(new_n1010), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1074), .A2(new_n1024), .B1(new_n756), .B2(new_n755), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n766), .B1(new_n1260), .B2(new_n1028), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1259), .A2(new_n1261), .B1(new_n990), .B2(new_n985), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1169), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1150), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1256), .A2(new_n1257), .A3(new_n1262), .A4(new_n1265), .ZN(G407));
  NAND2_X1  g1066(.A1(new_n694), .A2(G213), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT123), .Z(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1196), .A2(new_n1265), .A3(new_n1223), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(new_n1269), .C2(new_n1270), .ZN(G409));
  OAI211_X1 g1071(.A(G378), .B(new_n1223), .C1(new_n1191), .C2(new_n1195), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1171), .A2(new_n1187), .A3(new_n1029), .A4(new_n1189), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1197), .A3(new_n1222), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1265), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1153), .A2(KEYINPUT60), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1121), .B1(new_n1158), .B2(new_n1103), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1158), .A2(new_n1103), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(new_n1118), .B2(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1282), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1153), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1279), .A2(new_n1283), .A3(new_n759), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT60), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1225), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT124), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1166), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT60), .B1(new_n1282), .B2(new_n1153), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1282), .A2(new_n1153), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT124), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1284), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1251), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n868), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1279), .A2(new_n1283), .A3(new_n759), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1289), .A2(new_n1290), .A3(KEYINPUT124), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1287), .B1(new_n1286), .B2(new_n1166), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(G384), .A3(new_n1251), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1276), .A2(new_n1269), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT62), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1276), .A2(new_n1269), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1268), .A2(G2897), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1294), .A2(new_n1299), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1294), .B2(new_n1299), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1276), .A2(new_n1311), .A3(new_n1269), .A4(new_n1301), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1303), .A2(new_n1309), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1075), .A2(new_n1097), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1099), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1315), .B2(new_n1100), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(G387), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1262), .A2(G390), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G393), .A2(G396), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1255), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1317), .A2(new_n1318), .A3(new_n1320), .A4(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT126), .B1(new_n1262), .B2(G390), .ZN(new_n1324));
  AOI22_X1  g1124(.A1(new_n1324), .A2(new_n1320), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1313), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT61), .B1(new_n1304), .B2(new_n1308), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1324), .A2(new_n1320), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1322), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1302), .A2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1276), .A2(KEYINPUT63), .A3(new_n1269), .A4(new_n1301), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1328), .A2(new_n1332), .A3(new_n1334), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1327), .A2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(G375), .A2(G378), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1270), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1301), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT127), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1338), .A2(new_n1270), .A3(new_n1300), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1340), .A2(new_n1326), .A3(new_n1341), .A4(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1331), .A2(new_n1341), .A3(new_n1322), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1338), .A2(new_n1270), .A3(new_n1300), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1300), .B1(new_n1338), .B2(new_n1270), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1344), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1326), .A2(new_n1341), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1343), .B1(new_n1347), .B2(new_n1348), .ZN(G402));
endmodule


