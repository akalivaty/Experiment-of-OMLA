//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n212), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n215), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  XNOR2_X1  g0043(.A(KEYINPUT8), .B(G58), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n209), .A2(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G150), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  OAI22_X1  g0048(.A1(new_n244), .A2(new_n245), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n249), .B1(G20), .B2(new_n203), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n208), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OR2_X1    g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n252), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n258), .A2(new_n261), .B1(new_n202), .B2(new_n257), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT9), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G222), .A2(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G223), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n269), .B(new_n272), .C1(G77), .C2(new_n265), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT65), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT65), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n279), .A2(new_n255), .A3(G274), .A4(new_n271), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n271), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G226), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n273), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G200), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT70), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n264), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n286), .A2(new_n287), .B1(new_n290), .B2(new_n285), .ZN(new_n291));
  OR3_X1    g0091(.A1(new_n289), .A2(KEYINPUT10), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT10), .B1(new_n289), .B2(new_n291), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n263), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n285), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT66), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n285), .A2(G179), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n297), .B2(KEYINPUT66), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT73), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT3), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(G33), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(G223), .A2(G1698), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G226), .B2(new_n267), .ZN(new_n311));
  INV_X1    g0111(.A(G87), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n309), .A2(new_n311), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT75), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI221_X1 g0115(.A(KEYINPUT75), .B1(new_n307), .B2(new_n312), .C1(new_n309), .C2(new_n311), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n272), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n283), .A2(G232), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n280), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(G179), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n271), .B1(new_n313), .B2(new_n314), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n319), .B1(new_n322), .B2(new_n316), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n321), .B1(new_n296), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G58), .ZN(new_n325));
  INV_X1    g0125(.A(G68), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(G20), .B1(new_n327), .B2(new_n201), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n247), .A2(G159), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT7), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n309), .A2(new_n332), .A3(new_n209), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G68), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n332), .B1(new_n309), .B2(new_n209), .ZN(new_n335));
  OAI211_X1 g0135(.A(KEYINPUT16), .B(new_n331), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT74), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT7), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n332), .A2(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n265), .B2(G20), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n306), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(new_n209), .A3(new_n340), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n326), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n337), .B1(new_n346), .B2(new_n330), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n336), .A2(new_n347), .A3(new_n252), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n244), .B1(new_n255), .B2(G20), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n258), .B1(new_n257), .B2(new_n244), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n324), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT18), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT17), .ZN(new_n354));
  AOI211_X1 g0154(.A(G190), .B(new_n319), .C1(new_n322), .C2(new_n316), .ZN(new_n355));
  AOI21_X1  g0155(.A(G200), .B1(new_n317), .B2(new_n320), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n354), .B1(new_n357), .B2(new_n351), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n348), .A2(new_n350), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n317), .A2(new_n290), .A3(new_n320), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G200), .B2(new_n323), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(KEYINPUT17), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT18), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n324), .A2(new_n351), .A3(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n353), .A2(new_n358), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n248), .A2(new_n202), .B1(new_n209), .B2(G68), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n245), .A2(new_n217), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n252), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n368), .B(KEYINPUT11), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n257), .A2(new_n326), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT12), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n258), .A2(G68), .A3(new_n259), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(KEYINPUT71), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT71), .B1(new_n371), .B2(new_n372), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT72), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G97), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n229), .A2(G1698), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G226), .B2(G1698), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n378), .B1(new_n380), .B2(new_n344), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n272), .B1(new_n283), .B2(G238), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n280), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT13), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(G169), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n384), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n385), .B1(new_n384), .B2(G169), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n377), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n376), .B1(new_n384), .B2(new_n290), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n384), .A2(G200), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT69), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n280), .B1(new_n218), .B2(new_n282), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n397), .A2(KEYINPUT67), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n265), .A2(G238), .A3(G1698), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n265), .A2(G232), .A3(new_n267), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n219), .C2(new_n265), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n272), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(KEYINPUT67), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n398), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n404), .B2(G179), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n403), .A2(new_n402), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n406), .A2(KEYINPUT69), .A3(new_n387), .A4(new_n398), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n258), .A2(G77), .A3(new_n259), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT68), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G20), .A2(G77), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT15), .B(G87), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n411), .B1(new_n244), .B2(new_n248), .C1(new_n245), .C2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n252), .B1(new_n217), .B2(new_n257), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n404), .A2(new_n296), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n410), .A2(new_n414), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n404), .B2(G200), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n290), .B2(new_n404), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n302), .A2(new_n365), .A3(new_n395), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT84), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n305), .A2(new_n308), .A3(new_n209), .A4(new_n306), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT22), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n312), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n312), .A2(G20), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT22), .B1(new_n265), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n422), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n308), .A2(new_n306), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n431), .A2(new_n209), .A3(new_n305), .A4(new_n425), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n265), .A2(new_n428), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n424), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(KEYINPUT84), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G116), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(G20), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT23), .B1(new_n219), .B2(G20), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n219), .A2(KEYINPUT23), .A3(G20), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT24), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n436), .A2(KEYINPUT24), .A3(new_n442), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n252), .ZN(new_n447));
  OR3_X1    g0247(.A1(new_n256), .A2(KEYINPUT25), .A3(G107), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT25), .B1(new_n256), .B2(G107), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n255), .A2(G33), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n256), .A2(new_n450), .A3(new_n208), .A4(new_n251), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n448), .B(new_n449), .C1(new_n219), .C2(new_n451), .ZN(new_n452));
  XOR2_X1   g0252(.A(new_n452), .B(KEYINPUT85), .Z(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT80), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT5), .B1(new_n276), .B2(new_n278), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n255), .A2(G45), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT5), .ZN(new_n460));
  AND2_X1   g0260(.A1(KEYINPUT65), .A2(G41), .ZN(new_n461));
  NOR2_X1   g0261(.A1(KEYINPUT65), .A2(G41), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n458), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(KEYINPUT80), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n460), .A2(G41), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G264), .A3(new_n271), .ZN(new_n469));
  INV_X1    g0269(.A(G250), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n267), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(G257), .B2(new_n267), .ZN(new_n472));
  INV_X1    g0272(.A(G294), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n309), .A2(new_n472), .B1(new_n307), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n272), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT86), .ZN(new_n476));
  INV_X1    g0276(.A(G274), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n272), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n459), .A2(new_n465), .A3(new_n478), .A4(new_n467), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(new_n480), .A3(new_n272), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n469), .A2(new_n476), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G169), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n469), .A2(new_n475), .A3(new_n479), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n387), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n455), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n253), .B1(new_n443), .B2(new_n444), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n453), .B1(new_n487), .B2(new_n446), .ZN(new_n488));
  INV_X1    g0288(.A(G200), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(G190), .B2(new_n482), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n219), .A2(G97), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g0296(.A(G97), .B(G107), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n496), .A2(KEYINPUT77), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OR3_X1    g0298(.A1(new_n494), .A2(KEYINPUT77), .A3(new_n495), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n209), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n342), .A2(new_n345), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n501), .A2(new_n219), .B1(new_n217), .B2(new_n248), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n252), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n257), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT78), .ZN(new_n506));
  INV_X1    g0306(.A(new_n451), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(G97), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n468), .A2(G257), .A3(new_n271), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n218), .A2(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n305), .A2(new_n308), .A3(new_n511), .A4(new_n306), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT4), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n343), .A2(new_n306), .A3(G250), .A4(G1698), .ZN(new_n515));
  AND2_X1   g0315(.A1(KEYINPUT4), .A2(G244), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n343), .A2(new_n306), .A3(new_n516), .A4(new_n267), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n272), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n510), .A2(new_n479), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n296), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n509), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT79), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(KEYINPUT79), .B(new_n272), .C1(new_n514), .C2(new_n519), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n463), .A2(new_n464), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n466), .B1(new_n528), .B2(new_n456), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n272), .B1(new_n529), .B2(new_n465), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n459), .A2(new_n465), .A3(new_n467), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n530), .A2(G257), .B1(new_n531), .B2(new_n478), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n527), .A2(new_n532), .A3(new_n387), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT81), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n527), .A2(new_n532), .A3(new_n535), .A4(new_n387), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n523), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n503), .B(new_n508), .C1(new_n290), .C2(new_n521), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n527), .A2(new_n532), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(G200), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n412), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(new_n256), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n451), .A2(new_n312), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT82), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT82), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT19), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n209), .A2(G33), .A3(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n312), .A2(new_n504), .A3(new_n219), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n378), .A2(new_n209), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(new_n546), .A4(new_n548), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n551), .B(new_n554), .C1(new_n423), .C2(new_n326), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n543), .B(new_n544), .C1(new_n555), .C2(new_n252), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G238), .A2(G1698), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n218), .B2(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n558), .A2(new_n306), .A3(new_n305), .A4(new_n308), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n271), .B1(new_n559), .B2(new_n437), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n458), .A2(new_n470), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n255), .A2(new_n477), .A3(G45), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n561), .A2(new_n271), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(G200), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n218), .A2(G1698), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(G238), .B2(G1698), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n437), .B1(new_n309), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n567), .B2(new_n272), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G190), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n556), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n555), .A2(new_n252), .ZN(new_n571));
  INV_X1    g0371(.A(new_n543), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n507), .A2(new_n542), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n296), .B1(new_n560), .B2(new_n563), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n568), .A2(new_n387), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n570), .A2(new_n577), .A3(KEYINPUT83), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT83), .B1(new_n570), .B2(new_n577), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n518), .B(new_n209), .C1(G33), .C2(new_n504), .ZN(new_n581));
  INV_X1    g0381(.A(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G20), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n252), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT20), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n256), .A2(G116), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n507), .B2(G116), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n296), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n468), .A2(G270), .A3(new_n271), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n220), .A2(G1698), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(G257), .B2(G1698), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n309), .A2(new_n593), .B1(new_n594), .B2(new_n265), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n272), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n479), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n589), .B(KEYINPUT21), .C1(new_n591), .C2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n479), .A2(new_n596), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n586), .A2(new_n588), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n599), .A2(G179), .A3(new_n600), .A4(new_n590), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n590), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT21), .B1(new_n603), .B2(new_n589), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n600), .B1(new_n603), .B2(G200), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n290), .B2(new_n603), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n580), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n421), .A2(new_n493), .A3(new_n541), .A4(new_n608), .ZN(G372));
  AND2_X1   g0409(.A1(new_n509), .A2(new_n522), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n510), .A2(new_n479), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n525), .B2(new_n526), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n535), .B1(new_n612), .B2(new_n387), .ZN(new_n613));
  INV_X1    g0413(.A(new_n536), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n567), .A2(new_n272), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT87), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT87), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n567), .A2(new_n618), .A3(new_n272), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n563), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n569), .B(new_n556), .C1(new_n620), .C2(new_n489), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n543), .B1(new_n555), .B2(new_n252), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(new_n573), .B1(new_n568), .B2(new_n387), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n620), .B2(G169), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n488), .B2(new_n491), .ZN(new_n626));
  INV_X1    g0426(.A(new_n509), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n539), .A2(G200), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n627), .B(new_n628), .C1(new_n290), .C2(new_n521), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n615), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n603), .A2(new_n589), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(KEYINPUT88), .A3(new_n598), .A4(new_n601), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n602), .B2(new_n604), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n634), .A2(new_n636), .B1(new_n485), .B2(new_n455), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n534), .A2(new_n536), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n580), .A2(new_n639), .A3(new_n610), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  INV_X1    g0442(.A(new_n625), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n537), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n644), .A3(new_n624), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n421), .B1(new_n638), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n353), .A2(new_n364), .ZN(new_n647));
  INV_X1    g0447(.A(new_n390), .ZN(new_n648));
  INV_X1    g0448(.A(new_n416), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n394), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n358), .A2(new_n362), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n652), .A2(new_n294), .B1(new_n298), .B2(new_n300), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(KEYINPUT89), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n255), .A2(new_n209), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n455), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n493), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n486), .A2(new_n662), .A3(new_n492), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT89), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n486), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n661), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n661), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n586), .B2(new_n588), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n634), .A2(new_n636), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n605), .A2(new_n607), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n671), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n605), .A2(new_n661), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n663), .A2(new_n665), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n667), .A2(new_n670), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(G399));
  NOR2_X1   g0482(.A1(new_n461), .A2(new_n462), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n213), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n552), .A2(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n206), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  INV_X1    g0488(.A(G330), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n493), .A2(new_n541), .A3(new_n608), .A4(new_n670), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT31), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n469), .A2(new_n475), .A3(new_n568), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT90), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n603), .A2(new_n521), .A3(new_n387), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT92), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n693), .A2(KEYINPUT30), .A3(new_n694), .ZN(new_n699));
  AOI211_X1 g0499(.A(G179), .B(new_n620), .C1(new_n590), .C2(new_n599), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT91), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n539), .A2(new_n701), .A3(new_n484), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n539), .B2(new_n484), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT92), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n695), .A2(new_n705), .A3(new_n696), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n698), .A2(new_n699), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n661), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n691), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n704), .A2(new_n699), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n697), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n689), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n670), .B1(new_n645), .B2(new_n638), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT93), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT93), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n670), .C1(new_n645), .C2(new_n638), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT94), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n537), .A2(new_n720), .A3(KEYINPUT26), .A4(new_n643), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT94), .B1(new_n640), .B2(new_n642), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n615), .A2(new_n642), .A3(new_n625), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n624), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n615), .A2(new_n626), .A3(new_n629), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n486), .A2(new_n605), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n661), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT29), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n713), .B1(new_n719), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n688), .B1(new_n731), .B2(G1), .ZN(G364));
  INV_X1    g0532(.A(new_n684), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n209), .A2(G13), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n255), .B1(new_n734), .B2(G45), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n676), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G330), .B2(new_n674), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT95), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n265), .B(new_n213), .C1(new_n740), .C2(G355), .ZN(new_n741));
  AND2_X1   g0541(.A1(G355), .A2(new_n740), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n741), .A2(new_n742), .B1(G116), .B2(new_n213), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n239), .A2(new_n277), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n309), .A2(new_n213), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n207), .B2(new_n277), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n208), .B1(G20), .B2(new_n296), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n737), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n209), .A2(new_n387), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G322), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n209), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(new_n290), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n758), .A2(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n290), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n209), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(G294), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n755), .A2(new_n290), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT33), .B(G317), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n265), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n755), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n760), .A2(new_n772), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G311), .A2(new_n774), .B1(new_n776), .B2(G329), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n756), .A2(new_n489), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n778), .A2(G326), .B1(new_n780), .B2(G303), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n767), .A2(new_n771), .A3(new_n777), .A4(new_n781), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n265), .B1(new_n761), .B2(new_n219), .C1(new_n312), .C2(new_n779), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT97), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n768), .A2(new_n326), .B1(new_n773), .B2(new_n217), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT32), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT96), .B(G159), .Z(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n775), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n785), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n758), .A2(new_n325), .B1(new_n786), .B2(new_n788), .ZN(new_n790));
  INV_X1    g0590(.A(new_n778), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n791), .A2(new_n202), .B1(new_n504), .B2(new_n765), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n784), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n782), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n754), .B1(new_n795), .B2(new_n751), .ZN(new_n796));
  INV_X1    g0596(.A(new_n750), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n674), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n739), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  NAND3_X1  g0600(.A1(new_n408), .A2(new_n415), .A3(new_n661), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT100), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n408), .A2(new_n415), .A3(KEYINPUT100), .A4(new_n661), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n417), .A2(new_n661), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT99), .Z(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(new_n416), .A3(new_n419), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n748), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n751), .A2(new_n748), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n737), .B1(G77), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n769), .A2(KEYINPUT98), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G283), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n791), .A2(new_n594), .B1(new_n779), .B2(new_n219), .ZN(new_n819));
  INV_X1    g0619(.A(new_n761), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(G87), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n344), .B1(new_n775), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G116), .B2(new_n774), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G97), .A2(new_n766), .B1(new_n757), .B2(G294), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n818), .A2(new_n821), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n787), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G150), .A2(new_n769), .B1(new_n827), .B2(new_n774), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n829), .B2(new_n791), .C1(new_n830), .C2(new_n758), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n309), .B1(new_n776), .B2(G132), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n765), .A2(new_n325), .B1(new_n779), .B2(new_n202), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G68), .B2(new_n820), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n831), .A2(new_n832), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n826), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n813), .B1(new_n839), .B2(new_n751), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n810), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n715), .A2(new_n718), .A3(new_n809), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n805), .A2(new_n808), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n670), .B(new_n843), .C1(new_n645), .C2(new_n638), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n713), .ZN(new_n847));
  INV_X1    g0647(.A(new_n737), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(KEYINPUT101), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n713), .B2(new_n846), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT101), .B1(new_n847), .B2(new_n848), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n841), .B1(new_n850), .B2(new_n851), .ZN(G384));
  AND2_X1   g0652(.A1(new_n498), .A2(new_n499), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT35), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n855), .A2(G116), .A3(new_n210), .A4(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT36), .Z(new_n858));
  OR3_X1    g0658(.A1(new_n327), .A2(new_n206), .A3(new_n217), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n202), .A2(G68), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n255), .B(G13), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n377), .A2(new_n661), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n390), .A2(new_n394), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n377), .A2(new_n661), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n395), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n809), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n690), .A2(KEYINPUT31), .B1(new_n707), .B2(new_n661), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n359), .A2(new_n361), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(new_n659), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n351), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n871), .A2(new_n872), .A3(new_n352), .A4(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n876), .A2(new_n337), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n336), .A2(new_n252), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n350), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n324), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n873), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n871), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n875), .B1(new_n882), .B2(new_n872), .ZN(new_n883));
  INV_X1    g0683(.A(new_n881), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n365), .A2(KEYINPUT103), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT103), .B1(new_n365), .B2(new_n884), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT38), .B(new_n883), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n871), .A2(new_n352), .A3(new_n874), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n875), .ZN(new_n890));
  INV_X1    g0690(.A(new_n365), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n874), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n887), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT40), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n870), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n866), .A2(new_n864), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n843), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n899), .B1(new_n709), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n893), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT104), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n903), .A2(new_n904), .A3(new_n887), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n903), .B2(new_n887), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n709), .A2(new_n900), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n421), .ZN(new_n912));
  OAI21_X1  g0712(.A(G330), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n912), .B2(new_n910), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n719), .A2(new_n421), .A3(new_n730), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(new_n653), .ZN(new_n916));
  INV_X1    g0716(.A(new_n898), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n416), .A2(new_n661), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT102), .Z(new_n919));
  AOI21_X1  g0719(.A(new_n917), .B1(new_n844), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n905), .B2(new_n906), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n895), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n648), .A2(new_n670), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n647), .A2(new_n873), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n916), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n914), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n914), .A2(new_n930), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT105), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n931), .B1(new_n255), .B2(new_n734), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n932), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(KEYINPUT105), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n862), .B1(new_n934), .B2(new_n936), .ZN(G367));
  NOR2_X1   g0737(.A1(new_n627), .A2(new_n670), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n537), .A2(new_n540), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n615), .A2(new_n670), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT107), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n615), .B(new_n629), .C1(new_n627), .C2(new_n670), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n537), .A2(new_n661), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT107), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n679), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT42), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n942), .A2(new_n945), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n615), .B1(new_n951), .B2(new_n486), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n670), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n556), .A2(new_n670), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT106), .Z(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(new_n624), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n643), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n954), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n677), .A2(new_n951), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n950), .A2(new_n961), .A3(new_n960), .A4(new_n953), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n965), .B1(new_n964), .B2(new_n966), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n684), .B(KEYINPUT41), .ZN(new_n970));
  XOR2_X1   g0770(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n971));
  NAND3_X1  g0771(.A1(new_n681), .A2(new_n946), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n971), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n679), .A2(new_n680), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n973), .B1(new_n974), .B2(new_n951), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n974), .A2(new_n951), .A3(KEYINPUT44), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT44), .B1(new_n974), .B2(new_n951), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n972), .B(new_n975), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n677), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n669), .A2(new_n678), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n947), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n676), .A2(KEYINPUT111), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n676), .A2(KEYINPUT111), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n982), .A2(new_n984), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n980), .A2(new_n987), .A3(new_n731), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT109), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n677), .B1(new_n978), .B2(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n972), .A2(new_n975), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n992), .B(KEYINPUT109), .C1(new_n977), .C2(new_n976), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT110), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n994), .B1(new_n991), .B2(new_n993), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n989), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n970), .B1(new_n998), .B2(new_n731), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n969), .B1(new_n999), .B2(new_n736), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n960), .A2(new_n750), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n752), .B1(new_n213), .B2(new_n412), .C1(new_n235), .C2(new_n745), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT112), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n848), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n830), .A2(new_n791), .B1(new_n758), .B2(new_n246), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G58), .B2(new_n780), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n817), .A2(new_n827), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n265), .B1(new_n775), .B2(new_n829), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G50), .B2(new_n774), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n766), .A2(G68), .B1(new_n820), .B2(G77), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n779), .A2(new_n582), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT46), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n758), .A2(new_n594), .B1(new_n761), .B2(new_n504), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n791), .A2(new_n822), .B1(new_n219), .B2(new_n765), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(G317), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n773), .A2(new_n762), .B1(new_n775), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n309), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1017), .B(new_n1021), .C1(new_n473), .C2(new_n816), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1012), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT47), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1005), .B1(new_n1024), .B2(new_n751), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1001), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1000), .A2(new_n1026), .ZN(G387));
  INV_X1    g0827(.A(KEYINPUT113), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n987), .B2(new_n731), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n987), .A2(new_n731), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n731), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(KEYINPUT113), .C1(new_n985), .C2(new_n986), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1029), .A2(new_n733), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n666), .A2(new_n668), .A3(new_n750), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n685), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n213), .A3(new_n265), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(G107), .B2(new_n213), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n232), .A2(new_n277), .ZN(new_n1038));
  AOI211_X1 g0838(.A(G45), .B(new_n1035), .C1(G68), .C2(G77), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n244), .A2(G50), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n745), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1037), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n737), .B1(new_n1043), .B2(new_n753), .ZN(new_n1044));
  INV_X1    g0844(.A(G159), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n791), .A2(new_n1045), .B1(new_n779), .B2(new_n217), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n776), .A2(G150), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n326), .B2(new_n773), .C1(new_n244), .C2(new_n768), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n758), .A2(new_n202), .B1(new_n412), .B2(new_n765), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1020), .B1(new_n504), .B2(new_n761), .ZN(new_n1050));
  OR4_X1    g0850(.A1(new_n1046), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1020), .B1(G326), .B2(new_n776), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n765), .A2(new_n762), .B1(new_n779), .B2(new_n473), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n778), .A2(G322), .B1(new_n774), .B2(G303), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n1018), .B2(new_n758), .C1(new_n816), .C2(new_n822), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT49), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1052), .B1(new_n582), .B2(new_n761), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1051), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1044), .B1(new_n1062), .B2(new_n751), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n987), .A2(new_n736), .B1(new_n1034), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1033), .A2(new_n1064), .ZN(G393));
  XNOR2_X1  g0865(.A(new_n978), .B(new_n979), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n684), .B1(new_n1030), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n998), .A2(new_n1067), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1066), .A2(new_n735), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n752), .B1(new_n504), .B2(new_n213), .C1(new_n242), .C2(new_n745), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n737), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G311), .A2(new_n757), .B1(new_n778), .B2(G317), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT52), .Z(new_n1073));
  OAI22_X1  g0873(.A1(new_n219), .A2(new_n761), .B1(new_n779), .B2(new_n762), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G116), .B2(new_n766), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n344), .B1(new_n775), .B2(new_n759), .C1(new_n473), .C2(new_n773), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n817), .B2(G303), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G150), .A2(new_n778), .B1(new_n757), .B2(G159), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n765), .A2(new_n217), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1020), .B1(new_n244), .B2(new_n773), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(G87), .C2(new_n820), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n779), .A2(new_n326), .B1(new_n775), .B2(new_n830), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT114), .Z(new_n1085));
  OAI211_X1 g0885(.A(new_n1083), .B(new_n1085), .C1(new_n202), .C2(new_n816), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1078), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1071), .B1(new_n1087), .B2(new_n751), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n946), .B2(new_n797), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1068), .A2(new_n1069), .A3(new_n1089), .ZN(G390));
  NAND2_X1  g0890(.A1(new_n724), .A2(new_n728), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n670), .A3(new_n843), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n918), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n917), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n895), .A2(new_n925), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT115), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1095), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT115), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n918), .B1(new_n729), .B2(new_n843), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1097), .B(new_n1098), .C1(new_n1099), .C2(new_n917), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n713), .A2(new_n843), .A3(new_n898), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n844), .A2(new_n919), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n898), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1104), .A2(new_n925), .B1(new_n923), .B2(new_n924), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1101), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n911), .A2(G330), .A3(new_n867), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1105), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n911), .A2(new_n421), .A3(G330), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n915), .A2(new_n653), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1108), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n898), .B1(new_n713), .B2(new_n843), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1103), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n911), .A2(G330), .A3(new_n843), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n917), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n1102), .A3(new_n1099), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1112), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1110), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1107), .B(new_n1119), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n733), .A3(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1107), .B(new_n736), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n816), .A2(new_n219), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n344), .B1(new_n775), .B2(new_n473), .C1(new_n504), .C2(new_n773), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n326), .A2(new_n761), .B1(new_n779), .B2(new_n312), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1081), .B1(G116), .B2(new_n757), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n762), .C2(new_n791), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n344), .B1(new_n776), .B2(G125), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n773), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n817), .B2(G137), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n779), .A2(new_n246), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G159), .A2(new_n766), .B1(new_n757), .B2(G132), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n778), .A2(G128), .B1(new_n820), .B2(G50), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1130), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n751), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n848), .B1(new_n244), .B2(new_n811), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n923), .A2(new_n924), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1141), .B(new_n1142), .C1(new_n1143), .C2(new_n749), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1124), .A2(KEYINPUT116), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT116), .B1(new_n1124), .B2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1123), .B1(new_n1145), .B2(new_n1146), .ZN(G378));
  AND3_X1   g0947(.A1(new_n921), .A2(new_n927), .A3(new_n928), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n901), .A2(KEYINPUT40), .A3(new_n895), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n365), .A2(new_n884), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT103), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n365), .A2(KEYINPUT103), .A3(new_n884), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT38), .B1(new_n1154), .B2(new_n883), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n887), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT104), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n903), .A2(new_n904), .A3(new_n887), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n870), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(G330), .B(new_n1149), .C1(new_n1159), .C2(KEYINPUT40), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1148), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n909), .A2(G330), .A3(new_n929), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n263), .A2(new_n873), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT55), .Z(new_n1164));
  XNOR2_X1  g0964(.A(new_n302), .B(new_n1164), .ZN(new_n1165));
  XOR2_X1   g0965(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1161), .A2(new_n1162), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1167), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1168), .A2(new_n1169), .A3(new_n735), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n773), .A2(new_n829), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n779), .A2(new_n1132), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(G132), .C2(new_n769), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G150), .A2(new_n766), .B1(new_n778), .B2(G125), .ZN(new_n1174));
  INV_X1    g0974(.A(G128), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1174), .C1(new_n1175), .C2(new_n758), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n776), .A2(G124), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n307), .A2(new_n275), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT117), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(new_n761), .C2(new_n787), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1176), .B2(KEYINPUT59), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n309), .A2(new_n683), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1180), .A2(G50), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1177), .A2(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n779), .A2(new_n217), .B1(new_n775), .B2(new_n762), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1183), .B(new_n1186), .C1(G58), .C2(new_n820), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT118), .Z(new_n1188));
  OAI22_X1  g0988(.A1(new_n768), .A2(new_n504), .B1(new_n773), .B2(new_n412), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G68), .B2(new_n766), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G107), .A2(new_n757), .B1(new_n778), .B2(G116), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT58), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1185), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n751), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT119), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n737), .B1(G50), .B2(new_n812), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT120), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(new_n1167), .C2(new_n749), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT122), .ZN(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT123), .B1(new_n1170), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1201), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT123), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1167), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1148), .A2(new_n1160), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n929), .B1(new_n909), .B2(G330), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1161), .A2(new_n1162), .A3(new_n1167), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1203), .B(new_n1204), .C1(new_n1210), .C2(new_n735), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1202), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT57), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1108), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n709), .A2(new_n712), .ZN(new_n1215));
  AND4_X1   g1015(.A1(G330), .A2(new_n1215), .A3(new_n843), .A4(new_n898), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1216), .B(new_n1105), .C1(new_n1096), .C2(new_n1100), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1112), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1213), .B1(new_n1220), .B2(new_n1210), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1112), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1122), .A2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1223), .A2(KEYINPUT57), .A3(new_n1209), .A4(new_n1208), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1221), .A2(new_n733), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1212), .A2(new_n1225), .ZN(G375));
  NAND2_X1  g1026(.A1(new_n917), .A2(new_n748), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n737), .B1(G68), .B2(new_n812), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n817), .A2(G116), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n758), .A2(new_n762), .B1(new_n779), .B2(new_n504), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G294), .B2(new_n778), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n344), .B1(new_n775), .B2(new_n594), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G107), .B2(new_n774), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n766), .A2(new_n542), .B1(new_n820), .B2(G77), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1229), .A2(new_n1231), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n325), .A2(new_n761), .B1(new_n779), .B2(new_n1045), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1020), .B1(new_n1175), .B2(new_n775), .C1(new_n246), .C2(new_n773), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(G50), .C2(new_n766), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT124), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G132), .A2(new_n778), .B1(new_n757), .B2(G137), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n816), .B2(new_n1132), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1235), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1228), .B1(new_n1242), .B2(new_n751), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1219), .A2(new_n736), .B1(new_n1227), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n970), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1120), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1244), .B1(new_n1246), .B2(new_n1247), .ZN(G381));
  OR2_X1    g1048(.A1(G375), .A2(KEYINPUT125), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1033), .A2(new_n799), .A3(new_n1064), .ZN(new_n1250));
  OR3_X1    g1050(.A1(G381), .A2(new_n1250), .A3(G384), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1123), .A2(new_n1124), .A3(new_n1144), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(G387), .A2(new_n1251), .A3(G390), .A4(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G375), .A2(KEYINPUT125), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1249), .A2(new_n1253), .A3(new_n1254), .ZN(G407));
  INV_X1    g1055(.A(new_n1252), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n660), .A2(G213), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1249), .A2(new_n1254), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(G407), .A3(G213), .ZN(G409));
  NAND3_X1  g1060(.A1(new_n1212), .A2(new_n1225), .A3(G378), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1203), .B1(new_n1210), .B2(new_n735), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1220), .A2(new_n1210), .A3(new_n970), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1256), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1257), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1258), .A2(G2897), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1119), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n684), .B1(new_n1270), .B2(new_n1247), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1247), .B2(new_n1270), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(G384), .A3(new_n1244), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G384), .B1(new_n1272), .B2(new_n1244), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1268), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1244), .ZN(new_n1277));
  INV_X1    g1077(.A(G384), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n1273), .A3(new_n1267), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1266), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1283), .B1(new_n1266), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1258), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(KEYINPUT63), .A3(new_n1284), .ZN(new_n1288));
  INV_X1    g1088(.A(G390), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1000), .A2(new_n1026), .A3(G390), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1250), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G390), .B1(new_n1000), .B2(new_n1026), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1292), .A2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1290), .A2(new_n1296), .A3(new_n1291), .A4(new_n1294), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1282), .A2(new_n1286), .A3(new_n1288), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1287), .A2(new_n1302), .A3(new_n1284), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1304), .B1(new_n1287), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1302), .B1(new_n1287), .B2(new_n1284), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1303), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1301), .B1(new_n1308), .B2(new_n1300), .ZN(G405));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1300), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(G375), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1261), .B1(new_n1312), .B2(new_n1252), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1284), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1285), .B(new_n1261), .C1(new_n1312), .C2(new_n1252), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1298), .A2(KEYINPUT127), .A3(new_n1299), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1311), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1300), .A2(new_n1310), .A3(new_n1314), .A4(new_n1315), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(G402));
endmodule


