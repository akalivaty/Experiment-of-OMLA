//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(G472), .A3(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT65), .A2(G137), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT11), .A2(G134), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G137), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G137), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n204), .A2(new_n209), .A3(G131), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT11), .B1(new_n212), .B2(G134), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(G134), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT65), .A2(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n216), .A2(KEYINPUT11), .A3(G134), .A4(new_n200), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n211), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n199), .B1(new_n210), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT2), .B(G113), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G116), .B(G119), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G116), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G119), .ZN(new_n225));
  INV_X1    g039(.A(G119), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G116), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n220), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(G134), .B1(new_n216), .B2(new_n200), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n206), .A2(G137), .ZN(new_n232));
  OAI21_X1  g046(.A(G131), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n215), .A2(new_n217), .A3(new_n211), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n191), .B(new_n193), .C1(KEYINPUT1), .C2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n192), .A2(G146), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n190), .A2(G143), .ZN(new_n239));
  OAI211_X1 g053(.A(G128), .B(new_n237), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n233), .A2(new_n234), .A3(new_n236), .A4(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n219), .A2(new_n230), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(G237), .A2(G953), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G210), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT27), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n195), .B(new_n250), .C1(new_n196), .C2(new_n197), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n249), .B(new_n251), .C1(new_n210), .C2(new_n218), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n241), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT30), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n230), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n219), .A2(KEYINPUT30), .A3(new_n241), .ZN(new_n256));
  AOI211_X1 g070(.A(KEYINPUT31), .B(new_n248), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT31), .ZN(new_n258));
  INV_X1    g072(.A(new_n251), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n260), .B(new_n261), .C1(new_n238), .C2(new_n239), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n250), .B1(new_n262), .B2(new_n195), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(G131), .B1(new_n204), .B2(new_n209), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n234), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n240), .A2(new_n236), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n206), .B1(new_n201), .B2(new_n202), .ZN(new_n268));
  INV_X1    g082(.A(new_n232), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n211), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n264), .A2(new_n266), .B1(new_n234), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n229), .B(new_n256), .C1(new_n272), .C2(KEYINPUT30), .ZN(new_n273));
  INV_X1    g087(.A(new_n248), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n258), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n257), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n253), .A2(new_n229), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n242), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n219), .A2(new_n241), .A3(KEYINPUT28), .A4(new_n230), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n247), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n189), .B1(new_n276), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT30), .B1(new_n252), .B2(new_n241), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n219), .A2(KEYINPUT30), .A3(new_n241), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n285), .A2(new_n286), .A3(new_n230), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT31), .B1(new_n287), .B2(new_n248), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n273), .A2(new_n258), .A3(new_n274), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n189), .A3(new_n289), .A4(new_n283), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n188), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n293));
  INV_X1    g107(.A(new_n242), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n287), .A2(new_n247), .A3(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n281), .A2(new_n247), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n279), .A2(KEYINPUT67), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n230), .B1(new_n219), .B2(new_n241), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n278), .B1(new_n300), .B2(new_n242), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n279), .A2(KEYINPUT67), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n282), .A2(new_n293), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G472), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n292), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n288), .A2(new_n283), .A3(new_n289), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT66), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n290), .ZN(new_n311));
  NOR2_X1   g125(.A1(G472), .A2(G902), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT32), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT68), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n284), .B2(new_n291), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n187), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n311), .A2(new_n188), .B1(G472), .B2(new_n306), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G125), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G140), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT16), .ZN(new_n324));
  OR3_X1    g138(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G146), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G125), .B(G140), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n190), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT70), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n226), .A2(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n235), .A2(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n335), .A2(G110), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(G110), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n330), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n333), .A2(KEYINPUT70), .A3(new_n336), .A4(new_n337), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n235), .A2(KEYINPUT23), .A3(G119), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n226), .A2(G128), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n331), .B(new_n341), .C1(new_n342), .C2(KEYINPUT23), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n339), .B(new_n340), .C1(G110), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n329), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n343), .A2(G110), .B1(new_n334), .B2(new_n338), .ZN(new_n346));
  AOI21_X1  g160(.A(G146), .B1(new_n324), .B2(new_n325), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n346), .B(KEYINPUT69), .C1(new_n347), .C2(new_n327), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n347), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n326), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT69), .B1(new_n351), .B2(new_n346), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n345), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G953), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(G221), .A3(G234), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT71), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G137), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n358), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT72), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT72), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n345), .B(new_n362), .C1(new_n349), .C2(new_n352), .ZN(new_n366));
  INV_X1    g180(.A(G217), .ZN(new_n367));
  INV_X1    g181(.A(G902), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(G234), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT74), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n365), .A2(new_n366), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n373), .A2(new_n374), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n377), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n365), .A2(new_n379), .A3(new_n366), .A4(new_n375), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n380), .A3(new_n369), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n372), .A2(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n314), .A2(new_n319), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n384));
  OAI21_X1  g198(.A(G214), .B1(G237), .B2(G902), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G210), .B1(G237), .B2(G902), .ZN(new_n387));
  INV_X1    g201(.A(new_n267), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n322), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n199), .A2(G125), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n354), .A2(G224), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(KEYINPUT7), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(KEYINPUT7), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT80), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G104), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT3), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G107), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n399), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G101), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT75), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(KEYINPUT75), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(G104), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n404), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n403), .B2(new_n399), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n222), .A2(KEYINPUT5), .ZN(new_n414));
  INV_X1    g228(.A(G113), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n225), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n223), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n411), .A2(new_n418), .A3(new_n223), .A4(new_n412), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G110), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT8), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT80), .A4(new_n394), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n393), .A2(new_n397), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n400), .A2(KEYINPUT3), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n401), .B1(new_n403), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n402), .A2(G107), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n407), .B2(new_n409), .ZN(new_n431));
  OAI21_X1  g245(.A(G101), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n432), .A2(KEYINPUT4), .A3(new_n411), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n434), .B(G101), .C1(new_n429), .C2(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n229), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n423), .B(new_n421), .C1(new_n433), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n368), .B1(new_n427), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n421), .B1(new_n433), .B2(new_n436), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n442));
  INV_X1    g256(.A(new_n423), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n437), .A2(KEYINPUT6), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n432), .A2(KEYINPUT4), .A3(new_n411), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n229), .A3(new_n435), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n423), .B1(new_n447), .B2(new_n421), .ZN(new_n448));
  OAI211_X1 g262(.A(KEYINPUT79), .B(new_n444), .C1(new_n445), .C2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n448), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT79), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT6), .A4(new_n437), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n391), .B(new_n392), .Z(new_n454));
  OAI211_X1 g268(.A(new_n387), .B(new_n440), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n387), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n449), .B2(new_n452), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n439), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n386), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G113), .B(G122), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(G104), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G237), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n354), .A3(G214), .ZN(new_n464));
  NOR2_X1   g278(.A1(KEYINPUT82), .A2(G143), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n243), .B(G214), .C1(KEYINPUT82), .C2(G143), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT18), .A3(G131), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n328), .B(new_n190), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT18), .A2(G131), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n327), .A2(new_n347), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n466), .A2(new_n467), .A3(new_n211), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n211), .B1(new_n466), .B2(new_n467), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT17), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n474), .B1(new_n477), .B2(KEYINPUT85), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n468), .A2(G131), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n466), .A2(new_n467), .A3(new_n211), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n479), .A2(KEYINPUT85), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n476), .A2(new_n483), .A3(KEYINPUT17), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n476), .B2(KEYINPUT17), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n462), .B(new_n473), .C1(new_n478), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n468), .A2(KEYINPUT17), .A3(G131), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT84), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n476), .A2(new_n483), .A3(KEYINPUT17), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n491), .A2(new_n495), .A3(new_n474), .A4(new_n482), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n462), .B1(new_n496), .B2(new_n473), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n368), .B1(new_n488), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G475), .ZN(new_n499));
  NAND2_X1  g313(.A1(G234), .A2(G237), .ZN(new_n500));
  INV_X1    g314(.A(G952), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n501), .A2(KEYINPUT90), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(KEYINPUT90), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n354), .B(new_n500), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n500), .A2(G902), .A3(G953), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT21), .B(G898), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT19), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT19), .B1(new_n321), .B2(new_n323), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n190), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n512), .B(new_n326), .C1(new_n475), .C2(new_n476), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n473), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n461), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT83), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT83), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n517), .A3(new_n461), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n487), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n519), .B2(new_n521), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n499), .B(new_n509), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT9), .B(G234), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n526), .A2(new_n367), .A3(G953), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n235), .B2(G143), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n235), .A2(G143), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT87), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n192), .A2(G128), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n192), .A2(G128), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n533), .B(new_n534), .C1(new_n535), .C2(new_n529), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(KEYINPUT13), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n538), .A2(new_n539), .A3(G134), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n538), .B2(G134), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n235), .A2(G143), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n534), .A2(new_n542), .A3(new_n206), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n224), .A2(G122), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT86), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n224), .A3(G122), .ZN(new_n546));
  INV_X1    g360(.A(G122), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT86), .B1(new_n547), .B2(G116), .ZN(new_n548));
  AOI211_X1 g362(.A(G107), .B(new_n544), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n546), .ZN(new_n550));
  INV_X1    g364(.A(new_n544), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n398), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n543), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n540), .A2(new_n541), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G134), .B1(new_n531), .B2(new_n535), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n543), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n398), .A3(new_n551), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n544), .B1(new_n550), .B2(KEYINPUT14), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(KEYINPUT14), .B2(new_n550), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n560), .B2(G107), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n528), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n538), .A2(G134), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT88), .ZN(new_n564));
  INV_X1    g378(.A(new_n543), .ZN(new_n565));
  INV_X1    g379(.A(new_n552), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(new_n557), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n538), .A2(new_n539), .A3(G134), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n561), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT89), .A4(new_n527), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n541), .A2(new_n553), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n561), .B1(new_n573), .B2(new_n568), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT89), .B1(new_n574), .B2(new_n527), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n368), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G478), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(KEYINPUT15), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n570), .A3(new_n527), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n562), .A3(new_n571), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n583), .B(new_n368), .C1(KEYINPUT15), .C2(new_n577), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n525), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n459), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G221), .B1(new_n526), .B2(G902), .ZN(new_n588));
  XNOR2_X1  g402(.A(G110), .B(G140), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n354), .A2(G227), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n446), .A2(new_n199), .A3(new_n435), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n413), .B2(new_n267), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n388), .A2(KEYINPUT10), .A3(new_n411), .A4(new_n412), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n266), .ZN(new_n598));
  INV_X1    g412(.A(new_n266), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n593), .A2(new_n595), .A3(new_n599), .A4(new_n596), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n592), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n592), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n413), .A2(new_n267), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n411), .A2(new_n412), .B1(new_n236), .B2(new_n240), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n266), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT76), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT12), .B1(new_n266), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n607), .B(new_n266), .C1(new_n603), .C2(new_n604), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n601), .A2(KEYINPUT78), .B1(new_n602), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n600), .A2(new_n592), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT78), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n609), .A4(new_n610), .ZN(new_n615));
  AOI211_X1 g429(.A(G469), .B(G902), .C1(new_n612), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n602), .A2(KEYINPUT77), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT77), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n600), .A2(new_n618), .A3(new_n592), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n598), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n609), .A2(new_n610), .A3(new_n600), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n591), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(G469), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(G469), .A2(G902), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n588), .B1(new_n616), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n384), .B1(new_n587), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n588), .ZN(new_n628));
  INV_X1    g442(.A(new_n625), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n612), .A2(new_n615), .ZN(new_n630));
  INV_X1    g444(.A(G469), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n368), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n628), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n633), .A2(KEYINPUT91), .A3(new_n459), .A4(new_n586), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n383), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT92), .B(G101), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G3));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n572), .B2(new_n575), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT93), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n569), .A2(new_n570), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n639), .B1(new_n642), .B2(new_n528), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n580), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n577), .A2(G902), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n640), .A2(new_n641), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n576), .A2(new_n577), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n583), .A2(new_n639), .B1(new_n580), .B2(new_n643), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n641), .B1(new_n649), .B2(new_n645), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n499), .B1(new_n522), .B2(new_n524), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n653), .A2(new_n459), .A3(new_n509), .ZN(new_n654));
  AOI21_X1  g468(.A(G902), .B1(new_n310), .B2(new_n290), .ZN(new_n655));
  INV_X1    g469(.A(G472), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n315), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n382), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n657), .A2(new_n658), .A3(new_n626), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT94), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  AND3_X1   g477(.A1(new_n519), .A2(new_n523), .A3(new_n521), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n524), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(G475), .B2(new_n498), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n508), .B(KEYINPUT95), .Z(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n459), .A2(new_n666), .A3(new_n585), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n659), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  INV_X1    g486(.A(KEYINPUT96), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n364), .A2(new_n361), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT36), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  AOI211_X1 g491(.A(KEYINPUT96), .B(KEYINPUT36), .C1(new_n364), .C2(new_n361), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n353), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n353), .B1(new_n676), .B2(new_n678), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n370), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n381), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT97), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n381), .A2(KEYINPUT97), .A3(new_n683), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n657), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n627), .A2(new_n689), .A3(new_n634), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT37), .B(G110), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  INV_X1    g506(.A(new_n688), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n314), .A2(new_n319), .A3(new_n633), .A4(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(G900), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n505), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n504), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n666), .A2(new_n585), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT98), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT98), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n666), .A2(new_n700), .A3(new_n585), .A4(new_n697), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n459), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  XNOR2_X1  g518(.A(new_n697), .B(KEYINPUT39), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n626), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n282), .B1(new_n273), .B2(new_n242), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n294), .A2(new_n299), .A3(new_n247), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT100), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n368), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n710), .A2(KEYINPUT100), .A3(new_n711), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n316), .A2(new_n715), .A3(new_n292), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n381), .A3(new_n683), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n455), .A2(new_n458), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(new_n385), .A3(new_n585), .A4(new_n652), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n709), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(KEYINPUT40), .B2(new_n708), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G143), .ZN(G45));
  INV_X1    g538(.A(KEYINPUT101), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n652), .B(new_n697), .C1(new_n648), .C2(new_n650), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n725), .B1(new_n727), .B2(new_n459), .ZN(new_n728));
  INV_X1    g542(.A(new_n459), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n726), .A2(new_n729), .A3(KEYINPUT101), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n694), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n190), .ZN(G48));
  NAND3_X1  g546(.A1(new_n314), .A2(new_n319), .A3(new_n382), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n631), .B1(new_n630), .B2(new_n368), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n616), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT102), .B1(new_n735), .B2(new_n588), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(KEYINPUT102), .A3(new_n588), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n733), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n654), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n669), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  NAND2_X1  g558(.A1(new_n314), .A2(new_n319), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n688), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n738), .A2(new_n736), .A3(new_n729), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n586), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  OAI21_X1  g563(.A(new_n276), .B1(new_n247), .B2(new_n303), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n312), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n382), .B(new_n751), .C1(new_n655), .C2(new_n656), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n630), .A2(new_n368), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(G469), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n588), .A3(new_n632), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT102), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n718), .A2(new_n385), .A3(new_n668), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n585), .A2(new_n652), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n753), .A2(new_n758), .A3(new_n761), .A4(new_n737), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  OAI211_X1 g577(.A(new_n684), .B(new_n751), .C1(new_n655), .C2(new_n656), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n726), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n459), .A3(new_n758), .A4(new_n737), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n622), .A2(KEYINPUT103), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT103), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n621), .A2(new_n770), .A3(new_n591), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(G469), .A3(new_n620), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n624), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n588), .B1(new_n616), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n455), .A2(new_n385), .A3(new_n458), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n314), .A2(new_n319), .A3(new_n776), .A4(new_n382), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n768), .B1(new_n777), .B2(new_n726), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n658), .B1(new_n316), .B2(new_n317), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(KEYINPUT42), .A3(new_n776), .A4(new_n727), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  AND4_X1   g596(.A1(new_n314), .A2(new_n319), .A3(new_n382), .A4(new_n776), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n699), .A2(new_n701), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(KEYINPUT104), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT104), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(new_n777), .B2(new_n784), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G134), .ZN(G36));
  NAND4_X1  g604(.A1(new_n769), .A2(KEYINPUT45), .A3(new_n620), .A4(new_n771), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n620), .A2(new_n622), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n791), .B(G469), .C1(new_n792), .C2(KEYINPUT45), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n624), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n616), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n588), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n706), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n652), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n651), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT43), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n657), .A3(new_n684), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n775), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n805), .B2(new_n806), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n800), .B(new_n807), .C1(KEYINPUT105), .C2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(KEYINPUT105), .B2(new_n809), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  NOR2_X1   g626(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n813));
  AND2_X1   g627(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n798), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n798), .B2(new_n814), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n745), .A2(new_n658), .A3(new_n727), .A4(new_n808), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n320), .ZN(G42));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n314), .A2(new_n319), .A3(new_n633), .A4(new_n693), .ZN(new_n821));
  INV_X1    g635(.A(new_n585), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n808), .A2(new_n822), .A3(new_n666), .A4(new_n697), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n821), .A2(new_n824), .B1(new_n765), .B2(new_n776), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT104), .B1(new_n783), .B2(new_n785), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n777), .A2(new_n787), .A3(new_n784), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT109), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n738), .A2(new_n736), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n383), .B(new_n831), .C1(new_n654), .C2(new_n669), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n748), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT108), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n801), .A2(new_n585), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n759), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n651), .A2(new_n459), .A3(new_n652), .A4(new_n668), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n822), .A2(new_n652), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n459), .A3(KEYINPUT108), .A4(new_n668), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n659), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n636), .A2(new_n690), .A3(new_n762), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n833), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n789), .A2(KEYINPUT109), .A3(new_n825), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n830), .A2(new_n843), .A3(new_n781), .A4(new_n844), .ZN(new_n845));
  OR3_X1    g659(.A1(new_n694), .A2(new_n728), .A3(new_n730), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n729), .A2(new_n760), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n632), .A2(new_n624), .A3(new_n772), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n588), .A3(new_n697), .A4(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n717), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n846), .A2(new_n703), .A3(new_n766), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT52), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n766), .B1(new_n694), .B2(new_n702), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n731), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n851), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  OR3_X1    g673(.A1(new_n845), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n765), .A2(new_n776), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(new_n694), .B2(new_n823), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n829), .B(new_n862), .C1(new_n788), .C2(new_n786), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n627), .A2(new_n634), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n690), .B(new_n762), .C1(new_n733), .C2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n840), .A2(new_n659), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n748), .A3(new_n781), .A4(new_n832), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g683(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n855), .B2(new_n851), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n731), .A2(new_n854), .A3(new_n850), .A4(KEYINPUT52), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n869), .A2(new_n873), .A3(new_n830), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n859), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n820), .B1(new_n860), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n859), .B1(new_n845), .B2(new_n858), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n869), .A2(new_n873), .A3(KEYINPUT53), .A4(new_n830), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n820), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT111), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n831), .A2(new_n808), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT114), .Z(new_n885));
  NOR2_X1   g699(.A1(new_n716), .A2(new_n658), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n885), .A2(new_n504), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n651), .A2(new_n652), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT115), .Z(new_n891));
  NOR2_X1   g705(.A1(new_n720), .A2(new_n385), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n831), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT113), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n752), .A2(new_n504), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n803), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT50), .ZN(new_n898));
  INV_X1    g712(.A(new_n764), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n885), .A2(new_n504), .A3(new_n803), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n735), .B(KEYINPUT107), .Z(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n816), .B1(new_n588), .B2(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n803), .A2(new_n775), .A3(new_n895), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n891), .A2(KEYINPUT51), .A3(new_n901), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n888), .A2(new_n653), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n354), .B1(new_n502), .B2(new_n503), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n896), .B2(new_n747), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n900), .A2(new_n779), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT48), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(KEYINPUT116), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n911), .B(new_n914), .C1(new_n912), .C2(new_n915), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n906), .B(KEYINPUT112), .Z(new_n917));
  AND3_X1   g731(.A1(new_n891), .A2(new_n901), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n907), .B(new_n916), .C1(new_n918), .C2(KEYINPUT51), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n883), .A2(new_n919), .B1(G952), .B2(G953), .ZN(new_n920));
  NOR4_X1   g734(.A1(new_n887), .A2(new_n628), .A3(new_n386), .A4(new_n720), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n801), .A3(new_n651), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n902), .B(KEYINPUT49), .Z(new_n923));
  OAI21_X1  g737(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G75));
  NAND2_X1  g738(.A1(new_n501), .A2(G953), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n877), .A2(new_n878), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT119), .B1(new_n926), .B2(G902), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n928), .B(new_n368), .C1(new_n877), .C2(new_n878), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n927), .A2(new_n929), .A3(new_n387), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n453), .B(new_n454), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT56), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n925), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n926), .A2(G210), .A3(G902), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(KEYINPUT117), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n935), .B2(KEYINPUT117), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n932), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT118), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n934), .B1(new_n941), .B2(new_n942), .ZN(G51));
  XOR2_X1   g757(.A(new_n624), .B(KEYINPUT57), .Z(new_n944));
  AOI21_X1  g758(.A(new_n820), .B1(new_n877), .B2(new_n878), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n880), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n630), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n927), .A2(new_n929), .A3(new_n793), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR4_X1   g764(.A1(new_n927), .A2(new_n929), .A3(KEYINPUT120), .A4(new_n793), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n925), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT121), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT121), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n954), .B(new_n925), .C1(new_n950), .C2(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G54));
  NOR2_X1   g770(.A1(new_n927), .A2(new_n929), .ZN(new_n957));
  NAND2_X1  g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT122), .Z(new_n959));
  AND2_X1   g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(new_n519), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n519), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n961), .A2(new_n925), .A3(new_n962), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT59), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n649), .B1(new_n883), .B2(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n649), .B(new_n966), .C1(new_n880), .C2(new_n945), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n925), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n877), .B2(new_n878), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n681), .A3(new_n682), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n365), .A2(new_n366), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT123), .Z(new_n976));
  OAI211_X1 g790(.A(new_n974), .B(new_n925), .C1(new_n973), .C2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT61), .B1(new_n974), .B2(KEYINPUT124), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G66));
  INV_X1    g793(.A(G224), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n506), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n843), .A2(G953), .ZN(new_n983));
  MUX2_X1   g797(.A(new_n982), .B(KEYINPUT125), .S(new_n983), .Z(new_n984));
  OAI21_X1  g798(.A(new_n453), .B1(G898), .B2(new_n354), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(G69));
  INV_X1    g800(.A(new_n818), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n723), .A2(new_n855), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT62), .Z(new_n989));
  NOR3_X1   g803(.A1(new_n733), .A2(new_n708), .A3(new_n775), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n653), .B2(new_n838), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n811), .A2(new_n987), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n285), .A2(new_n286), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT126), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n510), .A2(new_n511), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n992), .A2(new_n354), .A3(new_n997), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n987), .A2(new_n781), .A3(new_n789), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n799), .A2(new_n779), .A3(new_n847), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT127), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n811), .A2(new_n855), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  MUX2_X1   g816(.A(new_n695), .B(new_n1002), .S(new_n354), .Z(new_n1003));
  OAI21_X1  g817(.A(new_n998), .B1(new_n1003), .B2(new_n997), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n354), .B1(G227), .B2(G900), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1004), .B(new_n1005), .Z(G72));
  INV_X1    g820(.A(new_n295), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g824(.A(new_n710), .B(new_n1010), .C1(new_n860), .C2(new_n875), .ZN(new_n1011));
  INV_X1    g825(.A(new_n843), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1009), .B1(new_n1002), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n295), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n925), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1009), .B1(new_n992), .B2(new_n1012), .ZN(new_n1016));
  AOI211_X1 g830(.A(new_n1011), .B(new_n1015), .C1(new_n710), .C2(new_n1016), .ZN(G57));
endmodule


