//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n542, new_n543,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(new_n453), .B2(G567), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  NAND3_X1  g032(.A1(new_n457), .A2(G101), .A3(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g035(.A1(new_n457), .A2(KEYINPUT68), .A3(G101), .A4(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n457), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n457), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n457), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(G100), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n480), .A2(new_n457), .A3(KEYINPUT70), .ZN(new_n481));
  AOI21_X1  g056(.A(KEYINPUT70), .B1(new_n480), .B2(new_n457), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G112), .B2(new_n457), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n477), .A2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(G136), .B2(new_n485), .ZN(G162));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  AND2_X1   g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n463), .B2(new_n464), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n463), .B2(new_n464), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n464), .C2(new_n463), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(new_n505), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n506), .A2(new_n516), .ZN(G166));
  AOI22_X1  g092(.A1(new_n513), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n501), .A2(new_n502), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(new_n511), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n520), .A2(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n505), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n511), .A2(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n514), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G171));
  AOI22_X1  g107(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n505), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n501), .A2(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G81), .B1(new_n511), .B2(G43), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  NAND4_X1  g114(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT71), .Z(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(G188));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n545));
  NAND2_X1  g120(.A1(G53), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n513), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n535), .A2(G91), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n546), .B1(new_n509), .B2(new_n510), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT72), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT72), .B1(new_n553), .B2(new_n545), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n551), .B(new_n552), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n519), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n561), .A2(KEYINPUT74), .A3(G651), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n564), .B2(new_n505), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n558), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n535), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n511), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(new_n511), .A2(G48), .ZN(new_n575));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n514), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n503), .A2(G61), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n505), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  AND2_X1   g157(.A1(new_n503), .A2(G60), .ZN(new_n583));
  AND2_X1   g158(.A1(G72), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT76), .B(G85), .Z(new_n588));
  AOI22_X1  g163(.A1(new_n535), .A2(new_n588), .B1(new_n511), .B2(G47), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n585), .A2(new_n586), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NOR2_X1   g168(.A1(G301), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n519), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G54), .B2(new_n511), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n514), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n535), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n594), .B1(new_n606), .B2(new_n593), .ZN(G284));
  AOI21_X1  g182(.A(new_n594), .B1(new_n606), .B2(new_n593), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n562), .A2(new_n565), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n557), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n609), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G559), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(G860), .B2(new_n606), .ZN(G148));
  NAND2_X1  g191(.A1(new_n537), .A2(new_n593), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n615), .B2(new_n593), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI21_X1  g194(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G2104), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n485), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n478), .A2(G123), .ZN(new_n627));
  OR2_X1    g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n628), .B(G2104), .C1(G111), .C2(new_n457), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(G2096), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n625), .A2(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n637), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n647), .A3(G14), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT80), .Z(new_n651));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT17), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT81), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(new_n652), .ZN(new_n657));
  INV_X1    g232(.A(new_n654), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n657), .B(new_n658), .C1(new_n653), .C2(new_n651), .ZN(new_n659));
  INV_X1    g234(.A(new_n652), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n650), .A3(new_n654), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n656), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n669), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(KEYINPUT82), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT83), .ZN(new_n680));
  XOR2_X1   g255(.A(G1981), .B(G1986), .Z(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n680), .B(new_n685), .ZN(G229));
  NOR2_X1   g261(.A1(G6), .A2(G16), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n581), .B2(G16), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G23), .ZN(new_n692));
  INV_X1    g267(.A(G288), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT33), .B(G1976), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(G22), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n691), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1971), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n690), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT34), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n691), .A2(G24), .ZN(new_n703));
  INV_X1    g278(.A(G290), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n691), .ZN(new_n705));
  INV_X1    g280(.A(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(new_n701), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G25), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n485), .A2(G131), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n478), .A2(G119), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n457), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n710), .B1(new_n716), .B2(new_n709), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT35), .B(G1991), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT84), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n717), .B(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n702), .A2(new_n707), .A3(new_n708), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT36), .ZN(new_n722));
  NOR2_X1   g297(.A1(G16), .A2(G19), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n538), .B2(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(G164), .A2(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G27), .B2(G29), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT91), .B(G2078), .Z(new_n727));
  AOI22_X1  g302(.A1(new_n724), .A2(G1341), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G168), .A2(new_n691), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n691), .B2(G21), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT88), .B(G1966), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n728), .B1(new_n730), .B2(new_n731), .C1(new_n726), .C2(new_n727), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n724), .A2(G1341), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n731), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT31), .B(G11), .Z(new_n735));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n709), .B1(new_n736), .B2(G28), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT89), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n738), .A2(KEYINPUT89), .B1(new_n736), .B2(G28), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n735), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n630), .A2(new_n709), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n733), .A2(new_n734), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n732), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n485), .A2(G141), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n478), .A2(G129), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT26), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n457), .A2(G2104), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n749), .A2(new_n750), .B1(G105), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n745), .A2(new_n746), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(new_n709), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n709), .B2(G32), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n691), .A2(G5), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G171), .B2(new_n691), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT90), .ZN(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n756), .A2(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n709), .A2(G26), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n457), .A2(G116), .ZN(new_n766));
  OAI21_X1  g341(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n478), .A2(G128), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n485), .A2(G140), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n709), .B1(new_n774), .B2(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n774), .B2(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G160), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n709), .A2(G33), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n781));
  NAND3_X1  g356(.A1(new_n457), .A2(G103), .A3(G2104), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n457), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G139), .B2(new_n485), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n780), .B1(new_n786), .B2(new_n709), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n779), .B1(new_n787), .B2(G2072), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G2072), .B2(new_n787), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n744), .A2(new_n762), .A3(new_n773), .A4(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n756), .A2(new_n757), .ZN(new_n791));
  NAND2_X1  g366(.A1(G162), .A2(G29), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G29), .B2(G35), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT29), .B(G2090), .Z(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n760), .A2(new_n761), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n791), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n691), .A2(G20), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT23), .Z(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G299), .B2(G16), .ZN(new_n801));
  INV_X1    g376(.A(G1956), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G4), .A2(G16), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n606), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT85), .B(G1348), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n790), .A2(new_n798), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n722), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT92), .Z(G311));
  XOR2_X1   g385(.A(new_n809), .B(KEYINPUT93), .Z(G150));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n505), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n511), .A2(G55), .ZN(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n514), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n812), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n535), .A2(G93), .B1(new_n511), .B2(G55), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n819), .B(KEYINPUT94), .C1(new_n505), .C2(new_n813), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n606), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n818), .A2(new_n537), .A3(new_n820), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n534), .B(new_n536), .C1(new_n814), .C2(new_n817), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT95), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n826), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n825), .B(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n834));
  INV_X1    g409(.A(G860), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n833), .B2(KEYINPUT39), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n823), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT96), .Z(G145));
  XNOR2_X1  g413(.A(G162), .B(new_n630), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G160), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(G118), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(G2105), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n478), .B2(G130), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n485), .A2(KEYINPUT97), .A3(G142), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT97), .B1(new_n485), .B2(G142), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT98), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n622), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n849), .A2(new_n622), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n851), .A2(new_n715), .A3(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n848), .B(KEYINPUT98), .Z(new_n854));
  INV_X1    g429(.A(new_n622), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n716), .B1(new_n856), .B2(new_n850), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n841), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n471), .A2(new_n491), .B1(new_n860), .B2(new_n489), .ZN(new_n861));
  INV_X1    g436(.A(new_n499), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n498), .B1(new_n471), .B2(new_n495), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n771), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n769), .A2(G164), .A3(new_n770), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(new_n754), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n754), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n869), .A2(new_n786), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n786), .B1(new_n869), .B2(new_n870), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n715), .B1(new_n851), .B2(new_n852), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n856), .A2(new_n716), .A3(new_n850), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(KEYINPUT99), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n858), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n873), .B1(new_n858), .B2(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n840), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n853), .A2(new_n857), .A3(new_n841), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT99), .B1(new_n874), .B2(new_n875), .ZN(new_n881));
  OAI22_X1  g456(.A1(new_n880), .A2(new_n881), .B1(new_n871), .B2(new_n872), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n853), .A2(new_n857), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n840), .B1(new_n883), .B2(new_n873), .ZN(new_n884));
  AOI21_X1  g459(.A(G37), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n879), .A2(new_n885), .A3(KEYINPUT40), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT40), .B1(new_n879), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(G395));
  NOR2_X1   g463(.A1(new_n821), .A2(G868), .ZN(new_n889));
  XNOR2_X1  g464(.A(G290), .B(G305), .ZN(new_n890));
  XNOR2_X1  g465(.A(G166), .B(G288), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT42), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n893), .A2(KEYINPUT102), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n615), .B(new_n832), .ZN(new_n895));
  INV_X1    g470(.A(new_n604), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT100), .B1(G299), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n611), .A2(new_n604), .ZN(new_n898));
  NAND2_X1  g473(.A1(G299), .A2(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n897), .B1(new_n900), .B2(KEYINPUT100), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n901), .A2(new_n904), .B1(new_n905), .B2(new_n900), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n903), .B1(new_n906), .B2(new_n895), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n894), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n893), .B2(KEYINPUT102), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n894), .B2(new_n907), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n889), .B1(new_n908), .B2(new_n910), .ZN(G295));
  AOI21_X1  g486(.A(new_n889), .B1(new_n908), .B2(new_n910), .ZN(G331));
  AND3_X1   g487(.A1(new_n826), .A2(new_n830), .A3(new_n827), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n830), .B1(new_n826), .B2(new_n827), .ZN(new_n914));
  OAI21_X1  g489(.A(G171), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n829), .A2(G301), .A3(new_n831), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(G286), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n916), .A3(G168), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n900), .A2(new_n905), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT103), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n901), .B1(new_n920), .B2(new_n904), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n892), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n915), .A2(new_n916), .A3(G168), .ZN(new_n926));
  AOI21_X1  g501(.A(G168), .B1(new_n915), .B2(new_n916), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n906), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n918), .A2(new_n901), .A3(new_n919), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n892), .ZN(new_n931));
  AOI21_X1  g506(.A(G37), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n925), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n925), .A2(new_n932), .A3(KEYINPUT105), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(KEYINPUT43), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n931), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n928), .A2(new_n929), .A3(new_n892), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n925), .A2(new_n932), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT104), .B1(new_n949), .B2(new_n943), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n951));
  AOI211_X1 g526(.A(new_n951), .B(KEYINPUT44), .C1(new_n946), .C2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n945), .B1(new_n950), .B2(new_n952), .ZN(G397));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT45), .B1(new_n864), .B2(new_n954), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n620), .A2(G137), .B1(new_n460), .B2(new_n461), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n467), .A2(new_n468), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n956), .B(G40), .C1(new_n957), .C2(new_n457), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n955), .A2(KEYINPUT114), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(G164), .B2(G1384), .ZN(new_n962));
  INV_X1    g537(.A(G40), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n466), .A2(new_n469), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n960), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n959), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT122), .ZN(new_n967));
  INV_X1    g542(.A(G2078), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n969));
  NAND3_X1  g544(.A1(new_n864), .A2(new_n954), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n497), .A2(new_n499), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n973), .B2(new_n861), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT115), .A3(new_n969), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT114), .B1(new_n955), .B2(new_n958), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n962), .A2(new_n960), .A3(new_n964), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n976), .A2(new_n978), .A3(new_n968), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT122), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n981), .A3(KEYINPUT53), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n864), .A2(new_n954), .ZN(new_n983));
  INV_X1    g558(.A(new_n969), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n958), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n968), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n864), .A2(new_n990), .A3(new_n954), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n964), .A3(new_n991), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n987), .A2(new_n988), .B1(new_n761), .B2(new_n992), .ZN(new_n993));
  AOI211_X1 g568(.A(KEYINPUT123), .B(G301), .C1(new_n982), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT123), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n980), .A2(KEYINPUT122), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT53), .B1(new_n980), .B2(KEYINPUT122), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n998), .B2(G171), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n993), .B1(new_n988), .B2(new_n987), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(G171), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n994), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT124), .B1(new_n1002), .B2(KEYINPUT54), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT124), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n998), .A2(G171), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT123), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n998), .A2(new_n995), .A3(G171), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1004), .B(new_n1005), .C1(new_n1009), .C2(new_n1001), .ZN(new_n1010));
  INV_X1    g585(.A(G2067), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n983), .A2(new_n958), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT118), .B1(new_n974), .B2(new_n964), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1348), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n992), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(KEYINPUT60), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n614), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1015), .A2(new_n606), .A3(KEYINPUT60), .A4(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT60), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1017), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1012), .B1(new_n983), .B2(new_n958), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n974), .A2(new_n964), .A3(KEYINPUT118), .ZN(new_n1024));
  AOI21_X1  g599(.A(G2067), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1019), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT58), .B(G1341), .Z(new_n1028));
  NAND3_X1  g603(.A1(new_n1023), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n984), .B1(G164), .B2(G1384), .ZN(new_n1030));
  INV_X1    g605(.A(G1996), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n986), .A2(new_n1030), .A3(new_n1031), .A4(new_n964), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT59), .B1(new_n1033), .B2(new_n538), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1035), .B(new_n537), .C1(new_n1029), .C2(new_n1032), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n992), .A2(new_n802), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT56), .B(G2072), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n985), .A2(new_n986), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1041), .A2(KEYINPUT117), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(KEYINPUT117), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1042), .B(new_n1043), .C1(new_n610), .C2(new_n557), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n558), .A2(KEYINPUT117), .A3(new_n566), .A4(new_n1041), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1038), .A2(new_n1040), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT61), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT120), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT61), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1038), .A2(new_n1040), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1046), .B(new_n1048), .C1(new_n1054), .C2(KEYINPUT61), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1027), .A2(new_n1037), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1050), .A2(KEYINPUT119), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1038), .A2(new_n1040), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n1051), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n606), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1046), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1056), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n974), .A2(new_n964), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT110), .B(G8), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1066), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT49), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n577), .A2(new_n580), .A3(G1981), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1981), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n578), .A2(new_n579), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G651), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n535), .A2(G86), .B1(new_n511), .B2(G48), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1072), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1073), .A2(new_n1079), .A3(KEYINPUT49), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1070), .A2(new_n1071), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n693), .A2(G1976), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT52), .B1(G288), .B2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1084), .B(new_n1086), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1071), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1069), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1089), .B1(new_n1091), .B2(new_n1084), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G303), .A2(G8), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1971), .B1(new_n985), .B2(new_n986), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT108), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1098), .A2(new_n1099), .B1(G2090), .B2(new_n992), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1097), .B(G8), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n992), .A2(KEYINPUT113), .ZN(new_n1103));
  AOI21_X1  g678(.A(G2090), .B1(new_n992), .B2(KEYINPUT113), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1098), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1096), .B1(new_n1105), .B2(new_n1067), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1093), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1005), .B1(new_n1000), .B2(G171), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n998), .B2(G171), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1064), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n992), .A2(G2084), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n976), .A2(new_n979), .A3(new_n978), .ZN(new_n1112));
  INV_X1    g687(.A(G1966), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G168), .A2(new_n1067), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1966), .B1(new_n966), .B2(new_n976), .ZN(new_n1118));
  OAI211_X1 g693(.A(KEYINPUT121), .B(new_n1068), .C1(new_n1118), .C2(new_n1111), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1114), .B2(new_n1067), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1115), .A2(KEYINPUT51), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G8), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1116), .B1(new_n1114), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT51), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1117), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1110), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1003), .A2(new_n1010), .A3(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1083), .A2(new_n1085), .A3(new_n693), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1073), .B(KEYINPUT112), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1091), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1093), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1102), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1093), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1111), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1067), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(G168), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1135), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT116), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1093), .A2(new_n1102), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1145));
  OAI21_X1  g720(.A(G8), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(new_n1096), .B2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1141), .A2(new_n1142), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1134), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1117), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1107), .B1(new_n994), .B2(new_n999), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1127), .A2(new_n1151), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1150), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1122), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1139), .B2(KEYINPUT121), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1160), .A2(new_n1121), .B1(KEYINPUT51), .B2(new_n1125), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT62), .B1(new_n1161), .B2(new_n1117), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1136), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1163));
  AND4_X1   g738(.A1(new_n1150), .A2(new_n1162), .A3(new_n1157), .A4(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1129), .B(new_n1149), .C1(new_n1158), .C2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1030), .A2(new_n958), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n771), .B(new_n1011), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n753), .B(new_n1031), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n715), .B(new_n719), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1167), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n704), .A2(new_n706), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(KEYINPUT107), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n704), .A2(new_n706), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1167), .B1(new_n1174), .B2(KEYINPUT107), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1173), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1165), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1167), .B1(new_n1168), .B2(new_n754), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT127), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1166), .A2(new_n1031), .ZN(new_n1183));
  XNOR2_X1  g758(.A(KEYINPUT126), .B(KEYINPUT46), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1182), .B(new_n1185), .C1(new_n1183), .C2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g762(.A(new_n1187), .B(KEYINPUT47), .Z(new_n1188));
  NOR2_X1   g763(.A1(new_n1176), .A2(new_n1167), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT48), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1190), .A2(new_n1173), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n716), .A2(new_n719), .ZN(new_n1192));
  OAI22_X1  g767(.A1(new_n1170), .A2(new_n1192), .B1(G2067), .B2(new_n771), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1193), .A2(new_n1166), .ZN(new_n1194));
  NOR3_X1   g769(.A1(new_n1188), .A2(new_n1191), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1180), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g771(.A1(new_n648), .A2(G319), .A3(new_n665), .ZN(new_n1198));
  OR2_X1    g772(.A1(G229), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g773(.A(new_n1199), .B1(new_n879), .B2(new_n885), .ZN(new_n1200));
  AND2_X1   g774(.A1(new_n1200), .A2(new_n949), .ZN(G308));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n949), .ZN(G225));
endmodule


