

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U553 ( .A(n714), .B(KEYINPUT97), .ZN(n806) );
  XOR2_X1 U554 ( .A(KEYINPUT17), .B(n516), .Z(n887) );
  NOR2_X1 U555 ( .A1(n520), .A2(G2104), .ZN(n884) );
  INV_X1 U556 ( .A(KEYINPUT107), .ZN(n741) );
  NOR2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n516) );
  AND2_X1 U558 ( .A1(n537), .A2(n536), .ZN(G160) );
  OR2_X1 U559 ( .A1(n739), .A2(n738), .ZN(n514) );
  XNOR2_X1 U560 ( .A(KEYINPUT32), .B(n734), .ZN(n515) );
  INV_X1 U561 ( .A(n727), .ZN(n708) );
  INV_X1 U562 ( .A(KEYINPUT28), .ZN(n686) );
  NOR2_X1 U563 ( .A1(n721), .A2(n720), .ZN(n722) );
  AND2_X1 U564 ( .A1(n733), .A2(n732), .ZN(n734) );
  INV_X1 U565 ( .A(n979), .ZN(n743) );
  NOR2_X1 U566 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U567 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U568 ( .A1(G651), .A2(n618), .ZN(n646) );
  AND2_X1 U569 ( .A1(G138), .A2(n887), .ZN(n518) );
  AND2_X1 U570 ( .A1(n822), .A2(n821), .ZN(n823) );
  INV_X1 U571 ( .A(KEYINPUT89), .ZN(n517) );
  XNOR2_X1 U572 ( .A(n518), .B(n517), .ZN(n526) );
  INV_X1 U573 ( .A(G2105), .ZN(n520) );
  NAND2_X1 U574 ( .A1(G126), .A2(n884), .ZN(n519) );
  XNOR2_X1 U575 ( .A(n519), .B(KEYINPUT88), .ZN(n524) );
  AND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NAND2_X1 U577 ( .A1(G114), .A2(n883), .ZN(n522) );
  AND2_X1 U578 ( .A1(n520), .A2(G2104), .ZN(n888) );
  NAND2_X1 U579 ( .A1(G102), .A2(n888), .ZN(n521) );
  AND2_X1 U580 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U582 ( .A1(n526), .A2(n525), .ZN(G164) );
  NAND2_X1 U583 ( .A1(n883), .A2(G113), .ZN(n528) );
  NAND2_X1 U584 ( .A1(n887), .A2(G137), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U586 ( .A1(n529), .A2(KEYINPUT65), .ZN(n531) );
  OR2_X1 U587 ( .A1(n529), .A2(KEYINPUT65), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n531), .A2(n530), .ZN(n537) );
  AND2_X1 U589 ( .A1(G125), .A2(n884), .ZN(n535) );
  NAND2_X1 U590 ( .A1(G101), .A2(n888), .ZN(n532) );
  XNOR2_X1 U591 ( .A(n532), .B(KEYINPUT23), .ZN(n533) );
  XNOR2_X1 U592 ( .A(n533), .B(KEYINPUT64), .ZN(n534) );
  NOR2_X1 U593 ( .A1(n535), .A2(n534), .ZN(n536) );
  INV_X1 U594 ( .A(G651), .ZN(n541) );
  NOR2_X1 U595 ( .A1(G543), .A2(n541), .ZN(n538) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n538), .Z(n638) );
  NAND2_X1 U597 ( .A1(G64), .A2(n638), .ZN(n540) );
  XOR2_X1 U598 ( .A(KEYINPUT0), .B(G543), .Z(n618) );
  NAND2_X1 U599 ( .A1(G52), .A2(n646), .ZN(n539) );
  NAND2_X1 U600 ( .A1(n540), .A2(n539), .ZN(n546) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U602 ( .A1(G90), .A2(n639), .ZN(n543) );
  NOR2_X1 U603 ( .A1(n618), .A2(n541), .ZN(n642) );
  NAND2_X1 U604 ( .A1(G77), .A2(n642), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n544), .Z(n545) );
  NOR2_X1 U607 ( .A1(n546), .A2(n545), .ZN(G171) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U609 ( .A1(G123), .A2(n884), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT78), .ZN(n548) );
  XNOR2_X1 U611 ( .A(n548), .B(KEYINPUT18), .ZN(n550) );
  NAND2_X1 U612 ( .A1(G111), .A2(n883), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G135), .A2(n887), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G99), .A2(n888), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n926) );
  XNOR2_X1 U618 ( .A(n926), .B(G2096), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n555), .B(KEYINPUT79), .ZN(n556) );
  OR2_X1 U620 ( .A1(G2100), .A2(n556), .ZN(G156) );
  INV_X1 U621 ( .A(G82), .ZN(G220) );
  NAND2_X1 U622 ( .A1(n639), .A2(G89), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT4), .B(n557), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n642), .A2(G76), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT75), .B(n558), .Z(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT5), .ZN(n566) );
  NAND2_X1 U628 ( .A1(G63), .A2(n638), .ZN(n563) );
  NAND2_X1 U629 ( .A1(G51), .A2(n646), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT10), .ZN(n569) );
  XNOR2_X1 U637 ( .A(KEYINPUT70), .B(n569), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n835) );
  NAND2_X1 U639 ( .A1(n835), .A2(G567), .ZN(n570) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U641 ( .A1(G56), .A2(n638), .ZN(n571) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n571), .Z(n578) );
  NAND2_X1 U643 ( .A1(G81), .A2(n639), .ZN(n572) );
  XOR2_X1 U644 ( .A(KEYINPUT71), .B(n572), .Z(n573) );
  XNOR2_X1 U645 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G68), .A2(n642), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n646), .A2(G43), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n973) );
  INV_X1 U652 ( .A(G860), .ZN(n602) );
  OR2_X1 U653 ( .A1(n973), .A2(n602), .ZN(G153) );
  XOR2_X1 U654 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U655 ( .A1(G66), .A2(n638), .ZN(n582) );
  NAND2_X1 U656 ( .A1(G92), .A2(n639), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U658 ( .A1(G79), .A2(n642), .ZN(n584) );
  NAND2_X1 U659 ( .A1(G54), .A2(n646), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U662 ( .A(KEYINPUT15), .B(n587), .Z(n976) );
  INV_X1 U663 ( .A(n976), .ZN(n844) );
  INV_X1 U664 ( .A(G868), .ZN(n658) );
  NAND2_X1 U665 ( .A1(n844), .A2(n658), .ZN(n588) );
  XNOR2_X1 U666 ( .A(KEYINPUT74), .B(n588), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n589) );
  XOR2_X1 U668 ( .A(KEYINPUT73), .B(n589), .Z(n590) );
  NAND2_X1 U669 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U670 ( .A1(G65), .A2(n638), .ZN(n593) );
  NAND2_X1 U671 ( .A1(G53), .A2(n646), .ZN(n592) );
  NAND2_X1 U672 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U673 ( .A1(G91), .A2(n639), .ZN(n595) );
  NAND2_X1 U674 ( .A1(G78), .A2(n642), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U676 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U677 ( .A(n598), .B(KEYINPUT67), .ZN(G299) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n599) );
  XNOR2_X1 U679 ( .A(n599), .B(KEYINPUT76), .ZN(n601) );
  NOR2_X1 U680 ( .A1(n658), .A2(G286), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n603), .A2(n976), .ZN(n604) );
  XNOR2_X1 U684 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n973), .ZN(n605) );
  XOR2_X1 U686 ( .A(KEYINPUT77), .B(n605), .Z(n608) );
  NAND2_X1 U687 ( .A1(G868), .A2(n976), .ZN(n606) );
  NOR2_X1 U688 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U689 ( .A1(n608), .A2(n607), .ZN(G282) );
  XNOR2_X1 U690 ( .A(n973), .B(KEYINPUT80), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n976), .A2(G559), .ZN(n609) );
  XNOR2_X1 U692 ( .A(n610), .B(n609), .ZN(n655) );
  NOR2_X1 U693 ( .A1(G860), .A2(n655), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G67), .A2(n638), .ZN(n612) );
  NAND2_X1 U695 ( .A1(G93), .A2(n639), .ZN(n611) );
  NAND2_X1 U696 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G80), .A2(n642), .ZN(n614) );
  NAND2_X1 U698 ( .A1(G55), .A2(n646), .ZN(n613) );
  NAND2_X1 U699 ( .A1(n614), .A2(n613), .ZN(n615) );
  OR2_X1 U700 ( .A1(n616), .A2(n615), .ZN(n659) );
  XOR2_X1 U701 ( .A(n617), .B(n659), .Z(G145) );
  NAND2_X1 U702 ( .A1(G49), .A2(n646), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G87), .A2(n618), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U705 ( .A1(n638), .A2(n621), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n622) );
  XOR2_X1 U707 ( .A(KEYINPUT81), .B(n622), .Z(n623) );
  NAND2_X1 U708 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U709 ( .A1(G60), .A2(n638), .ZN(n626) );
  NAND2_X1 U710 ( .A1(G85), .A2(n639), .ZN(n625) );
  NAND2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n642), .A2(G72), .ZN(n627) );
  XOR2_X1 U713 ( .A(KEYINPUT66), .B(n627), .Z(n628) );
  NOR2_X1 U714 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n646), .A2(G47), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G88), .A2(n639), .ZN(n633) );
  NAND2_X1 U718 ( .A1(G75), .A2(n642), .ZN(n632) );
  NAND2_X1 U719 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U720 ( .A1(G62), .A2(n638), .ZN(n635) );
  NAND2_X1 U721 ( .A1(G50), .A2(n646), .ZN(n634) );
  NAND2_X1 U722 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U723 ( .A1(n637), .A2(n636), .ZN(G166) );
  NAND2_X1 U724 ( .A1(G61), .A2(n638), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G86), .A2(n639), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n642), .A2(G73), .ZN(n643) );
  XOR2_X1 U728 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n646), .A2(G48), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n648), .A2(n647), .ZN(G305) );
  XOR2_X1 U732 ( .A(n659), .B(G288), .Z(n654) );
  XOR2_X1 U733 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n650) );
  INV_X1 U734 ( .A(G299), .ZN(n970) );
  XNOR2_X1 U735 ( .A(n970), .B(G166), .ZN(n649) );
  XNOR2_X1 U736 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U737 ( .A(n651), .B(G305), .Z(n652) );
  XNOR2_X1 U738 ( .A(G290), .B(n652), .ZN(n653) );
  XNOR2_X1 U739 ( .A(n654), .B(n653), .ZN(n841) );
  XNOR2_X1 U740 ( .A(n841), .B(n655), .ZN(n656) );
  NAND2_X1 U741 ( .A1(n656), .A2(G868), .ZN(n657) );
  XOR2_X1 U742 ( .A(KEYINPUT83), .B(n657), .Z(n661) );
  NAND2_X1 U743 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n665), .A2(G2072), .ZN(n666) );
  XNOR2_X1 U750 ( .A(KEYINPUT84), .B(n666), .ZN(G158) );
  XNOR2_X1 U751 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U753 ( .A(KEYINPUT68), .B(G57), .Z(G237) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n668) );
  XNOR2_X1 U755 ( .A(KEYINPUT22), .B(KEYINPUT85), .ZN(n667) );
  XNOR2_X1 U756 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U757 ( .A1(n669), .A2(G218), .ZN(n670) );
  XNOR2_X1 U758 ( .A(KEYINPUT86), .B(n670), .ZN(n671) );
  NAND2_X1 U759 ( .A1(n671), .A2(G96), .ZN(n840) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n840), .ZN(n675) );
  NAND2_X1 U761 ( .A1(G108), .A2(G120), .ZN(n672) );
  NOR2_X1 U762 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U763 ( .A1(G69), .A2(n673), .ZN(n839) );
  NAND2_X1 U764 ( .A1(G567), .A2(n839), .ZN(n674) );
  NAND2_X1 U765 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U766 ( .A(KEYINPUT87), .B(n676), .ZN(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n678) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n677) );
  NOR2_X1 U769 ( .A1(n678), .A2(n677), .ZN(n838) );
  NAND2_X1 U770 ( .A1(n838), .A2(G36), .ZN(G176) );
  XOR2_X1 U771 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n776) );
  AND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n679) );
  NAND2_X2 U774 ( .A1(n776), .A2(n679), .ZN(n727) );
  NAND2_X1 U775 ( .A1(G2072), .A2(n708), .ZN(n680) );
  XNOR2_X1 U776 ( .A(n680), .B(KEYINPUT27), .ZN(n682) );
  INV_X1 U777 ( .A(KEYINPUT101), .ZN(n681) );
  XNOR2_X1 U778 ( .A(n682), .B(n681), .ZN(n685) );
  XOR2_X1 U779 ( .A(G1956), .B(KEYINPUT102), .Z(n997) );
  NOR2_X1 U780 ( .A1(n708), .A2(n997), .ZN(n683) );
  XOR2_X1 U781 ( .A(KEYINPUT103), .B(n683), .Z(n684) );
  NOR2_X1 U782 ( .A1(n685), .A2(n684), .ZN(n688) );
  NOR2_X1 U783 ( .A1(n970), .A2(n688), .ZN(n687) );
  XNOR2_X1 U784 ( .A(n687), .B(n686), .ZN(n704) );
  NAND2_X1 U785 ( .A1(n970), .A2(n688), .ZN(n702) );
  NAND2_X1 U786 ( .A1(G1348), .A2(n727), .ZN(n690) );
  NAND2_X1 U787 ( .A1(n708), .A2(G2067), .ZN(n689) );
  NAND2_X1 U788 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U789 ( .A(KEYINPUT104), .B(n691), .Z(n698) );
  OR2_X1 U790 ( .A1(n976), .A2(n698), .ZN(n697) );
  INV_X1 U791 ( .A(G1996), .ZN(n946) );
  NOR2_X1 U792 ( .A1(n727), .A2(n946), .ZN(n692) );
  XOR2_X1 U793 ( .A(n692), .B(KEYINPUT26), .Z(n694) );
  NAND2_X1 U794 ( .A1(n727), .A2(G1341), .ZN(n693) );
  NAND2_X1 U795 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U796 ( .A1(n973), .A2(n695), .ZN(n696) );
  NAND2_X1 U797 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n698), .A2(n976), .ZN(n699) );
  AND2_X1 U799 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n706) );
  XNOR2_X1 U802 ( .A(KEYINPUT105), .B(KEYINPUT29), .ZN(n705) );
  XNOR2_X1 U803 ( .A(n706), .B(n705), .ZN(n713) );
  XOR2_X1 U804 ( .A(G2078), .B(KEYINPUT25), .Z(n707) );
  XNOR2_X1 U805 ( .A(KEYINPUT99), .B(n707), .ZN(n945) );
  NAND2_X1 U806 ( .A1(n708), .A2(n945), .ZN(n709) );
  XNOR2_X1 U807 ( .A(n709), .B(KEYINPUT100), .ZN(n711) );
  INV_X1 U808 ( .A(G1961), .ZN(n991) );
  NAND2_X1 U809 ( .A1(n991), .A2(n727), .ZN(n710) );
  NAND2_X1 U810 ( .A1(n711), .A2(n710), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n719), .A2(G171), .ZN(n712) );
  NAND2_X1 U812 ( .A1(n713), .A2(n712), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n727), .A2(G8), .ZN(n714) );
  INV_X1 U814 ( .A(n806), .ZN(n810) );
  NOR2_X1 U815 ( .A1(n810), .A2(G1966), .ZN(n739) );
  INV_X1 U816 ( .A(G8), .ZN(n715) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n727), .ZN(n735) );
  OR2_X1 U818 ( .A1(n715), .A2(n735), .ZN(n716) );
  OR2_X1 U819 ( .A1(n739), .A2(n716), .ZN(n717) );
  XNOR2_X1 U820 ( .A(n717), .B(KEYINPUT30), .ZN(n718) );
  NOR2_X1 U821 ( .A1(G168), .A2(n718), .ZN(n721) );
  NOR2_X1 U822 ( .A1(G171), .A2(n719), .ZN(n720) );
  XOR2_X1 U823 ( .A(KEYINPUT31), .B(n722), .Z(n723) );
  NAND2_X1 U824 ( .A1(n724), .A2(n723), .ZN(n737) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n725) );
  NAND2_X1 U826 ( .A1(n737), .A2(n725), .ZN(n733) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n810), .ZN(n726) );
  XNOR2_X1 U828 ( .A(n726), .B(KEYINPUT106), .ZN(n729) );
  NOR2_X1 U829 ( .A1(n727), .A2(G2090), .ZN(n728) );
  NOR2_X1 U830 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U831 ( .A1(G303), .A2(n730), .ZN(n731) );
  OR2_X1 U832 ( .A1(n715), .A2(n731), .ZN(n732) );
  NAND2_X1 U833 ( .A1(G8), .A2(n735), .ZN(n736) );
  NAND2_X1 U834 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U835 ( .A1(n515), .A2(n514), .ZN(n800) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U837 ( .A1(G303), .A2(G1971), .ZN(n740) );
  NOR2_X1 U838 ( .A1(n749), .A2(n740), .ZN(n971) );
  NAND2_X1 U839 ( .A1(n800), .A2(n971), .ZN(n742) );
  XNOR2_X1 U840 ( .A(n742), .B(n741), .ZN(n746) );
  NAND2_X1 U841 ( .A1(n806), .A2(KEYINPUT108), .ZN(n744) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n979) );
  NOR2_X1 U843 ( .A1(KEYINPUT33), .A2(n747), .ZN(n755) );
  INV_X1 U844 ( .A(KEYINPUT108), .ZN(n748) );
  NAND2_X1 U845 ( .A1(n748), .A2(n749), .ZN(n752) );
  NAND2_X1 U846 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NAND2_X1 U847 ( .A1(n750), .A2(KEYINPUT108), .ZN(n751) );
  NAND2_X1 U848 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U849 ( .A1(n810), .A2(n753), .ZN(n754) );
  NOR2_X1 U850 ( .A1(n755), .A2(n754), .ZN(n779) );
  XOR2_X1 U851 ( .A(G1981), .B(G305), .Z(n967) );
  NAND2_X1 U852 ( .A1(G107), .A2(n883), .ZN(n757) );
  NAND2_X1 U853 ( .A1(G119), .A2(n884), .ZN(n756) );
  NAND2_X1 U854 ( .A1(n757), .A2(n756), .ZN(n760) );
  NAND2_X1 U855 ( .A1(G131), .A2(n887), .ZN(n758) );
  XNOR2_X1 U856 ( .A(KEYINPUT93), .B(n758), .ZN(n759) );
  NOR2_X1 U857 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U858 ( .A1(n888), .A2(G95), .ZN(n761) );
  NAND2_X1 U859 ( .A1(n762), .A2(n761), .ZN(n894) );
  NAND2_X1 U860 ( .A1(G1991), .A2(n894), .ZN(n763) );
  XOR2_X1 U861 ( .A(KEYINPUT94), .B(n763), .Z(n774) );
  NAND2_X1 U862 ( .A1(G105), .A2(n888), .ZN(n764) );
  XNOR2_X1 U863 ( .A(n764), .B(KEYINPUT38), .ZN(n771) );
  NAND2_X1 U864 ( .A1(G141), .A2(n887), .ZN(n766) );
  NAND2_X1 U865 ( .A1(G117), .A2(n883), .ZN(n765) );
  NAND2_X1 U866 ( .A1(n766), .A2(n765), .ZN(n769) );
  NAND2_X1 U867 ( .A1(G129), .A2(n884), .ZN(n767) );
  XNOR2_X1 U868 ( .A(KEYINPUT95), .B(n767), .ZN(n768) );
  NOR2_X1 U869 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U870 ( .A1(n771), .A2(n770), .ZN(n898) );
  NAND2_X1 U871 ( .A1(G1996), .A2(n898), .ZN(n772) );
  XOR2_X1 U872 ( .A(KEYINPUT96), .B(n772), .Z(n773) );
  NOR2_X1 U873 ( .A1(n774), .A2(n773), .ZN(n922) );
  XOR2_X1 U874 ( .A(G1986), .B(G290), .Z(n980) );
  NAND2_X1 U875 ( .A1(n922), .A2(n980), .ZN(n777) );
  NAND2_X1 U876 ( .A1(G160), .A2(G40), .ZN(n775) );
  NOR2_X1 U877 ( .A1(n776), .A2(n775), .ZN(n820) );
  NAND2_X1 U878 ( .A1(n777), .A2(n820), .ZN(n799) );
  AND2_X1 U879 ( .A1(n967), .A2(n799), .ZN(n778) );
  NAND2_X1 U880 ( .A1(n779), .A2(n778), .ZN(n818) );
  NOR2_X1 U881 ( .A1(G1996), .A2(n898), .ZN(n919) );
  INV_X1 U882 ( .A(n922), .ZN(n782) );
  NOR2_X1 U883 ( .A1(G1986), .A2(G290), .ZN(n780) );
  NOR2_X1 U884 ( .A1(G1991), .A2(n894), .ZN(n927) );
  NOR2_X1 U885 ( .A1(n780), .A2(n927), .ZN(n781) );
  NOR2_X1 U886 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U887 ( .A1(n919), .A2(n783), .ZN(n784) );
  XNOR2_X1 U888 ( .A(KEYINPUT39), .B(n784), .ZN(n785) );
  NAND2_X1 U889 ( .A1(n785), .A2(n820), .ZN(n798) );
  XOR2_X1 U890 ( .A(G2067), .B(KEYINPUT37), .Z(n819) );
  NAND2_X1 U891 ( .A1(G140), .A2(n887), .ZN(n787) );
  NAND2_X1 U892 ( .A1(G104), .A2(n888), .ZN(n786) );
  NAND2_X1 U893 ( .A1(n787), .A2(n786), .ZN(n789) );
  XOR2_X1 U894 ( .A(KEYINPUT91), .B(KEYINPUT34), .Z(n788) );
  XNOR2_X1 U895 ( .A(n789), .B(n788), .ZN(n794) );
  NAND2_X1 U896 ( .A1(G116), .A2(n883), .ZN(n791) );
  NAND2_X1 U897 ( .A1(G128), .A2(n884), .ZN(n790) );
  NAND2_X1 U898 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U899 ( .A(KEYINPUT35), .B(n792), .Z(n793) );
  NOR2_X1 U900 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U901 ( .A(n795), .B(KEYINPUT36), .ZN(n796) );
  XOR2_X1 U902 ( .A(n796), .B(KEYINPUT92), .Z(n907) );
  NOR2_X1 U903 ( .A1(n819), .A2(n907), .ZN(n924) );
  NAND2_X1 U904 ( .A1(n924), .A2(n820), .ZN(n797) );
  AND2_X1 U905 ( .A1(n798), .A2(n797), .ZN(n816) );
  INV_X1 U906 ( .A(n799), .ZN(n814) );
  INV_X1 U907 ( .A(n800), .ZN(n804) );
  INV_X1 U908 ( .A(G2090), .ZN(n801) );
  NAND2_X1 U909 ( .A1(G8), .A2(n801), .ZN(n802) );
  NOR2_X1 U910 ( .A1(n802), .A2(G303), .ZN(n803) );
  NOR2_X1 U911 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U912 ( .A1(n806), .A2(n805), .ZN(n812) );
  NOR2_X1 U913 ( .A1(G1981), .A2(G305), .ZN(n807) );
  XOR2_X1 U914 ( .A(n807), .B(KEYINPUT24), .Z(n808) );
  XNOR2_X1 U915 ( .A(KEYINPUT98), .B(n808), .ZN(n809) );
  NOR2_X1 U916 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U917 ( .A1(n812), .A2(n811), .ZN(n813) );
  OR2_X1 U918 ( .A1(n814), .A2(n813), .ZN(n815) );
  AND2_X1 U919 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U920 ( .A1(n818), .A2(n817), .ZN(n822) );
  AND2_X1 U921 ( .A1(n907), .A2(n819), .ZN(n925) );
  NAND2_X1 U922 ( .A1(n925), .A2(n820), .ZN(n821) );
  XNOR2_X1 U923 ( .A(n823), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U924 ( .A(G2443), .B(G2435), .ZN(n833) );
  XOR2_X1 U925 ( .A(G2454), .B(G2430), .Z(n825) );
  XNOR2_X1 U926 ( .A(G2446), .B(KEYINPUT109), .ZN(n824) );
  XNOR2_X1 U927 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U928 ( .A(G2451), .B(G2427), .Z(n827) );
  XNOR2_X1 U929 ( .A(G1341), .B(G1348), .ZN(n826) );
  XNOR2_X1 U930 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U931 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U932 ( .A(G2438), .B(KEYINPUT110), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U935 ( .A1(n834), .A2(G14), .ZN(n913) );
  XNOR2_X1 U936 ( .A(KEYINPUT111), .B(n913), .ZN(G401) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U939 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U941 ( .A1(n838), .A2(n837), .ZN(G188) );
  XOR2_X1 U942 ( .A(G96), .B(KEYINPUT112), .Z(G221) );
  INV_X1 U944 ( .A(G120), .ZN(G236) );
  INV_X1 U945 ( .A(G108), .ZN(G238) );
  INV_X1 U946 ( .A(G69), .ZN(G235) );
  NOR2_X1 U947 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U948 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U949 ( .A(G286), .B(n841), .ZN(n843) );
  XNOR2_X1 U950 ( .A(n973), .B(G171), .ZN(n842) );
  XNOR2_X1 U951 ( .A(n843), .B(n842), .ZN(n846) );
  XOR2_X1 U952 ( .A(n844), .B(KEYINPUT119), .Z(n845) );
  XNOR2_X1 U953 ( .A(n846), .B(n845), .ZN(n847) );
  NOR2_X1 U954 ( .A1(G37), .A2(n847), .ZN(G397) );
  XOR2_X1 U955 ( .A(KEYINPUT113), .B(G2078), .Z(n849) );
  XNOR2_X1 U956 ( .A(G2072), .B(G2067), .ZN(n848) );
  XNOR2_X1 U957 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U958 ( .A(n850), .B(G2100), .Z(n852) );
  XNOR2_X1 U959 ( .A(G2084), .B(G2090), .ZN(n851) );
  XNOR2_X1 U960 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U961 ( .A(G2096), .B(KEYINPUT43), .Z(n854) );
  XNOR2_X1 U962 ( .A(KEYINPUT42), .B(G2678), .ZN(n853) );
  XNOR2_X1 U963 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U964 ( .A(n856), .B(n855), .Z(G227) );
  XOR2_X1 U965 ( .A(G1986), .B(G1991), .Z(n858) );
  XNOR2_X1 U966 ( .A(G1996), .B(G1971), .ZN(n857) );
  XNOR2_X1 U967 ( .A(n858), .B(n857), .ZN(n868) );
  XOR2_X1 U968 ( .A(KEYINPUT116), .B(G2474), .Z(n860) );
  XNOR2_X1 U969 ( .A(G1956), .B(KEYINPUT114), .ZN(n859) );
  XNOR2_X1 U970 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U971 ( .A(G1976), .B(G1981), .Z(n862) );
  XNOR2_X1 U972 ( .A(G1966), .B(G1961), .ZN(n861) );
  XNOR2_X1 U973 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U974 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U975 ( .A(KEYINPUT41), .B(KEYINPUT115), .ZN(n865) );
  XNOR2_X1 U976 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U977 ( .A(n868), .B(n867), .ZN(G229) );
  NAND2_X1 U978 ( .A1(G124), .A2(n884), .ZN(n869) );
  XNOR2_X1 U979 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U980 ( .A1(n883), .A2(G112), .ZN(n870) );
  NAND2_X1 U981 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U982 ( .A1(G136), .A2(n887), .ZN(n873) );
  NAND2_X1 U983 ( .A1(G100), .A2(n888), .ZN(n872) );
  NAND2_X1 U984 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U985 ( .A1(n875), .A2(n874), .ZN(G162) );
  NAND2_X1 U986 ( .A1(G139), .A2(n887), .ZN(n877) );
  NAND2_X1 U987 ( .A1(G103), .A2(n888), .ZN(n876) );
  NAND2_X1 U988 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U989 ( .A1(G115), .A2(n883), .ZN(n879) );
  NAND2_X1 U990 ( .A1(G127), .A2(n884), .ZN(n878) );
  NAND2_X1 U991 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U993 ( .A1(n882), .A2(n881), .ZN(n930) );
  NAND2_X1 U994 ( .A1(G118), .A2(n883), .ZN(n886) );
  NAND2_X1 U995 ( .A1(G130), .A2(n884), .ZN(n885) );
  NAND2_X1 U996 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U997 ( .A1(G142), .A2(n887), .ZN(n890) );
  NAND2_X1 U998 ( .A1(G106), .A2(n888), .ZN(n889) );
  NAND2_X1 U999 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U1000 ( .A(n891), .B(KEYINPUT45), .Z(n892) );
  NOR2_X1 U1001 ( .A1(n893), .A2(n892), .ZN(n895) );
  XNOR2_X1 U1002 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U1003 ( .A(n930), .B(n896), .ZN(n906) );
  XOR2_X1 U1004 ( .A(KEYINPUT118), .B(KEYINPUT48), .Z(n897) );
  XNOR2_X1 U1005 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U1006 ( .A(n899), .B(KEYINPUT117), .Z(n901) );
  XNOR2_X1 U1007 ( .A(G164), .B(KEYINPUT46), .ZN(n900) );
  XNOR2_X1 U1008 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1009 ( .A(n902), .B(n926), .Z(n904) );
  XNOR2_X1 U1010 ( .A(G160), .B(G162), .ZN(n903) );
  XNOR2_X1 U1011 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1012 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1013 ( .A(n908), .B(n907), .Z(n909) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n909), .ZN(G395) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n910) );
  XOR2_X1 U1016 ( .A(KEYINPUT49), .B(n910), .Z(n911) );
  XNOR2_X1 U1017 ( .A(n911), .B(KEYINPUT121), .ZN(n912) );
  NOR2_X1 U1018 ( .A1(G397), .A2(n912), .ZN(n917) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1020 ( .A(KEYINPUT120), .B(n914), .ZN(n915) );
  NOR2_X1 U1021 ( .A1(G395), .A2(n915), .ZN(n916) );
  NAND2_X1 U1022 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1025 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n920), .Z(n921) );
  XNOR2_X1 U1027 ( .A(KEYINPUT122), .B(n921), .ZN(n923) );
  NAND2_X1 U1028 ( .A1(n923), .A2(n922), .ZN(n940) );
  NOR2_X1 U1029 ( .A1(n925), .A2(n924), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(G160), .B(G2084), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G2072), .B(n930), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(G164), .B(G2078), .ZN(n931) );
  NAND2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1036 ( .A(KEYINPUT50), .B(n933), .Z(n934) );
  XNOR2_X1 U1037 ( .A(KEYINPUT123), .B(n934), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n941), .ZN(n942) );
  XOR2_X1 U1042 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n963) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n963), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n943), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G35), .ZN(n958) );
  XOR2_X1 U1046 ( .A(G2072), .B(G33), .Z(n944) );
  NAND2_X1 U1047 ( .A1(n944), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(n945), .B(G27), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(n946), .B(G32), .ZN(n947) );
  NAND2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(KEYINPUT125), .B(n949), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1053 ( .A(G1991), .B(G25), .ZN(n950) );
  NOR2_X1 U1054 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1062 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1063 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n966), .ZN(n1020) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G168), .ZN(n968) );
  NAND2_X1 U1068 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1069 ( .A(n969), .B(KEYINPUT57), .ZN(n988) );
  XNOR2_X1 U1070 ( .A(n970), .B(G1956), .ZN(n972) );
  NAND2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n986) );
  XNOR2_X1 U1072 ( .A(G1341), .B(n973), .ZN(n975) );
  XNOR2_X1 U1073 ( .A(G171), .B(n991), .ZN(n974) );
  NOR2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n976), .B(G1348), .ZN(n978) );
  NAND2_X1 U1076 ( .A1(G1971), .A2(G303), .ZN(n977) );
  NAND2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n1018) );
  INV_X1 U1084 ( .A(G16), .ZN(n1016) );
  XNOR2_X1 U1085 ( .A(n991), .B(G5), .ZN(n1012) );
  XOR2_X1 U1086 ( .A(G1966), .B(G21), .Z(n1003) );
  XNOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .ZN(n992) );
  XNOR2_X1 U1088 ( .A(n992), .B(G4), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n994) );
  XNOR2_X1 U1090 ( .A(G1981), .B(G6), .ZN(n993) );
  NOR2_X1 U1091 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n1000) );
  XOR2_X1 U1093 ( .A(G20), .B(n997), .Z(n998) );
  XNOR2_X1 U1094 ( .A(KEYINPUT126), .B(n998), .ZN(n999) );
  NOR2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1096 ( .A(KEYINPUT60), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1004) );
  NOR2_X1 U1100 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1101 ( .A(G1986), .B(G24), .Z(n1006) );
  NAND2_X1 U1102 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1104 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1106 ( .A(n1013), .B(KEYINPUT127), .ZN(n1014) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

