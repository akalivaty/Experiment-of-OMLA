//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n604, new_n605, new_n606, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n640, new_n641, new_n644, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT67), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT68), .B(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n465), .A2(new_n467), .A3(G137), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT71), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G137), .A4(new_n468), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT70), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n471), .A2(new_n478), .A3(G125), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AOI221_X4 g055(.A(new_n464), .B1(new_n470), .B2(new_n473), .C1(new_n480), .C2(G2105), .ZN(G160));
  NAND2_X1  g056(.A1(new_n471), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n474), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT73), .B(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n465), .A2(new_n467), .A3(G126), .A4(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT72), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n471), .A2(new_n496), .A3(G126), .A4(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n468), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT74), .A3(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT74), .A2(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n471), .A2(G138), .A3(new_n468), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  AND3_X1   g080(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(G543), .B1(KEYINPUT75), .B2(KEYINPUT5), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT76), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(new_n520), .A3(KEYINPUT76), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n506), .A2(new_n507), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(G651), .B1(G50), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n523), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  XNOR2_X1  g106(.A(KEYINPUT79), .B(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n512), .A2(new_n521), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(G51), .ZN(new_n537));
  NAND2_X1  g112(.A1(G63), .A2(G651), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(KEYINPUT77), .B1(new_n517), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n541));
  AOI211_X1 g116(.A(new_n541), .B(new_n538), .C1(new_n515), .C2(new_n516), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n537), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT78), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n539), .B1(new_n506), .B2(new_n507), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(new_n541), .ZN(new_n546));
  OAI211_X1 g121(.A(KEYINPUT77), .B(new_n539), .C1(new_n506), .C2(new_n507), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(new_n549), .A3(new_n537), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n536), .B1(new_n544), .B2(new_n550), .ZN(G168));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n525), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n528), .A2(G52), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n512), .A2(new_n521), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n515), .B2(new_n516), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT80), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n566), .B(new_n563), .C1(new_n525), .C2(new_n561), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n567), .A3(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT81), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n565), .A2(new_n567), .A3(new_n570), .A4(G651), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n569), .A2(new_n571), .B1(G43), .B2(new_n528), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT82), .B(G81), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n522), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G860), .ZN(G153));
  AND3_X1   g152(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G36), .ZN(G176));
  NAND2_X1  g154(.A1(G1), .A2(G3), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT8), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(G188));
  INV_X1    g157(.A(KEYINPUT85), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT84), .B1(new_n506), .B2(new_n507), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT84), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n515), .A2(new_n586), .A3(new_n516), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G65), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(G91), .A2(new_n522), .B1(new_n590), .B2(G651), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT83), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n528), .A2(new_n592), .A3(G53), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT9), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT9), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n528), .A2(new_n592), .A3(new_n595), .A4(G53), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n583), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n590), .A2(G651), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n512), .A2(G91), .A3(new_n521), .ZN(new_n600));
  AND4_X1   g175(.A1(new_n583), .A2(new_n599), .A3(new_n597), .A4(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G299));
  AND2_X1   g178(.A1(new_n533), .A2(new_n535), .ZN(new_n604));
  AOI221_X4 g179(.A(KEYINPUT78), .B1(G51), .B2(new_n528), .C1(new_n546), .C2(new_n547), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n549), .B1(new_n548), .B2(new_n537), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(G286));
  NAND3_X1  g182(.A1(new_n512), .A2(G87), .A3(new_n521), .ZN(new_n608));
  OAI21_X1  g183(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n528), .A2(G49), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(KEYINPUT86), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(KEYINPUT86), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(G288));
  NAND2_X1  g189(.A1(new_n522), .A2(G86), .ZN(new_n615));
  NAND2_X1  g190(.A1(G73), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G61), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n525), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n618), .A2(G651), .B1(G48), .B2(new_n528), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(G305));
  NAND2_X1  g195(.A1(new_n528), .A2(G47), .ZN(new_n621));
  INV_X1    g196(.A(G651), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n623));
  INV_X1    g198(.A(G85), .ZN(new_n624));
  OAI221_X1 g199(.A(new_n621), .B1(new_n622), .B2(new_n623), .C1(new_n557), .C2(new_n624), .ZN(G290));
  NAND2_X1  g200(.A1(G301), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n522), .B2(G92), .ZN(new_n628));
  INV_X1    g203(.A(G92), .ZN(new_n629));
  NOR3_X1   g204(.A1(new_n557), .A2(KEYINPUT10), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(G79), .A2(G543), .ZN(new_n632));
  INV_X1    g207(.A(G66), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n588), .B2(new_n633), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n634), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n626), .B1(new_n637), .B2(G868), .ZN(G284));
  OAI21_X1  g213(.A(new_n626), .B1(new_n637), .B2(G868), .ZN(G321));
  INV_X1    g214(.A(G868), .ZN(new_n640));
  NOR2_X1   g215(.A1(G286), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n602), .B2(new_n640), .ZN(G297));
  AOI21_X1  g217(.A(new_n641), .B1(new_n602), .B2(new_n640), .ZN(G280));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n637), .B1(new_n644), .B2(G860), .ZN(G148));
  NAND2_X1  g220(.A1(new_n575), .A2(new_n640), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n636), .A2(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n647), .B2(new_n640), .ZN(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n471), .A2(new_n462), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n483), .A2(G123), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n485), .A2(G135), .ZN(new_n656));
  NOR2_X1   g231(.A1(G99), .A2(G2105), .ZN(new_n657));
  OAI21_X1  g232(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n655), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(G2096), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n660), .ZN(G156));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2435), .ZN(new_n663));
  XOR2_X1   g238(.A(G2427), .B(G2438), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT14), .ZN(new_n666));
  XOR2_X1   g241(.A(G2451), .B(G2454), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1341), .B(G1348), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G14), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(KEYINPUT88), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n671), .A2(new_n678), .A3(new_n672), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G401));
  XNOR2_X1  g256(.A(G2084), .B(G2090), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT89), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2067), .B(G2678), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  OR3_X1    g263(.A1(new_n687), .A2(KEYINPUT18), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n683), .A2(new_n688), .A3(new_n685), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n684), .A2(new_n686), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(KEYINPUT17), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n687), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(KEYINPUT18), .B1(new_n687), .B2(new_n688), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n689), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT90), .B(G2096), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G2100), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(G227));
  XOR2_X1   g273(.A(G1961), .B(G1966), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  XOR2_X1   g275(.A(G1956), .B(G2474), .Z(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1971), .B(G1976), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT19), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n700), .A2(new_n701), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n705), .A2(new_n706), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n702), .A2(new_n707), .A3(new_n704), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n708), .B(new_n709), .C1(new_n706), .C2(new_n705), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n710), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT92), .B(G1986), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(G229));
  NAND2_X1  g293(.A1(new_n637), .A2(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G4), .B2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G1348), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NOR2_X1   g299(.A1(G164), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G27), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n722), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G29), .A2(G32), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n483), .A2(G129), .B1(new_n485), .B2(G141), .ZN(new_n729));
  INV_X1    g304(.A(G105), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n468), .A2(G2104), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT99), .B(KEYINPUT26), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n728), .B1(new_n736), .B2(G29), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT27), .B(G1996), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT100), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n737), .B(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(KEYINPUT24), .A2(G34), .ZN(new_n743));
  NOR2_X1   g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n743), .A2(new_n744), .A3(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n480), .A2(G2105), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n470), .A2(new_n473), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n746), .A2(new_n463), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n745), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT98), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G103), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT97), .B1(new_n731), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n462), .A2(new_n755), .A3(G103), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n754), .A2(new_n756), .A3(KEYINPUT25), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  INV_X1    g337(.A(G139), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n471), .A2(new_n468), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n762), .A2(new_n468), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(G29), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G33), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(G29), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2072), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n724), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n471), .A2(G128), .A3(G2105), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n471), .A2(G140), .A3(new_n468), .ZN(new_n774));
  OR2_X1    g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n775), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n772), .B1(new_n777), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2067), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(G28), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(G28), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n781), .A2(new_n782), .A3(new_n724), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n779), .B(new_n783), .C1(new_n724), .C2(new_n659), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n769), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n742), .A2(new_n752), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n720), .A2(new_n721), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n727), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G21), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G168), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT101), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1966), .ZN(new_n792));
  INV_X1    g367(.A(G16), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G5), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G171), .B2(new_n793), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1961), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n723), .B2(new_n726), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n750), .A2(new_n751), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n788), .A2(new_n792), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n793), .A2(G23), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n793), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT94), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT33), .B(G1976), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n803), .A2(new_n805), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n793), .B2(G22), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n808), .A2(new_n793), .A3(G22), .ZN(new_n810));
  AOI211_X1 g385(.A(new_n809), .B(new_n810), .C1(G303), .C2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1971), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n793), .A2(G6), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n615), .A2(new_n619), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n793), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT32), .B(G1981), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n806), .A2(new_n807), .A3(new_n812), .A4(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT34), .Z(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G24), .ZN(new_n820));
  XOR2_X1   g395(.A(G290), .B(KEYINPUT93), .Z(new_n821));
  AOI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(G16), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(G1986), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n483), .A2(G119), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n485), .A2(G131), .ZN(new_n825));
  NOR2_X1   g400(.A1(G95), .A2(G2105), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(new_n468), .B2(G107), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  MUX2_X1   g403(.A(G25), .B(new_n828), .S(G29), .Z(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT35), .B(G1991), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n829), .B(new_n830), .Z(new_n831));
  NAND3_X1  g406(.A1(new_n819), .A2(new_n823), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n819), .A2(new_n834), .A3(new_n823), .A4(new_n831), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n799), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n793), .A2(KEYINPUT23), .A3(G20), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT23), .ZN(new_n838));
  INV_X1    g413(.A(G20), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(G16), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n837), .B(new_n840), .C1(new_n602), .C2(new_n793), .ZN(new_n841));
  INV_X1    g416(.A(G1956), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n724), .A2(G35), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G162), .B2(new_n724), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT29), .B(G2090), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n793), .A2(G19), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n576), .B2(new_n793), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(G1341), .Z(new_n850));
  NAND4_X1  g425(.A1(new_n836), .A2(new_n843), .A3(new_n847), .A4(new_n850), .ZN(G150));
  INV_X1    g426(.A(G150), .ZN(G311));
  NAND2_X1  g427(.A1(new_n522), .A2(G93), .ZN(new_n853));
  NAND2_X1  g428(.A1(G80), .A2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G67), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n525), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n856), .A2(G651), .B1(G55), .B2(new_n528), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n644), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT39), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n862), .B(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n572), .A2(new_n574), .A3(new_n858), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n858), .B1(new_n572), .B2(new_n574), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n865), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n861), .B1(new_n870), .B2(G860), .ZN(G145));
  XOR2_X1   g446(.A(new_n828), .B(new_n652), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n483), .A2(G130), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n485), .A2(G142), .ZN(new_n874));
  OR2_X1    g449(.A1(G106), .A2(G2105), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n875), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n872), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n500), .A2(new_n880), .A3(new_n502), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n500), .B2(new_n502), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n498), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT105), .ZN(new_n884));
  INV_X1    g459(.A(new_n777), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n761), .B2(new_n765), .ZN(new_n886));
  NAND2_X1  g461(.A1(G115), .A2(G2104), .ZN(new_n887));
  INV_X1    g462(.A(G127), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n474), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n889), .A2(G2105), .B1(new_n485), .B2(G139), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n890), .A2(new_n760), .A3(new_n759), .A4(new_n777), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n893), .B(new_n498), .C1(new_n881), .C2(new_n882), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n884), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n892), .B1(new_n884), .B2(new_n894), .ZN(new_n897));
  INV_X1    g472(.A(new_n736), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n892), .ZN(new_n900));
  INV_X1    g475(.A(new_n882), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n500), .A2(new_n880), .A3(new_n502), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n893), .B1(new_n903), .B2(new_n498), .ZN(new_n904));
  INV_X1    g479(.A(new_n894), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n736), .B1(new_n906), .B2(new_n895), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n879), .B1(new_n899), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n872), .B(new_n877), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n898), .B1(new_n896), .B2(new_n897), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n736), .A3(new_n895), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n748), .B(new_n489), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n659), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n910), .A2(new_n911), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(new_n879), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n913), .B2(new_n918), .ZN(new_n921));
  INV_X1    g496(.A(new_n915), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT106), .B1(new_n908), .B2(new_n912), .ZN(new_n924));
  NOR4_X1   g499(.A1(new_n924), .A2(new_n920), .A3(KEYINPUT107), .A4(new_n915), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n916), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT108), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(new_n916), .C1(new_n923), .C2(new_n925), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n927), .A2(KEYINPUT40), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT40), .B1(new_n927), .B2(new_n929), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(G395));
  XNOR2_X1  g507(.A(new_n869), .B(new_n647), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n598), .B2(new_n601), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n591), .A2(new_n583), .A3(new_n597), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n599), .A2(new_n597), .A3(new_n600), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT85), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n938), .A3(KEYINPUT109), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(new_n636), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n602), .A2(new_n637), .A3(KEYINPUT109), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT41), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT41), .B1(new_n940), .B2(new_n941), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n933), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n946));
  INV_X1    g521(.A(new_n858), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n575), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n866), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(new_n647), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n940), .A2(new_n941), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n945), .A2(new_n946), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n946), .B1(new_n945), .B2(new_n952), .ZN(new_n954));
  XNOR2_X1  g529(.A(G303), .B(new_n801), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(G305), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(G290), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n953), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT41), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n951), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n950), .B1(new_n942), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n951), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n933), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT42), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n945), .A2(new_n946), .A3(new_n952), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n957), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(G868), .B1(new_n959), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n947), .A2(G868), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(G295));
  OAI21_X1  g546(.A(new_n958), .B1(new_n953), .B2(new_n954), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n965), .A2(new_n957), .A3(new_n966), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n640), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT110), .B1(new_n974), .B2(new_n969), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n968), .A2(new_n976), .A3(new_n970), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n975), .A2(new_n977), .ZN(G331));
  NAND2_X1  g553(.A1(new_n961), .A2(new_n942), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT112), .B1(G168), .B2(G301), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n982));
  NAND3_X1  g557(.A1(G286), .A2(new_n982), .A3(G171), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n604), .B(G301), .C1(new_n606), .C2(new_n605), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT111), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n987));
  NAND3_X1  g562(.A1(G168), .A2(new_n987), .A3(G301), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n949), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n984), .A2(new_n989), .A3(new_n948), .A4(new_n866), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n981), .A2(new_n983), .B1(new_n986), .B2(new_n988), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n869), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n993), .B2(new_n994), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n980), .A2(new_n993), .B1(new_n997), .B2(new_n963), .ZN(new_n998));
  AOI21_X1  g573(.A(G37), .B1(new_n998), .B2(new_n958), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(new_n993), .B2(new_n951), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n963), .A2(KEYINPUT114), .A3(new_n992), .A4(new_n991), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1001), .B(new_n1002), .C1(new_n997), .C2(new_n979), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1003), .A2(KEYINPUT115), .A3(new_n957), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT115), .B1(new_n1003), .B2(new_n957), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT43), .B(new_n999), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n980), .A2(new_n993), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n997), .A2(new_n963), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n958), .ZN(new_n1010));
  INV_X1    g585(.A(G37), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n998), .A2(new_n958), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1007), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1006), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT44), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1007), .B(new_n999), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT43), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1016), .A2(new_n1021), .ZN(G397));
  AOI21_X1  g597(.A(G1384), .B1(new_n884), .B2(new_n894), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(KEYINPUT45), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n746), .A2(G40), .A3(new_n463), .A4(new_n747), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G1996), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OR3_X1    g604(.A1(new_n1029), .A2(KEYINPUT116), .A3(new_n898), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1027), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n828), .A2(new_n830), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n828), .A2(new_n830), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G2067), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n777), .B(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1996), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1036), .B1(new_n736), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT116), .B1(new_n1029), .B2(new_n898), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1030), .A2(new_n1034), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(G290), .B(G1986), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1031), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1384), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n504), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1026), .B1(new_n1046), .B2(KEYINPUT45), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1023), .B2(KEYINPUT45), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n883), .A2(new_n1049), .A3(new_n1044), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(KEYINPUT50), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1026), .A3(new_n1051), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n1048), .A2(G1971), .B1(G2090), .B2(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G303), .A2(G8), .ZN(new_n1056));
  MUX2_X1   g631(.A(new_n1054), .B(new_n1055), .S(new_n1056), .Z(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(G8), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1023), .A2(KEYINPUT45), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1047), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n723), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  INV_X1    g637(.A(G1961), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1061), .A2(new_n1062), .B1(new_n1063), .B2(new_n1052), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n1044), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(G160), .A3(G40), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT45), .B1(new_n883), .B2(new_n1044), .ZN(new_n1067));
  OR4_X1    g642(.A1(new_n1062), .A2(new_n1066), .A3(new_n1067), .A4(G2078), .ZN(new_n1068));
  AOI21_X1  g643(.A(G301), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1025), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1384), .B1(new_n903), .B2(new_n498), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1049), .B2(new_n1071), .ZN(new_n1072));
  OAI22_X1  g647(.A1(new_n1048), .A2(G1971), .B1(new_n1072), .B2(G2090), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1057), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(G160), .A2(new_n883), .A3(G40), .A4(new_n1044), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n801), .A2(G1976), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(G8), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1976), .B1(new_n612), .B2(new_n613), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT52), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n1079), .B2(KEYINPUT52), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1981), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n615), .B2(new_n619), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT119), .B(G1981), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1087), .B(new_n1088), .C1(G305), .C2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G305), .A2(new_n1089), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT49), .B1(new_n1091), .B2(new_n1086), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1077), .A2(G8), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NOR4_X1   g670(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .A4(KEYINPUT52), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1084), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AND4_X1   g672(.A1(new_n1058), .A2(new_n1069), .A3(new_n1076), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1966), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1050), .A2(new_n1051), .A3(new_n751), .A4(new_n1026), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT120), .B(new_n1099), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G286), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT51), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1102), .A2(G168), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G8), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1108), .B2(G8), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT62), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1105), .B2(G286), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1109), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n1113), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1098), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT126), .B(new_n1098), .C1(new_n1115), .C2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1093), .A2(G1976), .A3(G288), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1094), .B1(new_n1125), .B2(new_n1091), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1081), .A2(KEYINPUT118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1127), .B(new_n1128), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1126), .B1(new_n1129), .B2(new_n1058), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1105), .A2(G8), .A3(G168), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1131), .A2(KEYINPUT63), .A3(new_n1058), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1053), .A2(G8), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1075), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1097), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1057), .B1(new_n1053), .B2(G8), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT121), .B1(new_n1129), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1132), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1097), .A2(new_n1076), .A3(new_n1058), .A4(new_n1131), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1130), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT56), .B(G2072), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1059), .A2(new_n1060), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1072), .A2(new_n842), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT57), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n937), .B(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1077), .B2(G2067), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1071), .A2(new_n1026), .A3(KEYINPUT122), .A4(new_n1035), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1052), .A2(new_n721), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT123), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1160), .A3(new_n1157), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1145), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n637), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1152), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n636), .B1(new_n1162), .B2(KEYINPUT60), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1156), .A2(new_n1160), .A3(new_n1157), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1160), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1168));
  OAI211_X1 g743(.A(KEYINPUT60), .B(new_n636), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1166), .A2(new_n1170), .B1(KEYINPUT60), .B2(new_n1162), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1077), .ZN(new_n1173));
  XNOR2_X1  g748(.A(KEYINPUT58), .B(G1341), .ZN(new_n1174));
  OAI22_X1  g749(.A1(new_n1172), .A2(G1996), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1175), .A2(new_n1176), .A3(new_n576), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1178), .B1(new_n1048), .B2(new_n1037), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT59), .B1(new_n1179), .B2(new_n575), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1163), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1149), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1152), .A2(KEYINPUT61), .A3(new_n1163), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1181), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1165), .B1(new_n1171), .B2(new_n1187), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1189));
  XOR2_X1   g764(.A(G301), .B(KEYINPUT54), .Z(new_n1190));
  OR2_X1    g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1097), .A2(new_n1076), .A3(new_n1058), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1026), .B1(new_n1023), .B2(KEYINPUT45), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(KEYINPUT125), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1195), .A2(KEYINPUT53), .A3(new_n723), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1059), .B1(new_n1194), .B2(KEYINPUT125), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1064), .B(new_n1190), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1143), .B1(new_n1188), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1043), .B1(new_n1124), .B2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1030), .A2(new_n1033), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n885), .A2(new_n1035), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1027), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1028), .A2(KEYINPUT46), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1028), .A2(KEYINPUT46), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1027), .B1(new_n736), .B2(new_n1036), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1027), .A2(G1986), .A3(G290), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT48), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1041), .A2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1204), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1201), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g789(.A(new_n459), .ZN(new_n1216));
  NOR2_X1   g790(.A1(G227), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n680), .A2(new_n717), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n1219));
  NOR2_X1   g793(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1220), .B1(new_n927), .B2(new_n929), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1222));
  AND3_X1   g796(.A1(new_n1221), .A2(new_n1019), .A3(new_n1222), .ZN(G308));
  NAND3_X1  g797(.A1(new_n1221), .A2(new_n1019), .A3(new_n1222), .ZN(G225));
endmodule


