

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U555 ( .A1(n753), .A2(n946), .ZN(n522) );
  OR2_X1 U556 ( .A1(n685), .A2(n684), .ZN(n794) );
  NOR2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n552) );
  XNOR2_X1 U558 ( .A(n522), .B(KEYINPUT101), .ZN(n757) );
  NAND2_X1 U559 ( .A1(n523), .A2(n709), .ZN(n712) );
  NAND2_X1 U560 ( .A1(n704), .A2(n705), .ZN(n523) );
  NAND2_X1 U561 ( .A1(n693), .A2(G2067), .ZN(n695) );
  XNOR2_X1 U562 ( .A(n715), .B(KEYINPUT92), .ZN(n693) );
  AND2_X1 U563 ( .A1(n795), .A2(n686), .ZN(n715) );
  NOR2_X2 U564 ( .A1(G2105), .A2(n555), .ZN(n560) );
  XNOR2_X1 U565 ( .A(KEYINPUT29), .B(KEYINPUT96), .ZN(n711) );
  XNOR2_X1 U566 ( .A(n712), .B(n711), .ZN(n738) );
  NAND2_X1 U567 ( .A1(G8), .A2(n740), .ZN(n778) );
  INV_X1 U568 ( .A(KEYINPUT102), .ZN(n820) );
  NOR2_X1 U569 ( .A1(n645), .A2(G651), .ZN(n646) );
  XOR2_X1 U570 ( .A(KEYINPUT0), .B(G543), .Z(n645) );
  NAND2_X1 U571 ( .A1(n646), .A2(G51), .ZN(n524) );
  XNOR2_X1 U572 ( .A(n524), .B(KEYINPUT72), .ZN(n527) );
  INV_X1 U573 ( .A(G651), .ZN(n530) );
  NOR2_X1 U574 ( .A1(G543), .A2(n530), .ZN(n525) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n525), .Z(n650) );
  NAND2_X1 U576 ( .A1(G63), .A2(n650), .ZN(n526) );
  NAND2_X1 U577 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U578 ( .A(KEYINPUT6), .B(n528), .ZN(n536) );
  NOR2_X1 U579 ( .A1(G543), .A2(G651), .ZN(n637) );
  NAND2_X1 U580 ( .A1(n637), .A2(G89), .ZN(n529) );
  XNOR2_X1 U581 ( .A(n529), .B(KEYINPUT4), .ZN(n532) );
  NOR2_X1 U582 ( .A1(n645), .A2(n530), .ZN(n635) );
  NAND2_X1 U583 ( .A1(G76), .A2(n635), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U585 ( .A(KEYINPUT71), .B(n533), .ZN(n534) );
  XNOR2_X1 U586 ( .A(KEYINPUT5), .B(n534), .ZN(n535) );
  NOR2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U588 ( .A(KEYINPUT7), .B(n537), .Z(G168) );
  XOR2_X1 U589 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U590 ( .A1(G85), .A2(n637), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G72), .A2(n635), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G60), .A2(n650), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G47), .A2(n646), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U596 ( .A1(n543), .A2(n542), .ZN(G290) );
  NAND2_X1 U597 ( .A1(G64), .A2(n650), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G52), .A2(n646), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n545), .A2(n544), .ZN(n551) );
  NAND2_X1 U600 ( .A1(n635), .A2(G77), .ZN(n546) );
  XNOR2_X1 U601 ( .A(n546), .B(KEYINPUT64), .ZN(n548) );
  NAND2_X1 U602 ( .A1(G90), .A2(n637), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(G171) );
  INV_X1 U606 ( .A(G171), .ZN(G301) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  XOR2_X2 U611 ( .A(KEYINPUT17), .B(n552), .Z(n897) );
  NAND2_X1 U612 ( .A1(G138), .A2(n897), .ZN(n554) );
  INV_X1 U613 ( .A(G2104), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G102), .A2(n560), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n559) );
  AND2_X1 U616 ( .A1(n555), .A2(G2105), .ZN(n901) );
  NAND2_X1 U617 ( .A1(G126), .A2(n901), .ZN(n557) );
  AND2_X1 U618 ( .A1(G2105), .A2(G2104), .ZN(n904) );
  NAND2_X1 U619 ( .A1(G114), .A2(n904), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U621 ( .A1(n559), .A2(n558), .ZN(G164) );
  NAND2_X1 U622 ( .A1(n897), .A2(G137), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G101), .A2(n560), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT23), .B(n561), .Z(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n685) );
  NAND2_X1 U626 ( .A1(G125), .A2(n901), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G113), .A2(n904), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n683) );
  NOR2_X1 U629 ( .A1(n685), .A2(n683), .ZN(G160) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n566) );
  XOR2_X1 U631 ( .A(n566), .B(KEYINPUT10), .Z(n836) );
  NAND2_X1 U632 ( .A1(n836), .A2(G567), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U634 ( .A1(G43), .A2(n646), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT68), .ZN(n571) );
  NAND2_X1 U636 ( .A1(G56), .A2(n650), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(KEYINPUT14), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G81), .A2(n637), .ZN(n572) );
  XOR2_X1 U640 ( .A(KEYINPUT67), .B(n572), .Z(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G68), .A2(n635), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n936) );
  NAND2_X1 U646 ( .A1(n936), .A2(G860), .ZN(G153) );
  NAND2_X1 U647 ( .A1(G66), .A2(n650), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G92), .A2(n637), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G79), .A2(n635), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G54), .A2(n646), .ZN(n581) );
  XNOR2_X1 U652 ( .A(KEYINPUT69), .B(n581), .ZN(n582) );
  NOR2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n586), .B(KEYINPUT15), .ZN(n941) );
  NOR2_X1 U656 ( .A1(n941), .A2(G868), .ZN(n587) );
  XOR2_X1 U657 ( .A(KEYINPUT70), .B(n587), .Z(n589) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G65), .A2(n650), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G53), .A2(n646), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U663 ( .A(KEYINPUT66), .B(n592), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G91), .A2(n637), .ZN(n593) );
  XNOR2_X1 U665 ( .A(KEYINPUT65), .B(n593), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n635), .A2(G78), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G299) );
  INV_X1 U669 ( .A(G868), .ZN(n663) );
  NOR2_X1 U670 ( .A1(G286), .A2(n663), .ZN(n599) );
  NOR2_X1 U671 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U673 ( .A(KEYINPUT73), .B(n600), .Z(G297) );
  INV_X1 U674 ( .A(G860), .ZN(n626) );
  NAND2_X1 U675 ( .A1(n626), .A2(G559), .ZN(n601) );
  NAND2_X1 U676 ( .A1(n601), .A2(n941), .ZN(n602) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U678 ( .A1(n941), .A2(G868), .ZN(n603) );
  XNOR2_X1 U679 ( .A(KEYINPUT74), .B(n603), .ZN(n604) );
  NOR2_X1 U680 ( .A1(G559), .A2(n604), .ZN(n605) );
  XOR2_X1 U681 ( .A(KEYINPUT75), .B(n605), .Z(n607) );
  AND2_X1 U682 ( .A1(n663), .A2(n936), .ZN(n606) );
  NOR2_X1 U683 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U684 ( .A1(n901), .A2(G123), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n608), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G111), .A2(n904), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G135), .A2(n897), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G99), .A2(n560), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n1012) );
  XOR2_X1 U692 ( .A(n1012), .B(G2096), .Z(n615) );
  NOR2_X1 U693 ( .A1(G2100), .A2(n615), .ZN(n616) );
  XOR2_X1 U694 ( .A(KEYINPUT76), .B(n616), .Z(G156) );
  NAND2_X1 U695 ( .A1(G93), .A2(n637), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G80), .A2(n635), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n650), .A2(G67), .ZN(n619) );
  XOR2_X1 U699 ( .A(KEYINPUT78), .B(n619), .Z(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n646), .A2(G55), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n665) );
  XOR2_X1 U703 ( .A(n936), .B(KEYINPUT77), .Z(n625) );
  NAND2_X1 U704 ( .A1(G559), .A2(n941), .ZN(n624) );
  XNOR2_X1 U705 ( .A(n625), .B(n624), .ZN(n661) );
  NAND2_X1 U706 ( .A1(n626), .A2(n661), .ZN(n627) );
  XOR2_X1 U707 ( .A(KEYINPUT79), .B(n627), .Z(n628) );
  XNOR2_X1 U708 ( .A(n665), .B(n628), .ZN(G145) );
  NAND2_X1 U709 ( .A1(G88), .A2(n637), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G75), .A2(n635), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G62), .A2(n650), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G50), .A2(n646), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U715 ( .A1(n634), .A2(n633), .ZN(G166) );
  INV_X1 U716 ( .A(G166), .ZN(G303) );
  NAND2_X1 U717 ( .A1(G73), .A2(n635), .ZN(n636) );
  XNOR2_X1 U718 ( .A(n636), .B(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U719 ( .A1(G86), .A2(n637), .ZN(n639) );
  NAND2_X1 U720 ( .A1(G61), .A2(n650), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G48), .A2(n646), .ZN(n640) );
  XNOR2_X1 U723 ( .A(KEYINPUT81), .B(n640), .ZN(n641) );
  NOR2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G87), .A2(n645), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G49), .A2(n646), .ZN(n648) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U730 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U732 ( .A(n653), .B(KEYINPUT80), .ZN(G288) );
  XOR2_X1 U733 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n655) );
  XOR2_X1 U734 ( .A(G303), .B(KEYINPUT19), .Z(n654) );
  XNOR2_X1 U735 ( .A(n655), .B(n654), .ZN(n658) );
  XOR2_X1 U736 ( .A(G299), .B(G290), .Z(n656) );
  XNOR2_X1 U737 ( .A(n656), .B(n665), .ZN(n657) );
  XNOR2_X1 U738 ( .A(n658), .B(n657), .ZN(n660) );
  XNOR2_X1 U739 ( .A(G305), .B(G288), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n660), .B(n659), .ZN(n866) );
  XNOR2_X1 U741 ( .A(n866), .B(n661), .ZN(n662) );
  XNOR2_X1 U742 ( .A(n662), .B(KEYINPUT84), .ZN(n664) );
  NOR2_X1 U743 ( .A1(n664), .A2(n663), .ZN(n667) );
  NOR2_X1 U744 ( .A1(G868), .A2(n665), .ZN(n666) );
  NOR2_X1 U745 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n672) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n672), .Z(n673) );
  NOR2_X1 U754 ( .A1(G218), .A2(n673), .ZN(n674) );
  NAND2_X1 U755 ( .A1(G96), .A2(n674), .ZN(n843) );
  NAND2_X1 U756 ( .A1(G2106), .A2(n843), .ZN(n678) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n675) );
  NOR2_X1 U758 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U759 ( .A1(G108), .A2(n676), .ZN(n842) );
  NAND2_X1 U760 ( .A1(G567), .A2(n842), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U762 ( .A(KEYINPUT85), .B(n679), .Z(n841) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U764 ( .A1(n841), .A2(n680), .ZN(n838) );
  NAND2_X1 U765 ( .A1(n838), .A2(G36), .ZN(G176) );
  NOR2_X1 U766 ( .A1(G1976), .A2(G288), .ZN(n776) );
  NOR2_X1 U767 ( .A1(G1971), .A2(G303), .ZN(n681) );
  NOR2_X1 U768 ( .A1(n776), .A2(n681), .ZN(n946) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n795) );
  INV_X1 U770 ( .A(G40), .ZN(n682) );
  OR2_X1 U771 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U772 ( .A(n794), .B(KEYINPUT90), .Z(n686) );
  NAND2_X1 U773 ( .A1(n795), .A2(n686), .ZN(n740) );
  NOR2_X1 U774 ( .A1(G2084), .A2(n740), .ZN(n721) );
  NAND2_X1 U775 ( .A1(n721), .A2(G8), .ZN(n734) );
  NAND2_X1 U776 ( .A1(n693), .A2(G2072), .ZN(n687) );
  XNOR2_X1 U777 ( .A(n687), .B(KEYINPUT27), .ZN(n689) );
  XOR2_X1 U778 ( .A(KEYINPUT92), .B(n715), .Z(n714) );
  AND2_X1 U779 ( .A1(n714), .A2(G1956), .ZN(n688) );
  NOR2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n707) );
  INV_X1 U781 ( .A(G299), .ZN(n706) );
  NAND2_X1 U782 ( .A1(n707), .A2(n706), .ZN(n705) );
  NAND2_X1 U783 ( .A1(G1996), .A2(n715), .ZN(n690) );
  XNOR2_X1 U784 ( .A(n690), .B(KEYINPUT26), .ZN(n692) );
  NAND2_X1 U785 ( .A1(G1341), .A2(n740), .ZN(n691) );
  NAND2_X1 U786 ( .A1(n692), .A2(n691), .ZN(n698) );
  NAND2_X1 U787 ( .A1(G1348), .A2(n740), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U789 ( .A(KEYINPUT94), .B(n696), .Z(n700) );
  NOR2_X1 U790 ( .A1(n941), .A2(n700), .ZN(n697) );
  NOR2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n936), .A2(n699), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n941), .A2(n700), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U795 ( .A(n703), .B(KEYINPUT95), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U797 ( .A(n708), .B(KEYINPUT28), .Z(n709) );
  XNOR2_X1 U798 ( .A(G2078), .B(KEYINPUT93), .ZN(n713) );
  XNOR2_X1 U799 ( .A(n713), .B(KEYINPUT25), .ZN(n986) );
  NOR2_X1 U800 ( .A1(n986), .A2(n714), .ZN(n717) );
  NOR2_X1 U801 ( .A1(n715), .A2(G1961), .ZN(n716) );
  NOR2_X1 U802 ( .A1(n717), .A2(n716), .ZN(n719) );
  NOR2_X1 U803 ( .A1(n719), .A2(G301), .ZN(n736) );
  NOR2_X1 U804 ( .A1(G1966), .A2(n778), .ZN(n720) );
  OR2_X1 U805 ( .A1(n736), .A2(n720), .ZN(n718) );
  NOR2_X1 U806 ( .A1(n738), .A2(n718), .ZN(n732) );
  INV_X1 U807 ( .A(n720), .ZN(n730) );
  AND2_X1 U808 ( .A1(G301), .A2(n719), .ZN(n728) );
  NOR2_X1 U809 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U810 ( .A(KEYINPUT97), .B(n722), .Z(n723) );
  NAND2_X1 U811 ( .A1(G8), .A2(n723), .ZN(n725) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(KEYINPUT98), .ZN(n724) );
  XNOR2_X1 U813 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U814 ( .A1(G168), .A2(n726), .ZN(n727) );
  NOR2_X1 U815 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U816 ( .A(n729), .B(KEYINPUT31), .ZN(n739) );
  AND2_X1 U817 ( .A1(n730), .A2(n739), .ZN(n731) );
  OR2_X1 U818 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U819 ( .A1(n734), .A2(n733), .ZN(n761) );
  INV_X1 U820 ( .A(G286), .ZN(n735) );
  OR2_X1 U821 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U822 ( .A1(n738), .A2(n737), .ZN(n750) );
  INV_X1 U823 ( .A(G8), .ZN(n748) );
  AND2_X1 U824 ( .A1(n739), .A2(G286), .ZN(n746) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n740), .ZN(n742) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n778), .ZN(n741) );
  NOR2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U828 ( .A1(n743), .A2(G303), .ZN(n744) );
  XNOR2_X1 U829 ( .A(KEYINPUT99), .B(n744), .ZN(n745) );
  NOR2_X1 U830 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U831 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U832 ( .A1(n750), .A2(n749), .ZN(n752) );
  XNOR2_X1 U833 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n751) );
  XNOR2_X1 U834 ( .A(n752), .B(n751), .ZN(n763) );
  NAND2_X1 U835 ( .A1(n761), .A2(n763), .ZN(n753) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n945) );
  INV_X1 U837 ( .A(n778), .ZN(n755) );
  NAND2_X1 U838 ( .A1(n945), .A2(n755), .ZN(n756) );
  NOR2_X1 U839 ( .A1(n757), .A2(n756), .ZN(n774) );
  NOR2_X1 U840 ( .A1(G1981), .A2(G305), .ZN(n758) );
  XNOR2_X1 U841 ( .A(n758), .B(KEYINPUT24), .ZN(n759) );
  XNOR2_X1 U842 ( .A(KEYINPUT91), .B(n759), .ZN(n760) );
  NOR2_X1 U843 ( .A1(n778), .A2(n760), .ZN(n766) );
  OR2_X1 U844 ( .A1(n766), .A2(n778), .ZN(n764) );
  AND2_X1 U845 ( .A1(n761), .A2(n764), .ZN(n762) );
  NAND2_X1 U846 ( .A1(n763), .A2(n762), .ZN(n772) );
  INV_X1 U847 ( .A(n764), .ZN(n770) );
  NOR2_X1 U848 ( .A1(G2090), .A2(G303), .ZN(n765) );
  NAND2_X1 U849 ( .A1(G8), .A2(n765), .ZN(n768) );
  INV_X1 U850 ( .A(n766), .ZN(n767) );
  AND2_X1 U851 ( .A1(n768), .A2(n767), .ZN(n769) );
  OR2_X1 U852 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U853 ( .A1(n772), .A2(n771), .ZN(n775) );
  OR2_X1 U854 ( .A1(KEYINPUT33), .A2(n775), .ZN(n773) );
  NOR2_X1 U855 ( .A1(n774), .A2(n773), .ZN(n819) );
  INV_X1 U856 ( .A(n775), .ZN(n782) );
  XOR2_X1 U857 ( .A(G1981), .B(G305), .Z(n933) );
  INV_X1 U858 ( .A(n933), .ZN(n780) );
  NAND2_X1 U859 ( .A1(n776), .A2(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U860 ( .A1(n778), .A2(n777), .ZN(n779) );
  OR2_X1 U861 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U862 ( .A1(n782), .A2(n781), .ZN(n817) );
  XNOR2_X1 U863 ( .A(KEYINPUT34), .B(KEYINPUT86), .ZN(n786) );
  NAND2_X1 U864 ( .A1(G140), .A2(n897), .ZN(n784) );
  NAND2_X1 U865 ( .A1(G104), .A2(n560), .ZN(n783) );
  NAND2_X1 U866 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U867 ( .A(n786), .B(n785), .ZN(n791) );
  NAND2_X1 U868 ( .A1(G128), .A2(n901), .ZN(n788) );
  NAND2_X1 U869 ( .A1(G116), .A2(n904), .ZN(n787) );
  NAND2_X1 U870 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U871 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U872 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U873 ( .A(KEYINPUT36), .B(n792), .ZN(n911) );
  XNOR2_X1 U874 ( .A(KEYINPUT37), .B(G2067), .ZN(n829) );
  NOR2_X1 U875 ( .A1(n911), .A2(n829), .ZN(n793) );
  XNOR2_X1 U876 ( .A(n793), .B(KEYINPUT87), .ZN(n1008) );
  XOR2_X1 U877 ( .A(G1986), .B(G290), .Z(n940) );
  NAND2_X1 U878 ( .A1(n1008), .A2(n940), .ZN(n796) );
  NOR2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n831) );
  NAND2_X1 U880 ( .A1(n796), .A2(n831), .ZN(n815) );
  NAND2_X1 U881 ( .A1(G131), .A2(n897), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G119), .A2(n901), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U884 ( .A1(G95), .A2(n560), .ZN(n800) );
  NAND2_X1 U885 ( .A1(G107), .A2(n904), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n884) );
  NAND2_X1 U888 ( .A1(G1991), .A2(n884), .ZN(n803) );
  XOR2_X1 U889 ( .A(KEYINPUT88), .B(n803), .Z(n813) );
  NAND2_X1 U890 ( .A1(G105), .A2(n560), .ZN(n804) );
  XNOR2_X1 U891 ( .A(n804), .B(KEYINPUT38), .ZN(n811) );
  NAND2_X1 U892 ( .A1(G141), .A2(n897), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G117), .A2(n904), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n809) );
  NAND2_X1 U895 ( .A1(G129), .A2(n901), .ZN(n807) );
  XNOR2_X1 U896 ( .A(KEYINPUT89), .B(n807), .ZN(n808) );
  NOR2_X1 U897 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n881) );
  AND2_X1 U899 ( .A1(G1996), .A2(n881), .ZN(n812) );
  NOR2_X1 U900 ( .A1(n813), .A2(n812), .ZN(n1009) );
  INV_X1 U901 ( .A(n1009), .ZN(n814) );
  NAND2_X1 U902 ( .A1(n814), .A2(n831), .ZN(n822) );
  AND2_X1 U903 ( .A1(n815), .A2(n822), .ZN(n816) );
  NAND2_X1 U904 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U905 ( .A1(n819), .A2(n818), .ZN(n821) );
  XNOR2_X1 U906 ( .A(n821), .B(n820), .ZN(n834) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n881), .ZN(n1023) );
  INV_X1 U908 ( .A(n822), .ZN(n825) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n884), .ZN(n1013) );
  NOR2_X1 U911 ( .A1(n823), .A2(n1013), .ZN(n824) );
  NOR2_X1 U912 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U913 ( .A1(n1023), .A2(n826), .ZN(n827) );
  XNOR2_X1 U914 ( .A(n827), .B(KEYINPUT39), .ZN(n828) );
  NAND2_X1 U915 ( .A1(n828), .A2(n1008), .ZN(n830) );
  NAND2_X1 U916 ( .A1(n829), .A2(n911), .ZN(n1027) );
  NAND2_X1 U917 ( .A1(n830), .A2(n1027), .ZN(n832) );
  NAND2_X1 U918 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U919 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U920 ( .A(n835), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n836), .ZN(G217) );
  INV_X1 U922 ( .A(n836), .ZN(G223) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U924 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G1), .A2(G3), .ZN(n839) );
  NAND2_X1 U926 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U927 ( .A(n840), .B(KEYINPUT106), .ZN(G188) );
  INV_X1 U928 ( .A(n841), .ZN(G319) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U934 ( .A(n844), .B(KEYINPUT107), .Z(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n846) );
  XNOR2_X1 U937 ( .A(G2678), .B(G2096), .ZN(n845) );
  XNOR2_X1 U938 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U939 ( .A(n847), .B(KEYINPUT43), .Z(n849) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2084), .ZN(n848) );
  XNOR2_X1 U941 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U942 ( .A(G2100), .B(G2090), .Z(n851) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2072), .ZN(n850) );
  XNOR2_X1 U944 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U945 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U946 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n854) );
  XNOR2_X1 U947 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1956), .B(G1961), .Z(n857) );
  XNOR2_X1 U949 ( .A(G1991), .B(G1986), .ZN(n856) );
  XNOR2_X1 U950 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U951 ( .A(G1976), .B(G1981), .Z(n859) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1971), .ZN(n858) );
  XNOR2_X1 U953 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U954 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U955 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n862) );
  XNOR2_X1 U956 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U957 ( .A(G2474), .B(n864), .ZN(n865) );
  XOR2_X1 U958 ( .A(n865), .B(G1996), .Z(G229) );
  XOR2_X1 U959 ( .A(KEYINPUT117), .B(n866), .Z(n868) );
  XNOR2_X1 U960 ( .A(n941), .B(n936), .ZN(n867) );
  XNOR2_X1 U961 ( .A(n868), .B(n867), .ZN(n870) );
  XNOR2_X1 U962 ( .A(G301), .B(G286), .ZN(n869) );
  XNOR2_X1 U963 ( .A(n870), .B(n869), .ZN(n871) );
  NOR2_X1 U964 ( .A1(G37), .A2(n871), .ZN(G397) );
  NAND2_X1 U965 ( .A1(G124), .A2(n901), .ZN(n872) );
  XNOR2_X1 U966 ( .A(n872), .B(KEYINPUT44), .ZN(n873) );
  XNOR2_X1 U967 ( .A(KEYINPUT112), .B(n873), .ZN(n876) );
  NAND2_X1 U968 ( .A1(G136), .A2(n897), .ZN(n874) );
  XOR2_X1 U969 ( .A(KEYINPUT113), .B(n874), .Z(n875) );
  NAND2_X1 U970 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U971 ( .A1(G100), .A2(n560), .ZN(n878) );
  NAND2_X1 U972 ( .A1(G112), .A2(n904), .ZN(n877) );
  NAND2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U974 ( .A1(n880), .A2(n879), .ZN(G162) );
  XNOR2_X1 U975 ( .A(n1012), .B(n881), .ZN(n883) );
  XNOR2_X1 U976 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U977 ( .A(n883), .B(n882), .ZN(n888) );
  XNOR2_X1 U978 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n886) );
  XNOR2_X1 U979 ( .A(n884), .B(G162), .ZN(n885) );
  XNOR2_X1 U980 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U981 ( .A(n888), .B(n887), .Z(n910) );
  NAND2_X1 U982 ( .A1(G139), .A2(n897), .ZN(n890) );
  NAND2_X1 U983 ( .A1(G103), .A2(n560), .ZN(n889) );
  NAND2_X1 U984 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U985 ( .A(KEYINPUT115), .B(n891), .Z(n896) );
  NAND2_X1 U986 ( .A1(G127), .A2(n901), .ZN(n893) );
  NAND2_X1 U987 ( .A1(G115), .A2(n904), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n1017) );
  NAND2_X1 U991 ( .A1(G142), .A2(n897), .ZN(n899) );
  NAND2_X1 U992 ( .A1(G106), .A2(n560), .ZN(n898) );
  NAND2_X1 U993 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n900), .B(KEYINPUT45), .ZN(n903) );
  NAND2_X1 U995 ( .A1(G130), .A2(n901), .ZN(n902) );
  NAND2_X1 U996 ( .A1(n903), .A2(n902), .ZN(n907) );
  NAND2_X1 U997 ( .A1(n904), .A2(G118), .ZN(n905) );
  XOR2_X1 U998 ( .A(KEYINPUT114), .B(n905), .Z(n906) );
  NOR2_X1 U999 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1000 ( .A(n1017), .B(n908), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n910), .B(n909), .ZN(n912) );
  XOR2_X1 U1002 ( .A(n912), .B(n911), .Z(n913) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1004 ( .A(KEYINPUT116), .B(n914), .ZN(G395) );
  XOR2_X1 U1005 ( .A(KEYINPUT103), .B(G2446), .Z(n916) );
  XNOR2_X1 U1006 ( .A(G2430), .B(G2451), .ZN(n915) );
  XNOR2_X1 U1007 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1008 ( .A(n917), .B(KEYINPUT104), .Z(n919) );
  XNOR2_X1 U1009 ( .A(G1348), .B(G1341), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(n919), .B(n918), .ZN(n923) );
  XOR2_X1 U1011 ( .A(G2435), .B(KEYINPUT105), .Z(n921) );
  XNOR2_X1 U1012 ( .A(G2438), .B(G2454), .ZN(n920) );
  XNOR2_X1 U1013 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1014 ( .A(n923), .B(n922), .Z(n925) );
  XNOR2_X1 U1015 ( .A(G2443), .B(G2427), .ZN(n924) );
  XNOR2_X1 U1016 ( .A(n925), .B(n924), .ZN(n926) );
  NAND2_X1 U1017 ( .A1(n926), .A2(G14), .ZN(n932) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n932), .ZN(n929) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n927) );
  XNOR2_X1 U1020 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1021 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1022 ( .A1(G397), .A2(G395), .ZN(n930) );
  NAND2_X1 U1023 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(n932), .ZN(G401) );
  INV_X1 U1027 ( .A(G16), .ZN(n983) );
  XOR2_X1 U1028 ( .A(n983), .B(KEYINPUT56), .Z(n957) );
  XNOR2_X1 U1029 ( .A(G168), .B(G1966), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(n935), .B(KEYINPUT57), .ZN(n955) );
  XOR2_X1 U1032 ( .A(n936), .B(G1341), .Z(n938) );
  XNOR2_X1 U1033 ( .A(G299), .B(G1956), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n944) );
  XOR2_X1 U1036 ( .A(G1348), .B(n941), .Z(n942) );
  XNOR2_X1 U1037 ( .A(KEYINPUT122), .B(n942), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n951) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n948) );
  AND2_X1 U1040 ( .A1(G303), .A2(G1971), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1042 ( .A(KEYINPUT123), .B(n949), .Z(n950) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n953) );
  XOR2_X1 U1044 ( .A(G1961), .B(G171), .Z(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1047 ( .A1(n957), .A2(n956), .ZN(n985) );
  XNOR2_X1 U1048 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n981) );
  XOR2_X1 U1049 ( .A(G1966), .B(G21), .Z(n968) );
  XNOR2_X1 U1050 ( .A(G1348), .B(KEYINPUT59), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(n958), .B(G4), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(G1956), .B(G20), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(G19), .B(G1341), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1056 ( .A(KEYINPUT125), .B(G1981), .Z(n963) );
  XNOR2_X1 U1057 ( .A(G6), .B(n963), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT60), .B(n966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(KEYINPUT124), .B(G1961), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(G5), .B(n969), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(KEYINPUT126), .B(n972), .ZN(n979) );
  XOR2_X1 U1065 ( .A(G1976), .B(G23), .Z(n974) );
  XOR2_X1 U1066 ( .A(G1971), .B(G22), .Z(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(G24), .B(G1986), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(KEYINPUT58), .B(n977), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n981), .B(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n1038) );
  INV_X1 U1075 ( .A(KEYINPUT55), .ZN(n1032) );
  XNOR2_X1 U1076 ( .A(n986), .B(G27), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(G2072), .B(G33), .ZN(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n996) );
  XOR2_X1 U1079 ( .A(G2067), .B(G26), .Z(n990) );
  XOR2_X1 U1080 ( .A(G1996), .B(G32), .Z(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n994) );
  XOR2_X1 U1082 ( .A(G1991), .B(G25), .Z(n991) );
  NAND2_X1 U1083 ( .A1(n991), .A2(G28), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(KEYINPUT120), .B(n992), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(KEYINPUT53), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(G2084), .B(G34), .Z(n998) );
  XNOR2_X1 U1089 ( .A(KEYINPUT54), .B(n998), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(G35), .B(G2090), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1093 ( .A(n1032), .B(n1003), .Z(n1005) );
  INV_X1 U1094 ( .A(G29), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(G11), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT121), .ZN(n1036) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(G160), .B(G2084), .Z(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT118), .B(n1016), .ZN(n1030) );
  XNOR2_X1 U1104 ( .A(G2072), .B(n1017), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(G164), .B(G2078), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT119), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(n1021), .B(KEYINPUT50), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(G2090), .B(G162), .Z(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(n1024), .B(KEYINPUT51), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(KEYINPUT52), .B(n1031), .ZN(n1033) );
  NAND2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1117 ( .A1(n1034), .A2(G29), .ZN(n1035) );
  NAND2_X1 U1118 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1119 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1120 ( .A(n1039), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1121 ( .A(G150), .ZN(G311) );
endmodule

