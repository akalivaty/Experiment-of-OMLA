//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(G221), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT76), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n192), .B(new_n194), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT10), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G143), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n200), .B(new_n202), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n208), .A3(new_n204), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n201), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n208), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n199), .B1(new_n211), .B2(G146), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n205), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT77), .B1(new_n214), .B2(G104), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(G104), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G101), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(G107), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n214), .A2(KEYINPUT3), .A3(G104), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(new_n214), .B2(G104), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n222), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT78), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n213), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n213), .B2(new_n227), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n197), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT65), .A2(G134), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT65), .A2(G134), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  OAI22_X1  g048(.A1(new_n232), .A2(new_n233), .B1(new_n234), .B2(G137), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(G137), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT11), .A3(G134), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(G131), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n204), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n244), .B1(new_n209), .B2(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n247), .A2(new_n248), .B1(new_n212), .B2(new_n244), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G101), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n253), .A3(G101), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n245), .B1(new_n203), .B2(new_n204), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n201), .B1(new_n200), .B2(KEYINPUT1), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n205), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n227), .A2(new_n258), .A3(KEYINPUT10), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n231), .A2(new_n242), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n242), .B1(new_n231), .B2(new_n260), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n196), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(KEYINPUT81), .B(new_n196), .C1(new_n261), .C2(new_n262), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n242), .A2(KEYINPUT79), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n229), .A2(new_n230), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n227), .A2(new_n258), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT12), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n272), .B(new_n267), .C1(new_n268), .C2(new_n269), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n231), .A2(new_n242), .A3(new_n260), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n271), .A2(new_n273), .A3(new_n274), .A4(new_n195), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n265), .A2(new_n266), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G469), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n276), .A2(new_n277), .A3(new_n188), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n261), .B2(new_n196), .ZN(new_n280));
  INV_X1    g094(.A(new_n262), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n274), .A2(KEYINPUT80), .A3(new_n195), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n196), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n285), .A3(G469), .ZN(new_n286));
  NAND2_X1  g100(.A1(G469), .A2(G902), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n191), .B1(new_n278), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n276), .A2(new_n277), .A3(new_n188), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(new_n287), .A3(new_n286), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT82), .A3(new_n191), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G475), .ZN(new_n296));
  XNOR2_X1  g110(.A(G125), .B(G140), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT16), .ZN(new_n298));
  INV_X1    g112(.A(G125), .ZN(new_n299));
  OR3_X1    g113(.A1(new_n299), .A2(KEYINPUT16), .A3(G140), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(G146), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(G146), .B1(new_n298), .B2(new_n300), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G237), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n305), .A2(new_n193), .A3(G214), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT91), .B1(new_n203), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(G143), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT91), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(new_n193), .A3(G214), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n211), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G131), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT17), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n304), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT93), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n307), .A2(new_n311), .A3(new_n317), .A4(new_n308), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n313), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT93), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n304), .B(new_n320), .C1(new_n313), .C2(new_n314), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n316), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G113), .B(G122), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(new_n217), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n297), .B(new_n204), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT18), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(new_n317), .ZN(new_n327));
  OAI221_X1 g141(.A(new_n325), .B1(new_n327), .B2(new_n312), .C1(new_n313), .C2(new_n326), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n322), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n313), .A2(new_n318), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT92), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n301), .B(KEYINPUT73), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n297), .B(KEYINPUT19), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n204), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT92), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n313), .A2(new_n335), .A3(new_n318), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n331), .A2(new_n332), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n324), .B1(new_n337), .B2(new_n328), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n296), .B(new_n188), .C1(new_n329), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT20), .ZN(new_n340));
  INV_X1    g154(.A(new_n338), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n322), .A2(new_n324), .A3(new_n328), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n296), .A4(new_n188), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n324), .B1(new_n322), .B2(new_n328), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n188), .B1(new_n329), .B2(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n340), .A2(new_n345), .B1(new_n347), .B2(G475), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT70), .B(G217), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n187), .A2(new_n193), .A3(new_n349), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n201), .A2(KEYINPUT95), .A3(G143), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT95), .B1(new_n201), .B2(G143), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n201), .B1(new_n206), .B2(new_n208), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n232), .A2(new_n233), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G116), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G122), .ZN(new_n358));
  INV_X1    g172(.A(G122), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G116), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(G107), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT94), .B1(new_n354), .B2(KEYINPUT13), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT95), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n198), .B2(G128), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n201), .A2(KEYINPUT95), .A3(G143), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT94), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT13), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n368), .B(new_n369), .C1(new_n203), .C2(new_n201), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n354), .A2(KEYINPUT13), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n363), .A2(new_n367), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n356), .B(new_n362), .C1(new_n372), .C2(G134), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT97), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n358), .B2(KEYINPUT14), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT14), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(new_n357), .A3(KEYINPUT97), .A4(G122), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n358), .A2(KEYINPUT14), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n376), .A2(new_n360), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G107), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n361), .A2(new_n214), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n232), .A2(new_n233), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n207), .A2(G143), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n386));
  OAI21_X1  g200(.A(G128), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n384), .B1(new_n387), .B2(new_n367), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT96), .B1(new_n356), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n355), .B1(new_n353), .B2(new_n354), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n384), .A3(new_n367), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI211_X1 g207(.A(KEYINPUT98), .B(new_n383), .C1(new_n389), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT98), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n393), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n381), .A2(new_n382), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n374), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT99), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n391), .B1(new_n390), .B2(new_n392), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n397), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT98), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n395), .A3(new_n397), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT99), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n374), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n350), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n350), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n373), .B1(new_n404), .B2(new_n405), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(new_n407), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n188), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT15), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(G478), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(G478), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n188), .B(new_n416), .C1(new_n409), .C2(new_n412), .ZN(new_n417));
  INV_X1    g231(.A(G952), .ZN(new_n418));
  AOI211_X1 g232(.A(G953), .B(new_n418), .C1(G234), .C2(G237), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT21), .B(G898), .Z(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI211_X1 g235(.A(new_n188), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n348), .A2(new_n415), .A3(new_n417), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT100), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n413), .B(new_n416), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT100), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n348), .A4(new_n424), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G472), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n188), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT69), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT2), .B(G113), .ZN(new_n434));
  INV_X1    g248(.A(G119), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G116), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n357), .A2(G119), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT66), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n437), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n442), .A2(new_n434), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n249), .B1(new_n240), .B2(new_n241), .ZN(new_n445));
  NAND2_X1  g259(.A1(G134), .A2(G137), .ZN(new_n446));
  OAI211_X1 g260(.A(G131), .B(new_n446), .C1(new_n355), .C2(G137), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n258), .B(new_n447), .C1(G131), .C2(new_n239), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT30), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n449), .B1(new_n445), .B2(new_n448), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n444), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT31), .ZN(new_n454));
  INV_X1    g268(.A(new_n444), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n448), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n457));
  INV_X1    g271(.A(G210), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n458), .A2(G237), .A3(G953), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n457), .B(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT26), .B(G101), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n453), .A2(new_n454), .A3(new_n456), .A4(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT68), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n456), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n445), .A2(new_n448), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT30), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n450), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n469), .B2(new_n444), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n470), .A2(KEYINPUT68), .A3(new_n454), .A4(new_n462), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n462), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT28), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n455), .B1(new_n445), .B2(new_n448), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n476), .B2(new_n456), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n456), .A2(new_n474), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n473), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n480), .A2(new_n454), .B1(new_n470), .B2(new_n462), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n433), .B1(new_n472), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT32), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n470), .A2(new_n462), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT28), .B1(new_n466), .B2(new_n475), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n462), .B1(new_n485), .B2(new_n478), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n486), .B2(KEYINPUT31), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n465), .A3(new_n471), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT32), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n433), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n462), .A3(new_n478), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n470), .A2(new_n462), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n493), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n494), .B(new_n188), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G472), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT23), .B1(new_n201), .B2(G119), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT72), .B1(new_n435), .B2(G128), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n499), .B(new_n500), .Z(new_n501));
  XNOR2_X1  g315(.A(G119), .B(G128), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT24), .B(G110), .Z(new_n503));
  OAI22_X1  g317(.A1(new_n501), .A2(G110), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n297), .A2(new_n204), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n332), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(G110), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT71), .B1(new_n503), .B2(new_n502), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n503), .A2(KEYINPUT71), .A3(new_n502), .ZN(new_n509));
  OAI221_X1 g323(.A(new_n507), .B1(new_n302), .B2(new_n303), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT22), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(G137), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n506), .A2(new_n510), .A3(new_n514), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n188), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n521));
  INV_X1    g335(.A(new_n519), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n516), .A2(new_n188), .A3(new_n517), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n349), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(G234), .B2(new_n188), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n516), .A2(new_n517), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n526), .A2(G902), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT75), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n491), .A2(new_n498), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT84), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT5), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n439), .A2(new_n440), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G113), .B1(new_n436), .B2(KEYINPUT5), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n442), .A2(KEYINPUT66), .ZN(new_n542));
  XNOR2_X1  g356(.A(G116), .B(G119), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n438), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT5), .ZN(new_n545));
  INV_X1    g359(.A(new_n540), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(KEYINPUT84), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n541), .A2(new_n443), .A3(new_n227), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n252), .A2(new_n444), .A3(new_n254), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(G110), .B(G122), .Z(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n551), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n553), .A3(new_n549), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n552), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n548), .A2(new_n553), .A3(new_n549), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n553), .B1(new_n548), .B2(new_n549), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT6), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n550), .A2(new_n558), .A3(new_n551), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT85), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n555), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n258), .A2(G125), .ZN(new_n564));
  INV_X1    g378(.A(new_n249), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(G125), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n193), .A2(G224), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n567), .B(KEYINPUT86), .Z(new_n568));
  XNOR2_X1  g382(.A(new_n566), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(KEYINPUT7), .ZN(new_n571));
  AOI211_X1 g385(.A(new_n571), .B(new_n564), .C1(G125), .C2(new_n565), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n556), .B1(KEYINPUT89), .B2(new_n572), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n572), .A2(KEYINPUT89), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n566), .A2(KEYINPUT88), .ZN(new_n575));
  INV_X1    g389(.A(new_n564), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n575), .B(new_n571), .C1(KEYINPUT88), .C2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n442), .A2(new_n538), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT87), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n443), .B1(new_n579), .B2(new_n540), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n227), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n551), .B(KEYINPUT8), .Z(new_n582));
  NAND3_X1  g396(.A1(new_n541), .A2(new_n443), .A3(new_n547), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n581), .B(new_n582), .C1(new_n583), .C2(new_n227), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n573), .A2(new_n574), .A3(new_n577), .A4(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n570), .A2(new_n188), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(G210), .B1(G237), .B2(G902), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n563), .B2(new_n569), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n587), .A3(new_n585), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(KEYINPUT90), .A3(new_n591), .ZN(new_n592));
  OR3_X1    g406(.A1(new_n586), .A2(KEYINPUT90), .A3(new_n588), .ZN(new_n593));
  OAI21_X1  g407(.A(G214), .B1(G237), .B2(G902), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n594), .B(KEYINPUT83), .Z(new_n595));
  AND3_X1   g409(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n295), .A2(new_n430), .A3(new_n536), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  NAND2_X1  g412(.A1(new_n533), .A2(new_n535), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n431), .B1(new_n488), .B2(new_n188), .ZN(new_n600));
  INV_X1    g414(.A(new_n482), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n295), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n407), .B1(new_n406), .B2(new_n374), .ZN(new_n605));
  AOI211_X1 g419(.A(KEYINPUT99), .B(new_n373), .C1(new_n404), .C2(new_n405), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n410), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  INV_X1    g422(.A(new_n412), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n410), .B1(new_n411), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n399), .A2(KEYINPUT102), .A3(new_n350), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT33), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G478), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(G902), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n604), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n618), .ZN(new_n620));
  AOI211_X1 g434(.A(KEYINPUT103), .B(new_n620), .C1(new_n610), .C2(new_n615), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n413), .A2(new_n617), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n348), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n589), .A2(KEYINPUT101), .A3(new_n591), .ZN(new_n625));
  INV_X1    g439(.A(new_n594), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n587), .B1(new_n590), .B2(new_n585), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n624), .A2(new_n424), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n603), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n340), .A2(new_n345), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n347), .A2(G475), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n339), .A2(KEYINPUT104), .A3(KEYINPUT20), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n423), .B(KEYINPUT105), .Z(new_n640));
  NOR3_X1   g454(.A1(new_n427), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n630), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n603), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT35), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  XNOR2_X1  g459(.A(new_n511), .B(KEYINPUT106), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n646), .A2(KEYINPUT36), .A3(new_n515), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n529), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n651), .A2(new_n527), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n652), .A2(new_n600), .A3(new_n601), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n295), .A2(new_n430), .A3(new_n653), .A4(new_n596), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n527), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n625), .A2(new_n629), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n415), .A2(new_n417), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n638), .A2(new_n637), .ZN(new_n660));
  INV_X1    g474(.A(new_n422), .ZN(new_n661));
  OR3_X1    g475(.A1(new_n661), .A2(KEYINPUT107), .A3(G900), .ZN(new_n662));
  INV_X1    g476(.A(new_n419), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT107), .B1(new_n661), .B2(G900), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n659), .A2(new_n660), .A3(new_n636), .A4(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n491), .A2(new_n498), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n295), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XNOR2_X1  g484(.A(new_n665), .B(KEYINPUT39), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n295), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n673), .A2(new_n348), .A3(new_n427), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n592), .A2(new_n593), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n470), .A2(new_n473), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n466), .A2(new_n475), .ZN(new_n680));
  AOI21_X1  g494(.A(G902), .B1(new_n680), .B2(new_n473), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n431), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n483), .B2(new_n490), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n672), .B2(KEYINPUT40), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n657), .A2(new_n626), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n674), .A2(new_n677), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n203), .ZN(G45));
  AOI22_X1  g501(.A1(new_n483), .A2(new_n490), .B1(G472), .B2(new_n497), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n291), .B2(new_n294), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n400), .A2(new_n408), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n412), .B1(new_n691), .B2(new_n410), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n690), .B1(new_n692), .B2(new_n608), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT103), .B1(new_n693), .B2(new_n620), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n616), .A2(new_n604), .A3(new_n618), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n623), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n348), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n696), .A2(new_n697), .A3(new_n665), .ZN(new_n698));
  INV_X1    g512(.A(new_n658), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n689), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT108), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  INV_X1    g516(.A(new_n599), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n276), .A2(new_n188), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  INV_X1    g519(.A(new_n190), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n292), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n703), .A2(new_n688), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n424), .A3(new_n630), .A4(new_n624), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT41), .B(G113), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT109), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n709), .B(new_n711), .ZN(G15));
  INV_X1    g526(.A(new_n707), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n536), .A2(new_n630), .A3(new_n641), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NOR2_X1   g529(.A1(new_n658), .A2(new_n707), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n430), .A3(new_n668), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  INV_X1    g532(.A(new_n602), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n719), .A2(new_n531), .A3(new_n707), .ZN(new_n720));
  INV_X1    g534(.A(new_n640), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT110), .B1(new_n427), .B2(new_n348), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n697), .A2(new_n659), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n720), .A2(new_n630), .A3(new_n721), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NAND3_X1  g541(.A1(new_n698), .A2(new_n716), .A3(new_n602), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n626), .B1(new_n592), .B2(new_n593), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n697), .A3(new_n696), .A4(new_n665), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n293), .A2(new_n706), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n668), .A2(new_n733), .A3(new_n599), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n730), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n688), .A2(new_n730), .A3(new_n531), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n698), .A2(new_n736), .A3(new_n733), .A4(new_n731), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  INV_X1    g553(.A(new_n666), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n731), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n734), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(G134), .Z(G36));
  INV_X1    g557(.A(new_n731), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n696), .A2(new_n348), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT112), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n348), .B(KEYINPUT113), .Z(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT43), .A3(new_n696), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n745), .A2(new_n751), .A3(new_n746), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n748), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n719), .A3(new_n657), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n744), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n283), .A2(new_n285), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT45), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(G469), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n287), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT46), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n287), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n292), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n706), .A3(new_n671), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT111), .Z(new_n768));
  NAND4_X1  g582(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n719), .A4(new_n657), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n756), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  NAND2_X1  g585(.A1(new_n766), .A2(new_n706), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n766), .A2(KEYINPUT47), .A3(new_n706), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n668), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(new_n703), .A3(new_n698), .A4(new_n731), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n688), .A2(new_n531), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n731), .A2(new_n713), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n753), .A2(new_n419), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT48), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n599), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n683), .A2(new_n419), .ZN(new_n787));
  OR3_X1    g601(.A1(new_n786), .A2(KEYINPUT117), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT117), .B1(new_n786), .B2(new_n787), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n624), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n418), .A2(G953), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n753), .A2(new_n419), .A3(new_n630), .A4(new_n720), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n779), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n783), .B(KEYINPUT48), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n792), .A2(new_n791), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(KEYINPUT118), .A3(new_n790), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n753), .A2(new_n419), .A3(new_n720), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n799), .A2(new_n626), .A3(new_n676), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n753), .A2(new_n626), .A3(new_n419), .A4(new_n720), .ZN(new_n803));
  OAI211_X1 g617(.A(KEYINPUT116), .B(new_n800), .C1(new_n803), .C2(new_n677), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n696), .A2(new_n697), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n788), .A2(new_n789), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n753), .A2(new_n419), .A3(new_n653), .A4(new_n782), .ZN(new_n808));
  INV_X1    g622(.A(new_n191), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n705), .A2(new_n809), .A3(new_n292), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n774), .A2(new_n775), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n719), .A2(new_n531), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n753), .A2(new_n419), .A3(new_n731), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n805), .A2(new_n807), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n802), .B2(new_n804), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n820), .B2(new_n807), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n798), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n683), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n706), .A2(new_n293), .A3(new_n652), .A4(new_n665), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n725), .A2(new_n630), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n700), .A2(new_n728), .A3(new_n669), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n696), .A2(new_n602), .A3(new_n697), .A4(new_n665), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n716), .A2(new_n829), .B1(new_n689), .B2(new_n667), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n700), .A4(new_n825), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n742), .B1(new_n735), .B2(new_n737), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n293), .A2(KEYINPUT82), .A3(new_n191), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT82), .B1(new_n293), .B2(new_n191), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n668), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n639), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n659), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n415), .A2(new_n417), .A3(KEYINPUT114), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n838), .A2(new_n840), .A3(new_n665), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n733), .ZN(new_n843));
  OAI22_X1  g657(.A1(new_n837), .A2(new_n842), .B1(new_n828), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n657), .A3(new_n731), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n834), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n709), .A2(new_n714), .A3(new_n726), .A4(new_n717), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n697), .B1(new_n840), .B2(new_n841), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n596), .B(new_n721), .C1(new_n624), .C2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n597), .B(new_n654), .C1(new_n850), .C2(new_n603), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n833), .A2(KEYINPUT53), .A3(new_n847), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  INV_X1    g668(.A(new_n851), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n536), .A2(new_n713), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n725), .A2(new_n630), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n713), .A2(new_n532), .A3(new_n602), .A4(new_n721), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n631), .A2(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n717), .A2(new_n714), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n855), .A2(new_n861), .A3(new_n834), .A4(new_n845), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n827), .A2(new_n832), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n854), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n853), .A2(new_n864), .A3(KEYINPUT115), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n846), .A2(new_n848), .A3(new_n851), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT53), .A4(new_n833), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(KEYINPUT54), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n853), .A2(new_n864), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT119), .B1(new_n822), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n820), .A2(new_n819), .A3(new_n807), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n874), .A2(new_n875), .B1(new_n794), .B2(new_n797), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n869), .A4(new_n871), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n418), .A2(new_n193), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n677), .A2(new_n531), .A3(new_n809), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n705), .A2(new_n292), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT49), .Z(new_n883));
  AND3_X1   g697(.A1(new_n883), .A2(new_n595), .A3(new_n683), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n881), .A2(new_n696), .A3(new_n749), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n193), .A2(G952), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n563), .B(new_n569), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  XOR2_X1   g703(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n890));
  AOI21_X1  g704(.A(new_n188), .B1(new_n853), .B2(new_n864), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n889), .B(new_n890), .C1(new_n891), .C2(G210), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n853), .A2(new_n864), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(G902), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n895), .B2(new_n458), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n891), .A2(KEYINPUT120), .A3(G210), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n887), .B(new_n892), .C1(new_n899), .C2(new_n889), .ZN(G51));
  INV_X1    g714(.A(new_n887), .ZN(new_n901));
  INV_X1    g715(.A(new_n276), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n287), .A2(KEYINPUT57), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n866), .B2(new_n833), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n862), .A2(new_n863), .A3(new_n854), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT54), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(new_n907), .B2(new_n871), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n287), .A2(KEYINPUT57), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n902), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n895), .A2(new_n761), .ZN(new_n911));
  OAI211_X1 g725(.A(KEYINPUT122), .B(new_n901), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n853), .A2(new_n870), .A3(new_n864), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n870), .B1(new_n853), .B2(new_n864), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n909), .B(new_n903), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n911), .B1(new_n916), .B2(new_n276), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n913), .B1(new_n917), .B2(new_n887), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  INV_X1    g734(.A(new_n343), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n887), .ZN(G60));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n869), .B2(new_n871), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n901), .B1(new_n927), .B2(new_n616), .ZN(new_n928));
  INV_X1    g742(.A(new_n926), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n616), .B(new_n929), .C1(new_n914), .C2(new_n915), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(G63));
  XOR2_X1   g748(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n935), .B(new_n936), .Z(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n853), .B2(new_n864), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n649), .A2(new_n650), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n887), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n528), .B2(new_n938), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT61), .Z(G66));
  INV_X1    g757(.A(G224), .ZN(new_n944));
  OAI21_X1  g758(.A(G953), .B1(new_n421), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n852), .B2(G953), .ZN(new_n946));
  INV_X1    g760(.A(new_n563), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(G898), .B2(new_n193), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G69));
  XOR2_X1   g763(.A(new_n469), .B(new_n333), .Z(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(G900), .B2(G953), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n768), .A2(new_n630), .A3(new_n725), .A4(new_n780), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n952), .A2(new_n834), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n830), .A2(new_n700), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n770), .A2(KEYINPUT126), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT126), .B1(new_n770), .B2(new_n954), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n777), .B(new_n953), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n951), .B1(new_n957), .B2(G953), .ZN(new_n958));
  XOR2_X1   g772(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n686), .A2(new_n954), .A3(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n960), .A2(new_n777), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n536), .B1(new_n624), .B2(new_n849), .ZN(new_n962));
  OR3_X1    g776(.A1(new_n962), .A2(new_n672), .A3(new_n744), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n686), .A2(new_n954), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(KEYINPUT62), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n961), .A2(new_n770), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n193), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n950), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n958), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n971), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n958), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(new_n470), .A2(new_n473), .ZN(new_n976));
  INV_X1    g790(.A(new_n852), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n957), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  AOI21_X1  g794(.A(new_n976), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n967), .B2(new_n977), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n678), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n679), .A2(new_n980), .A3(new_n976), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT127), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n865), .A2(new_n868), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n901), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n981), .A2(new_n987), .ZN(G57));
endmodule


