//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967;
  NAND2_X1  g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G71gat), .B(G78gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT96), .B(G57gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G64gat), .ZN(new_n207));
  INV_X1    g006(.A(G64gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G57gat), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n207), .A2(KEYINPUT97), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT97), .B1(new_n207), .B2(new_n209), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n204), .B(new_n205), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n205), .B(KEYINPUT95), .ZN(new_n213));
  INV_X1    g012(.A(new_n209), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n208), .A2(G57gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n204), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G231gat), .A2(G233gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G127gat), .B(G155gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n218), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT98), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT98), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n218), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(KEYINPUT21), .A3(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G15gat), .B(G22gat), .Z(new_n232));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(G1gat), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT94), .Z(new_n236));
  INV_X1    g035(.A(G8gat), .ZN(new_n237));
  INV_X1    g036(.A(G1gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(KEYINPUT93), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n235), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G8gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n231), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n226), .B(new_n246), .Z(new_n247));
  XOR2_X1   g046(.A(G183gat), .B(G211gat), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n226), .B(new_n246), .ZN(new_n250));
  INV_X1    g049(.A(new_n248), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  OR3_X1    g052(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT91), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT88), .B(G29gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G36gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT92), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT15), .ZN(new_n262));
  XOR2_X1   g061(.A(KEYINPUT89), .B(G43gat), .Z(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G50gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT90), .B(G50gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(G43gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n254), .A2(KEYINPUT91), .A3(new_n255), .ZN(new_n268));
  XNOR2_X1  g067(.A(G43gat), .B(G50gat), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n258), .A2(KEYINPUT92), .B1(KEYINPUT15), .B2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n261), .A2(new_n267), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT87), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n254), .B1(new_n272), .B2(new_n255), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n255), .A2(new_n272), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n258), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT15), .A3(new_n269), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT17), .ZN(new_n278));
  NAND2_X1  g077(.A1(G85gat), .A2(G92gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT7), .ZN(new_n280));
  NAND2_X1  g079(.A1(G99gat), .A2(G106gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT8), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n280), .B(new_n282), .C1(G85gat), .C2(G92gat), .ZN(new_n283));
  XOR2_X1   g082(.A(G99gat), .B(G106gat), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  AND2_X1   g086(.A1(G232gat), .A2(G233gat), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n277), .A2(new_n287), .B1(KEYINPUT41), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G190gat), .B(G218gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT99), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT100), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT100), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n295), .A3(new_n292), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n290), .A2(new_n292), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n288), .A2(KEYINPUT41), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n299), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n294), .A2(new_n297), .A3(new_n301), .A4(new_n296), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G134gat), .B(G162gat), .Z(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n306), .B1(new_n300), .B2(new_n302), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n253), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G230gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n284), .A2(KEYINPUT102), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n283), .B(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n227), .A2(new_n313), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n218), .A2(KEYINPUT101), .A3(new_n285), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT101), .B1(new_n218), .B2(new_n285), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n311), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT103), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n228), .A2(KEYINPUT10), .A3(new_n230), .A4(new_n287), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n310), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT104), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(KEYINPUT104), .B(new_n310), .C1(new_n320), .C2(new_n321), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n315), .A2(new_n316), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n227), .B2(new_n313), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(new_n310), .ZN(new_n329));
  XNOR2_X1  g128(.A(G120gat), .B(G148gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT105), .ZN(new_n331));
  XOR2_X1   g130(.A(G176gat), .B(G204gat), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n319), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n336), .A2(new_n310), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n333), .B1(new_n337), .B2(new_n329), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT106), .B1(new_n309), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n278), .A2(new_n245), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n244), .A2(new_n277), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G229gat), .A2(G233gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT18), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(KEYINPUT18), .A3(new_n344), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n244), .B(new_n277), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n344), .B(KEYINPUT13), .Z(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G113gat), .B(G141gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT11), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(G197gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT12), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n352), .B(new_n358), .Z(new_n359));
  INV_X1    g158(.A(KEYINPUT106), .ZN(new_n360));
  INV_X1    g159(.A(new_n339), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n253), .A2(new_n360), .A3(new_n308), .A4(new_n361), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n340), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365));
  INV_X1    g164(.A(G211gat), .ZN(new_n366));
  INV_X1    g165(.A(G218gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n364), .A3(new_n368), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n376), .B(KEYINPUT71), .Z(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT27), .B(G183gat), .ZN(new_n378));
  INV_X1    g177(.A(G190gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(KEYINPUT28), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G183gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT27), .B1(new_n381), .B2(KEYINPUT66), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT66), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(G183gat), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n382), .A2(new_n385), .A3(new_n379), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n380), .B1(new_n386), .B2(KEYINPUT28), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT67), .ZN(new_n388));
  NOR3_X1   g187(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT26), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n389), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n388), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n390), .B1(new_n393), .B2(new_n392), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT67), .B(new_n396), .C1(new_n399), .C2(new_n389), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n387), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n390), .A2(KEYINPUT23), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT23), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n404), .B1(G169gat), .B2(G176gat), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n403), .B1(new_n405), .B2(new_n390), .ZN(new_n406));
  AND3_X1   g205(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n396), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(KEYINPUT64), .B(new_n402), .C1(new_n406), .C2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n396), .ZN(new_n412));
  OAI211_X1 g211(.A(G183gat), .B(G190gat), .C1(KEYINPUT65), .C2(KEYINPUT24), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n412), .B(new_n413), .C1(G183gat), .C2(G190gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n392), .A2(KEYINPUT23), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n391), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n414), .A2(KEYINPUT25), .A3(new_n403), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(new_n396), .ZN(new_n419));
  NAND3_X1  g218(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(new_n403), .A3(new_n416), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT64), .B1(new_n422), .B2(new_n402), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n401), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n377), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n377), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n402), .B1(new_n406), .B2(new_n409), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n410), .A3(new_n417), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n431), .B2(new_n401), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n375), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT72), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(new_n375), .C1(new_n426), .C2(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT73), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n426), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n432), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n426), .A2(new_n438), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n374), .A4(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n437), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT75), .B(KEYINPUT30), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n446), .B1(new_n437), .B2(new_n442), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n437), .A2(new_n442), .A3(KEYINPUT30), .A4(new_n446), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454));
  XOR2_X1   g253(.A(G155gat), .B(G162gat), .Z(new_n455));
  XNOR2_X1  g254(.A(G141gat), .B(G148gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(G148gat), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(G141gat), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT77), .B1(new_n459), .B2(G141gat), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT2), .ZN(new_n465));
  INV_X1    g264(.A(G155gat), .ZN(new_n466));
  INV_X1    g265(.A(G162gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G155gat), .A2(G162gat), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n458), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G127gat), .B(G134gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT1), .ZN(new_n473));
  INV_X1    g272(.A(G113gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(G120gat), .ZN(new_n475));
  INV_X1    g274(.A(G120gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(G113gat), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n472), .B(new_n473), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G113gat), .B(G120gat), .ZN(new_n479));
  INV_X1    g278(.A(G134gat), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n480), .A2(G127gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(G127gat), .ZN(new_n482));
  OAI22_X1  g281(.A1(new_n479), .A2(KEYINPUT1), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n454), .B1(new_n471), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n462), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n486), .A2(new_n460), .B1(new_n469), .B2(new_n468), .ZN(new_n487));
  XNOR2_X1  g286(.A(G155gat), .B(G162gat), .ZN(new_n488));
  INV_X1    g287(.A(G141gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G148gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n465), .A2(KEYINPUT76), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT76), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT2), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n488), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n478), .A2(new_n483), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n485), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT78), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n487), .B2(new_n496), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n458), .B(KEYINPUT78), .C1(new_n464), .C2(new_n470), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT3), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT3), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n498), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n500), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n507), .A2(KEYINPUT39), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G1gat), .B(G29gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT0), .ZN(new_n511));
  XNOR2_X1  g310(.A(G57gat), .B(G85gat), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n511), .B(new_n512), .Z(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n502), .A2(new_n503), .A3(new_n484), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n498), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n508), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT39), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(KEYINPUT85), .B(KEYINPUT39), .C1(new_n518), .C2(new_n519), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n522), .B(new_n523), .C1(new_n508), .C2(new_n507), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n515), .A2(KEYINPUT40), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n485), .A2(new_n499), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n504), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n526), .A2(new_n508), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT79), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n518), .B2(new_n519), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT5), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n518), .A2(new_n529), .A3(new_n519), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n526), .A2(new_n527), .A3(new_n508), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n535), .A3(new_n514), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n525), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT40), .B1(new_n515), .B2(new_n524), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n453), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n497), .A2(new_n505), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n374), .B1(new_n541), .B2(new_n425), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT29), .B1(new_n372), .B2(new_n373), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n471), .B1(new_n543), .B2(KEYINPUT3), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G228gat), .ZN(new_n546));
  INV_X1    g345(.A(G233gat), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n542), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n541), .A2(new_n425), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n375), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n546), .A2(new_n547), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n502), .B(new_n503), .C1(new_n543), .C2(KEYINPUT3), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G22gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n548), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n548), .B2(new_n553), .ZN(new_n557));
  XNOR2_X1  g356(.A(G78gat), .B(G106gat), .ZN(new_n558));
  INV_X1    g357(.A(G50gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n548), .A2(new_n553), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G22gat), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n564), .B2(new_n555), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT83), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n561), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n560), .B1(new_n556), .B2(new_n557), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n564), .A2(new_n555), .A3(new_n562), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n540), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT5), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n518), .A2(new_n519), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT79), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n575), .B1(new_n577), .B2(new_n534), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n507), .A2(new_n508), .B1(new_n532), .B2(KEYINPUT5), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n513), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n536), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n531), .A2(new_n535), .A3(new_n514), .A4(new_n581), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n447), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT38), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n437), .A2(new_n442), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n586), .B1(new_n587), .B2(KEYINPUT37), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n588), .B(new_n445), .C1(KEYINPUT37), .C2(new_n587), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n439), .A2(new_n440), .A3(new_n375), .A4(new_n441), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n374), .B1(new_n426), .B2(new_n432), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(KEYINPUT37), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n445), .B(new_n592), .C1(new_n587), .C2(KEYINPUT37), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n586), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n585), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n574), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT74), .ZN(new_n598));
  INV_X1    g397(.A(new_n452), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n450), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n451), .A2(KEYINPUT74), .A3(new_n452), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n583), .A2(new_n584), .B1(new_n447), .B2(new_n448), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT81), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT81), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n573), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT70), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT68), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n431), .A2(new_n612), .A3(new_n498), .A4(new_n401), .ZN(new_n613));
  INV_X1    g412(.A(G227gat), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT68), .B1(new_n424), .B2(new_n484), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n401), .B(new_n498), .C1(new_n418), .C2(new_n423), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI221_X1 g416(.A(new_n613), .B1(new_n614), .B2(new_n547), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT34), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT32), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n613), .B1(new_n615), .B2(new_n617), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n614), .A2(new_n547), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT33), .B1(new_n621), .B2(new_n622), .ZN(new_n624));
  XOR2_X1   g423(.A(G15gat), .B(G43gat), .Z(new_n625));
  XNOR2_X1  g424(.A(G71gat), .B(G99gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  AOI221_X4 g428(.A(new_n620), .B1(KEYINPUT33), .B2(new_n627), .C1(new_n621), .C2(new_n622), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n611), .B(new_n619), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n623), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n621), .A2(new_n622), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n635), .A3(new_n627), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT34), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n618), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n630), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n631), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n639), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n611), .B1(new_n642), .B2(new_n619), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n610), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n619), .B1(new_n629), .B2(new_n630), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT69), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT69), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n642), .A2(new_n647), .A3(new_n619), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n646), .A2(new_n648), .A3(KEYINPUT36), .A4(new_n640), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT84), .B1(new_n609), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n573), .B1(new_n604), .B2(new_n606), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n644), .A2(new_n649), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT84), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n597), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  AND4_X1   g455(.A1(new_n648), .A2(new_n646), .A3(new_n573), .A4(new_n640), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n604), .A3(new_n606), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT35), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT86), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n583), .A2(new_n584), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n453), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n599), .A2(new_n450), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n583), .A2(new_n584), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n663), .A2(KEYINPUT86), .A3(new_n664), .A4(new_n449), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n569), .A2(new_n572), .A3(KEYINPUT35), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n645), .A2(KEYINPUT70), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n667), .A2(new_n668), .A3(new_n640), .A4(new_n631), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n659), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n363), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n661), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  INV_X1    g476(.A(new_n453), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT107), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n233), .ZN(new_n681));
  OR3_X1    g480(.A1(new_n674), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(G8gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(G8gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n679), .B1(new_n674), .B2(new_n678), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(G15gat), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n641), .A2(new_n643), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n675), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n675), .A2(new_n653), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n691), .B2(new_n687), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n608), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  AOI21_X1  g494(.A(new_n308), .B1(new_n656), .B2(new_n672), .ZN(new_n696));
  INV_X1    g495(.A(new_n359), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n253), .A2(new_n697), .A3(new_n339), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n699), .A2(new_n664), .A3(new_n257), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT45), .Z(new_n701));
  INV_X1    g500(.A(new_n698), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  INV_X1    g502(.A(new_n308), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n652), .A2(new_n653), .A3(new_n596), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n670), .B1(new_n658), .B2(KEYINPUT35), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT108), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n609), .A2(new_n597), .A3(new_n650), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n672), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n703), .A4(new_n704), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n609), .A2(KEYINPUT84), .A3(new_n650), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n654), .B1(new_n652), .B2(new_n653), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n706), .B1(new_n716), .B2(new_n597), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT44), .B1(new_n717), .B2(new_n308), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n702), .B1(new_n713), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n257), .B1(new_n720), .B2(new_n664), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n701), .A2(new_n721), .ZN(G1328gat));
  NOR3_X1   g521(.A1(new_n699), .A2(G36gat), .A3(new_n678), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT46), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n720), .B2(new_n678), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1329gat));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n703), .B1(new_n673), .B2(new_n704), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n708), .A2(new_n712), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n653), .B(new_n698), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n263), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(KEYINPUT109), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n699), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n688), .A2(new_n263), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT109), .B1(new_n730), .B2(new_n731), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n727), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n719), .B2(new_n653), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n708), .B(new_n712), .C1(new_n696), .C2(new_n703), .ZN(new_n743));
  AND4_X1   g542(.A1(new_n741), .A2(new_n743), .A3(new_n653), .A4(new_n698), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n731), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n736), .A2(KEYINPUT47), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n740), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n730), .A2(KEYINPUT110), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n743), .A2(new_n741), .A3(new_n653), .A4(new_n698), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n263), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(KEYINPUT111), .A3(new_n746), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n739), .B1(new_n748), .B2(new_n752), .ZN(G1330gat));
  OAI21_X1  g552(.A(new_n265), .B1(new_n699), .B2(new_n573), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n573), .A2(new_n265), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n720), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g556(.A1(new_n309), .A2(new_n359), .A3(new_n361), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n758), .A2(new_n710), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n661), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(new_n206), .Z(G1332gat));
  AOI21_X1  g560(.A(new_n678), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n763), .B(new_n764), .Z(G1333gat));
  NAND2_X1  g564(.A1(new_n759), .A2(new_n653), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n641), .A2(new_n643), .A3(G71gat), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n766), .A2(G71gat), .B1(new_n759), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n759), .A2(new_n608), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g570(.A1(new_n253), .A2(new_n359), .A3(new_n361), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n743), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n774), .A2(G85gat), .A3(new_n661), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n253), .A2(new_n359), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n710), .A2(new_n776), .A3(new_n704), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n339), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n661), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n775), .A2(new_n783), .ZN(G1336gat));
  NAND3_X1  g583(.A1(new_n743), .A2(new_n453), .A3(new_n772), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n781), .A2(G92gat), .A3(new_n678), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n788));
  OR3_X1    g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n785), .A2(new_n790), .A3(G92gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n785), .B2(G92gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n791), .A2(new_n792), .A3(new_n787), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(G1337gat));
  AND3_X1   g594(.A1(new_n774), .A2(G99gat), .A3(new_n653), .ZN(new_n796));
  AOI21_X1  g595(.A(G99gat), .B1(new_n782), .B2(new_n688), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(G1338gat));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  AOI21_X1  g598(.A(G106gat), .B1(new_n782), .B2(new_n608), .ZN(new_n800));
  INV_X1    g599(.A(G106gat), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n773), .A2(new_n801), .A3(new_n573), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT53), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n799), .B(new_n805), .C1(new_n800), .C2(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1339gat));
  INV_X1    g606(.A(new_n253), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT54), .B1(new_n336), .B2(new_n310), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n324), .B2(new_n325), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n336), .A2(new_n811), .A3(new_n310), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n812), .A2(KEYINPUT115), .A3(new_n333), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT115), .B1(new_n812), .B2(new_n333), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n816), .A2(KEYINPUT55), .B1(new_n326), .B2(new_n334), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n810), .B2(new_n815), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT116), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n818), .C1(new_n810), .C2(new_n815), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n817), .A2(new_n359), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n347), .A2(new_n348), .A3(new_n351), .A4(new_n358), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n343), .A2(new_n344), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n349), .A2(new_n350), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n357), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n339), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n704), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n817), .A2(new_n822), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n828), .B1(new_n305), .B2(new_n307), .ZN(new_n832));
  INV_X1    g631(.A(new_n820), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n808), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n253), .A2(new_n697), .A3(new_n308), .A4(new_n361), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n453), .A2(new_n664), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n657), .ZN(new_n841));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n359), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n608), .A2(new_n641), .A3(new_n643), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(new_n474), .A3(new_n697), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n842), .A2(new_n845), .ZN(G1340gat));
  AOI21_X1  g645(.A(G120gat), .B1(new_n841), .B2(new_n339), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n844), .A2(new_n476), .A3(new_n361), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(G1341gat));
  AOI21_X1  g648(.A(G127gat), .B1(new_n841), .B2(new_n253), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n840), .A2(G127gat), .A3(new_n253), .A4(new_n843), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(G1342gat));
  OAI21_X1  g654(.A(G134gat), .B1(new_n844), .B2(new_n308), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT118), .Z(new_n857));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n480), .A3(new_n657), .A4(new_n704), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT56), .Z(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1343gat));
  AND2_X1   g659(.A1(new_n650), .A2(new_n838), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n837), .B2(new_n608), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n573), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n829), .B(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n817), .A2(new_n359), .A3(new_n819), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n704), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n808), .B1(new_n869), .B2(new_n834), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n865), .B1(new_n870), .B2(new_n836), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n359), .B(new_n861), .C1(new_n862), .C2(new_n871), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(KEYINPUT121), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(KEYINPUT121), .ZN(new_n874));
  OAI21_X1  g673(.A(G141gat), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n653), .A2(new_n573), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n839), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n489), .A3(new_n359), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n872), .A2(new_n883), .A3(G141gat), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n879), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n872), .B2(G141gat), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT58), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n882), .A2(new_n887), .ZN(G1344gat));
  NOR3_X1   g687(.A1(new_n453), .A2(G148gat), .A3(new_n664), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n837), .A2(new_n339), .A3(new_n876), .A4(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n340), .A2(new_n697), .A3(new_n362), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n867), .A2(new_n868), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n308), .ZN(new_n894));
  INV_X1    g693(.A(new_n834), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n253), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n863), .B(new_n608), .C1(new_n892), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n837), .A2(new_n608), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT57), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n339), .A3(new_n861), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n891), .B1(new_n901), .B2(G148gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n861), .B1(new_n862), .B2(new_n871), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n361), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(KEYINPUT59), .A3(new_n459), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n890), .B1(new_n902), .B2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(G155gat), .B1(new_n903), .B2(new_n808), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n878), .A2(new_n466), .A3(new_n253), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1346gat));
  NAND4_X1  g708(.A1(new_n840), .A2(new_n467), .A3(new_n704), .A4(new_n876), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT123), .ZN(new_n911));
  OAI21_X1  g710(.A(G162gat), .B1(new_n903), .B2(new_n308), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n678), .A2(new_n661), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n837), .A2(new_n843), .A3(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(new_n355), .A3(new_n697), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n661), .B1(new_n835), .B2(new_n836), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n657), .A2(new_n453), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n918), .B(KEYINPUT124), .Z(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n359), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n916), .B1(new_n922), .B2(new_n355), .ZN(G1348gat));
  OAI21_X1  g722(.A(G176gat), .B1(new_n915), .B2(new_n361), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n361), .A2(G176gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n920), .B2(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(G183gat), .B1(new_n915), .B2(new_n808), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n253), .A2(new_n378), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n920), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n921), .A2(new_n379), .A3(new_n704), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n837), .A2(new_n704), .A3(new_n843), .A4(new_n914), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G190gat), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n932), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n935), .A2(new_n937), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n931), .B1(new_n942), .B2(new_n943), .ZN(G1351gat));
  NAND4_X1  g743(.A1(new_n897), .A2(new_n899), .A3(new_n650), .A4(new_n914), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n359), .A2(G197gat), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n877), .A2(new_n678), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n917), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n697), .ZN(new_n949));
  OAI22_X1  g748(.A1(new_n945), .A2(new_n946), .B1(G197gat), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n900), .A2(new_n339), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n650), .A2(new_n914), .ZN(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n948), .A2(G204gat), .A3(new_n361), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1353gat));
  NAND4_X1  g756(.A1(new_n917), .A2(new_n366), .A3(new_n253), .A4(new_n947), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n945), .A2(new_n808), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n960));
  OAI211_X1 g759(.A(KEYINPUT63), .B(G211gat), .C1(new_n945), .C2(new_n808), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n960), .B2(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(new_n367), .B1(new_n948), .B2(new_n308), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n704), .A2(G218gat), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n945), .B2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(G1355gat));
endmodule


