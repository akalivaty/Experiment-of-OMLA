//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g0015(.A(KEYINPUT65), .B(G244), .Z(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G77), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n209), .B(new_n215), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G1), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n243), .A2(G13), .A3(G20), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT70), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g0046(.A1(new_n243), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n247));
  AND2_X1   g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT69), .B1(new_n206), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT69), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n251), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n212), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n213), .A2(G1), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(new_n257), .B1(new_n248), .B2(new_n255), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT66), .ZN(new_n259));
  AND2_X1   g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  OAI21_X1  g0060(.A(G274), .B1(new_n260), .B2(new_n212), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n243), .B1(G41), .B2(G45), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n262), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(KEYINPUT66), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(G223), .A2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G226), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G1698), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n271), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G87), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n260), .A2(new_n212), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT78), .B(G190), .Z(new_n281));
  NAND3_X1  g0081(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n282), .A2(G232), .A3(new_n262), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AND4_X1   g0084(.A1(new_n270), .A2(new_n280), .A3(new_n281), .A4(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G200), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n278), .B2(new_n279), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n270), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT7), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n249), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n290), .B1(new_n294), .B2(G20), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n293), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT77), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n274), .A2(new_n275), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT77), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT7), .A4(new_n213), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n295), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G68), .ZN(new_n302));
  INV_X1    g0102(.A(G58), .ZN(new_n303));
  INV_X1    g0103(.A(G68), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(G20), .B1(new_n305), .B2(new_n201), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G20), .A2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G159), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT16), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n253), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT67), .B1(new_n274), .B2(new_n275), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT67), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n292), .A2(new_n315), .A3(new_n293), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT7), .B1(new_n317), .B2(new_n213), .ZN(new_n318));
  INV_X1    g0118(.A(new_n296), .ZN(new_n319));
  OAI21_X1  g0119(.A(G68), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n309), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT16), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n258), .B(new_n289), .C1(new_n313), .C2(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT17), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT18), .ZN(new_n325));
  INV_X1    g0125(.A(new_n258), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT67), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n315), .B1(new_n292), .B2(new_n293), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n213), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n319), .B1(new_n329), .B2(new_n290), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n321), .B1(new_n330), .B2(new_n304), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n310), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n250), .A2(new_n212), .A3(new_n252), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n302), .B2(new_n311), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n326), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n287), .A2(G179), .A3(new_n270), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n287), .B2(new_n270), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n325), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n258), .B1(new_n313), .B2(new_n322), .ZN(new_n341));
  INV_X1    g0141(.A(new_n339), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT18), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n279), .A2(new_n268), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n216), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n270), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n270), .A2(KEYINPUT71), .A3(new_n346), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT68), .ZN(new_n352));
  INV_X1    g0152(.A(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n317), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT68), .A4(G1698), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G238), .A3(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n314), .A2(new_n316), .A3(new_n353), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(G232), .B1(G107), .B2(new_n317), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n282), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(G200), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n255), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n307), .B1(new_n217), .B2(G20), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(KEYINPUT72), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n213), .A2(G33), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n362), .B2(KEYINPUT72), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n333), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n256), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n254), .A2(G77), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n217), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT73), .B1(new_n248), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n246), .A2(new_n247), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n373), .A2(new_n374), .A3(new_n217), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n370), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT74), .B1(new_n360), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n360), .A2(KEYINPUT74), .A3(new_n377), .ZN(new_n379));
  INV_X1    g0179(.A(new_n359), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n349), .A2(new_n350), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(G190), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n324), .B(new_n344), .C1(new_n378), .C2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n354), .A2(G223), .A3(new_n355), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n357), .A2(G222), .B1(new_n217), .B2(new_n317), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n282), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n345), .A2(G226), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n270), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n337), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n203), .A2(G20), .ZN(new_n391));
  INV_X1    g0191(.A(G150), .ZN(new_n392));
  INV_X1    g0192(.A(new_n307), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n391), .B1(new_n392), .B2(new_n393), .C1(new_n255), .C2(new_n365), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n253), .B1(new_n202), .B2(new_n248), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n254), .A2(G50), .A3(new_n369), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n387), .A2(G179), .A3(new_n389), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n389), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n385), .A2(new_n386), .ZN(new_n402));
  OAI211_X1 g0202(.A(G190), .B(new_n401), .C1(new_n402), .C2(new_n282), .ZN(new_n403));
  OAI21_X1  g0203(.A(G200), .B1(new_n387), .B2(new_n389), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT9), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT9), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n403), .A2(new_n404), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT10), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT75), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n409), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n408), .A2(new_n411), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n400), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n307), .A2(G50), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT76), .ZN(new_n416));
  INV_X1    g0216(.A(G77), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n365), .A2(new_n417), .B1(new_n213), .B2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n253), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT11), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n254), .A2(G68), .A3(new_n369), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT12), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n373), .B2(G68), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n248), .A2(KEYINPUT12), .A3(new_n304), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n419), .C2(new_n420), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n345), .A2(G238), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n270), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G226), .A2(G1698), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n228), .B2(G1698), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n314), .A2(new_n433), .A3(new_n316), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n282), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n435), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n279), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT13), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n263), .A2(new_n269), .B1(new_n345), .B2(G238), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(G169), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n437), .A2(new_n442), .A3(G179), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n443), .B2(G169), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n429), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n431), .A2(KEYINPUT13), .A3(new_n436), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n451));
  OAI21_X1  g0251(.A(G200), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n437), .A2(new_n442), .A3(G190), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n428), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G179), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n380), .A2(new_n381), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n377), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n337), .B1(new_n351), .B2(new_n359), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n449), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n384), .A2(new_n414), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G107), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n330), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  INV_X1    g0264(.A(G97), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n464), .A2(new_n465), .A3(G107), .ZN(new_n466));
  XNOR2_X1  g0266(.A(G97), .B(G107), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n468), .A2(new_n213), .B1(new_n417), .B2(new_n393), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n253), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n243), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n333), .A2(new_n373), .A3(new_n471), .ZN(new_n472));
  MUX2_X1   g0272(.A(new_n373), .B(new_n472), .S(G97), .Z(new_n473));
  INV_X1    g0273(.A(G283), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n249), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(new_n353), .C1(new_n274), .C2(new_n275), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n353), .A2(G244), .ZN(new_n479));
  INV_X1    g0279(.A(G250), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n479), .A2(new_n477), .B1(new_n480), .B2(new_n353), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n314), .A3(new_n316), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n282), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  NAND2_X1  g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(G257), .A3(new_n282), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT5), .B(G41), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n267), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n483), .A2(new_n493), .A3(G190), .ZN(new_n494));
  INV_X1    g0294(.A(new_n482), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n479), .B1(new_n292), .B2(new_n293), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n496), .A2(KEYINPUT4), .B1(new_n249), .B2(new_n474), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n279), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n493), .ZN(new_n499));
  AOI21_X1  g0299(.A(G200), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n470), .B(new_n473), .C1(new_n494), .C2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(G169), .B1(new_n498), .B2(new_n499), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n483), .A2(new_n493), .A3(G179), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(G20), .B1(new_n314), .B2(new_n316), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n296), .B1(new_n505), .B2(KEYINPUT7), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n469), .B1(new_n506), .B2(G107), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n473), .B1(new_n507), .B2(new_n333), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT19), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n213), .B1(new_n435), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n465), .A3(new_n462), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n213), .B(G68), .C1(new_n274), .C2(new_n275), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n510), .B1(new_n365), .B2(new_n465), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n253), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n248), .A2(new_n364), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n472), .C2(new_n364), .ZN(new_n520));
  OR2_X1    g0320(.A1(G238), .A2(G1698), .ZN(new_n521));
  INV_X1    g0321(.A(G244), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G1698), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n523), .C1(new_n274), .C2(new_n275), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G116), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n282), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n480), .B1(new_n243), .B2(G45), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n282), .ZN(new_n528));
  INV_X1    g0328(.A(new_n485), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n261), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n455), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n520), .B(new_n532), .C1(G169), .C2(new_n531), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n267), .A2(new_n485), .B1(new_n282), .B2(new_n527), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G238), .A2(G1698), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n522), .B2(G1698), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(new_n294), .B1(G33), .B2(G116), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n534), .B1(new_n537), .B2(new_n282), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n531), .A2(G190), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n517), .A2(new_n253), .B1(new_n248), .B2(new_n364), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n333), .A2(G87), .A3(new_n373), .A4(new_n471), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n539), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n533), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n501), .A2(new_n509), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n472), .A2(G116), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n248), .A2(G116), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(G20), .B1(G33), .B2(G283), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n249), .A2(G97), .ZN(new_n551));
  INV_X1    g0351(.A(G116), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n550), .A2(new_n551), .B1(G20), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n253), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n253), .A2(KEYINPUT20), .A3(new_n553), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n547), .A2(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n317), .A2(G303), .ZN(new_n559));
  INV_X1    g0359(.A(G257), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n353), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n353), .A2(G264), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n294), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n282), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n489), .A2(G270), .A3(new_n282), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n492), .ZN(new_n566));
  OAI21_X1  g0366(.A(G169), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n546), .B1(new_n558), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n563), .ZN(new_n569));
  INV_X1    g0369(.A(G303), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n314), .B2(new_n316), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n279), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n566), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n337), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n556), .A2(new_n557), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n548), .B1(G116), .B2(new_n472), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(KEYINPUT21), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n565), .A2(G179), .A3(new_n492), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n564), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n575), .B2(new_n576), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n568), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n572), .A2(new_n573), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G200), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n572), .A2(new_n573), .A3(new_n281), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n583), .A2(new_n558), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n213), .B(G87), .C1(new_n274), .C2(new_n275), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n588));
  OR3_X1    g0388(.A1(new_n512), .A2(KEYINPUT22), .A3(G20), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n317), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n213), .A2(KEYINPUT23), .A3(G107), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  OAI22_X1  g0393(.A1(new_n592), .A2(KEYINPUT79), .B1(new_n593), .B2(new_n462), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n462), .A3(G20), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT79), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n597));
  OAI22_X1  g0397(.A1(new_n595), .A2(new_n596), .B1(new_n597), .B2(G20), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n590), .A2(new_n591), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n591), .B1(new_n590), .B2(new_n599), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n253), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n462), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT25), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n373), .B2(G107), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n462), .B2(new_n472), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n489), .A2(G264), .A3(new_n282), .ZN(new_n609));
  NOR2_X1   g0409(.A1(G250), .A2(G1698), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n560), .B2(G1698), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n294), .B1(G33), .B2(G294), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n609), .B(new_n492), .C1(new_n612), .C2(new_n282), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n286), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(G190), .B2(new_n613), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n602), .A2(new_n608), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n337), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(G179), .B2(new_n613), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n602), .B2(new_n608), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n545), .A2(new_n586), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n461), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n400), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT82), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n309), .B1(new_n506), .B2(G68), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n334), .B1(KEYINPUT16), .B2(new_n626), .ZN(new_n627));
  AOI211_X1 g0427(.A(new_n325), .B(new_n339), .C1(new_n627), .C2(new_n258), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT18), .B1(new_n341), .B2(new_n342), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n340), .A2(KEYINPUT82), .A3(new_n343), .ZN(new_n631));
  INV_X1    g0431(.A(new_n449), .ZN(new_n632));
  INV_X1    g0432(.A(new_n459), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n632), .B1(new_n454), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT17), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n323), .B(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n630), .B(new_n631), .C1(new_n634), .C2(new_n636), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n408), .B(new_n411), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n624), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT80), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n526), .A2(new_n640), .ZN(new_n641));
  AOI211_X1 g0441(.A(KEYINPUT80), .B(new_n282), .C1(new_n524), .C2(new_n525), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n534), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(G200), .B1(G190), .B2(new_n531), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n542), .A2(new_n518), .A3(new_n519), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT81), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n541), .A2(KEYINPUT81), .A3(new_n542), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n520), .A2(new_n532), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(new_n337), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n644), .A2(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n337), .B1(new_n483), .B2(new_n493), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n498), .A2(new_n499), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(G179), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n470), .B2(new_n473), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n652), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n504), .A2(new_n508), .A3(new_n533), .A4(new_n543), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n659), .A2(KEYINPUT26), .B1(new_n650), .B2(new_n651), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n616), .B(new_n652), .C1(new_n581), .C2(new_n620), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n501), .A2(new_n509), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n658), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n461), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n639), .A2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n243), .A2(new_n213), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n558), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT83), .ZN(new_n674));
  MUX2_X1   g0474(.A(new_n581), .B(new_n586), .S(new_n674), .Z(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n590), .A2(new_n599), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT24), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n590), .A2(new_n591), .A3(new_n599), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n333), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n671), .B1(new_n680), .B2(new_n607), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n621), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n620), .A2(new_n671), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n676), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n581), .A2(new_n672), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n688), .A2(new_n620), .A3(new_n617), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n620), .B2(new_n672), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n207), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n513), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n210), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT86), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n652), .A2(new_n656), .A3(new_n700), .A4(KEYINPUT26), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT80), .B1(new_n537), .B2(new_n282), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n526), .A2(new_n640), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n530), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n532), .B(new_n520), .C1(new_n704), .C2(G169), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n541), .A2(KEYINPUT81), .A3(new_n542), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT81), .B1(new_n541), .B2(new_n542), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n540), .B1(new_n704), .B2(new_n286), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n710), .A2(new_n657), .A3(new_n509), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT86), .B1(new_n659), .B2(new_n657), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n701), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n500), .A2(new_n494), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n508), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT87), .B1(new_n656), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n613), .A2(G179), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n337), .B2(new_n613), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n680), .B2(new_n607), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(new_n568), .A3(new_n580), .A4(new_n577), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n644), .A2(new_n649), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n721), .A2(new_n616), .A3(new_n705), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT87), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n501), .A2(new_n509), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n716), .A2(new_n720), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n713), .A2(new_n705), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n699), .B1(new_n726), .B2(new_n672), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n663), .A2(new_n672), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n613), .A2(new_n455), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n654), .A3(new_n643), .A4(new_n582), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n560), .A2(G1698), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G250), .B2(G1698), .ZN(new_n734));
  INV_X1    g0534(.A(G294), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(new_n298), .B1(new_n249), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n279), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n609), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n538), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n483), .A2(new_n493), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n579), .A2(new_n739), .A3(KEYINPUT30), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n732), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n579), .A2(new_n739), .A3(new_n740), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT30), .B1(new_n744), .B2(KEYINPUT84), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT84), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n579), .A2(new_n739), .A3(new_n746), .A4(new_n740), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT85), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n279), .B1(new_n485), .B2(new_n491), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n279), .A2(new_n736), .B1(new_n749), .B2(G264), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n498), .A2(new_n750), .A3(new_n499), .A4(new_n531), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n572), .A2(new_n573), .A3(G179), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT84), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n753), .A2(new_n747), .A3(KEYINPUT85), .A4(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n743), .B1(new_n748), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT31), .B1(new_n757), .B2(new_n671), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n545), .A2(new_n586), .A3(new_n621), .A4(new_n672), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n753), .A2(new_n754), .A3(new_n747), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n743), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT31), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n672), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(G330), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n730), .A2(new_n766), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT88), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT88), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n698), .B1(new_n770), .B2(G1), .ZN(G364));
  NAND2_X1  g0571(.A1(new_n213), .A2(G13), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n243), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n693), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n675), .B2(G330), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n675), .ZN(new_n778));
  INV_X1    g0578(.A(new_n776), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n212), .B1(G20), .B2(new_n337), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT90), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT90), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT32), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G179), .A2(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(new_n213), .A3(G190), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n785), .B1(new_n788), .B2(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n213), .A2(new_n455), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n286), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n281), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n281), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n202), .A2(new_n793), .B1(new_n795), .B2(new_n303), .ZN(new_n796));
  INV_X1    g0596(.A(new_n792), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G190), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n789), .B(new_n796), .C1(G68), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n213), .A2(G179), .ZN(new_n800));
  INV_X1    g0600(.A(G190), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n800), .A2(new_n801), .A3(G200), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n462), .ZN(new_n803));
  INV_X1    g0603(.A(new_n788), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n804), .A2(KEYINPUT32), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n794), .A2(new_n801), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n803), .B(new_n806), .C1(new_n217), .C2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n800), .A2(G190), .A3(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n317), .B1(G87), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT91), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(G20), .B1(new_n787), .B2(new_n801), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT92), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n820), .A2(G97), .B1(new_n813), .B2(new_n812), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n799), .A2(new_n809), .A3(new_n814), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n317), .ZN(new_n823));
  INV_X1    g0623(.A(G326), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n824), .A2(new_n793), .B1(new_n807), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n823), .B(new_n826), .C1(G329), .C2(new_n788), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n820), .A2(G294), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT33), .B(G317), .ZN(new_n829));
  INV_X1    g0629(.A(new_n802), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n798), .A2(new_n829), .B1(G283), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n795), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G322), .B1(G303), .B2(new_n811), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n827), .A2(new_n828), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n784), .B1(new_n822), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(G13), .A2(G33), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(G20), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n783), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n238), .A2(new_n484), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n692), .A2(new_n294), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n484), .B2(new_n211), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n317), .A2(new_n692), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G355), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(G116), .B2(new_n207), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n840), .A2(new_n843), .B1(new_n846), .B2(KEYINPUT89), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(KEYINPUT89), .B2(new_n846), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n779), .B(new_n835), .C1(new_n839), .C2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n838), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n675), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n778), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G396));
  NOR2_X1   g0653(.A1(new_n783), .A2(new_n836), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n820), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(new_n303), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n298), .B1(new_n788), .B2(G132), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n858), .B1(new_n202), .B2(new_n810), .C1(new_n304), .C2(new_n802), .ZN(new_n859));
  INV_X1    g0659(.A(new_n793), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G137), .A2(new_n860), .B1(new_n808), .B2(G159), .ZN(new_n861));
  INV_X1    g0661(.A(G143), .ZN(new_n862));
  INV_X1    g0662(.A(new_n798), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n861), .B1(new_n862), .B2(new_n795), .C1(new_n392), .C2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT34), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n857), .B(new_n859), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G283), .A2(new_n798), .B1(new_n860), .B2(G303), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n552), .B2(new_n807), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT93), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n317), .B1(new_n804), .B2(new_n825), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n832), .A2(G294), .B1(G87), .B2(new_n830), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n462), .B2(new_n810), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n871), .B(new_n873), .C1(G97), .C2(new_n820), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n866), .A2(new_n867), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n776), .B1(G77), .B2(new_n855), .C1(new_n875), .C2(new_n784), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n459), .A2(new_n671), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n383), .A2(new_n378), .B1(new_n377), .B2(new_n672), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n459), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n876), .B1(new_n880), .B2(new_n836), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n728), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n377), .A2(new_n672), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n379), .A2(new_n382), .ZN(new_n884));
  INV_X1    g0684(.A(new_n378), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n663), .A2(new_n886), .A3(new_n459), .A4(new_n672), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n888), .A2(new_n766), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n776), .B1(new_n888), .B2(new_n766), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n881), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(G384));
  AOI22_X1  g0692(.A1(new_n622), .A2(new_n672), .B1(new_n757), .B2(new_n763), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n757), .A2(new_n671), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT97), .B1(new_n894), .B2(new_n762), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT85), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n760), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n742), .B1(new_n897), .B2(new_n755), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT97), .B(new_n762), .C1(new_n898), .C2(new_n672), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n893), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n428), .A2(new_n672), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n449), .A2(new_n454), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(G169), .B1(new_n450), .B2(new_n451), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT14), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n454), .A2(new_n906), .A3(new_n446), .A4(new_n445), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT94), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n908), .A3(new_n902), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n908), .B1(new_n907), .B2(new_n902), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT95), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n911), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT95), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(new_n904), .A4(new_n909), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT16), .B1(new_n302), .B2(new_n321), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n258), .B1(new_n313), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n669), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n628), .A2(new_n629), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n636), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT37), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n323), .B1(new_n335), .B2(new_n669), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n339), .B1(new_n627), .B2(new_n258), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n918), .B1(new_n342), .B2(new_n919), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(KEYINPUT37), .A3(new_n323), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n923), .A2(KEYINPUT38), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT38), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n920), .B1(new_n324), .B2(new_n344), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n927), .A2(new_n929), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n901), .A2(new_n916), .A3(new_n935), .A4(new_n879), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n323), .B(new_n625), .C1(new_n335), .C2(new_n669), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT37), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n341), .A2(new_n342), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n941), .B(new_n323), .C1(new_n335), .C2(new_n669), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n323), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n669), .B1(new_n627), .B2(new_n258), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n946), .A2(KEYINPUT82), .A3(KEYINPUT37), .A4(new_n941), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n630), .A2(new_n324), .A3(new_n631), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n948), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n930), .B1(new_n950), .B2(KEYINPUT38), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n762), .B1(new_n898), .B2(new_n672), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT97), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n899), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n880), .B1(new_n955), .B2(new_n893), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n951), .A2(new_n956), .A3(KEYINPUT40), .A4(new_n916), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n938), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n901), .A2(new_n461), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  INV_X1    g0761(.A(G330), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT98), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT39), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n949), .A2(new_n945), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n946), .A2(new_n941), .B1(new_n939), .B2(KEYINPUT37), .ZN(new_n968));
  NOR4_X1   g0768(.A1(new_n925), .A2(new_n625), .A3(new_n926), .A4(new_n924), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT38), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n932), .A2(new_n933), .A3(new_n931), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n632), .A2(new_n672), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n930), .A2(new_n934), .A3(KEYINPUT39), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n973), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT96), .ZN(new_n978));
  INV_X1    g0778(.A(new_n877), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n887), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n916), .A2(new_n935), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n919), .B1(new_n630), .B2(new_n631), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n978), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n912), .A2(new_n915), .B1(new_n887), .B2(new_n979), .ZN(new_n986));
  AOI211_X1 g0786(.A(KEYINPUT96), .B(new_n982), .C1(new_n986), .C2(new_n935), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n461), .B1(new_n727), .B2(new_n729), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n639), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n989), .B(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n965), .A2(new_n992), .B1(G1), .B2(new_n772), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n965), .B2(new_n992), .ZN(new_n994));
  INV_X1    g0794(.A(new_n468), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT35), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(KEYINPUT35), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n996), .A2(G116), .A3(new_n214), .A4(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT36), .Z(new_n999));
  OAI211_X1 g0799(.A(new_n217), .B(new_n211), .C1(new_n303), .C2(new_n304), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n202), .A2(G68), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n243), .B(G13), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n994), .A2(new_n1003), .ZN(G367));
  NAND2_X1  g0804(.A1(new_n508), .A2(new_n671), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n716), .A2(new_n724), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n656), .A2(new_n671), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n1006), .A2(KEYINPUT99), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT99), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n689), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT42), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n620), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n671), .B1(new_n1014), .B2(new_n509), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT43), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n708), .A2(new_n671), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(new_n705), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n652), .B2(new_n1017), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1013), .A2(new_n1015), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1016), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n687), .A2(new_n1010), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n693), .B(KEYINPUT41), .Z(new_n1026));
  INV_X1    g0826(.A(new_n690), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1010), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT44), .Z(new_n1029));
  NOR2_X1   g0829(.A1(new_n1010), .A2(new_n1027), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT45), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n687), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n687), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n685), .A2(new_n688), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1036), .A2(KEYINPUT100), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(KEYINPUT100), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n689), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(new_n676), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1035), .A2(new_n770), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1026), .B1(new_n1042), .B2(new_n770), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1024), .B(new_n1025), .C1(new_n1043), .C2(new_n775), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n839), .B1(new_n207), .B2(new_n364), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n234), .A2(new_n842), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n776), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G311), .A2(new_n860), .B1(new_n808), .B2(G283), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n830), .A2(G97), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n570), .C2(new_n795), .ZN(new_n1050));
  INV_X1    g0850(.A(G317), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n298), .B1(new_n804), .B2(new_n1051), .C1(new_n863), .C2(new_n735), .ZN(new_n1052));
  AOI21_X1  g0852(.A(KEYINPUT46), .B1(new_n811), .B2(G116), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n811), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT101), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n820), .A2(G107), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(KEYINPUT101), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n856), .A2(new_n304), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G150), .A2(new_n832), .B1(new_n808), .B2(G50), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n798), .A2(G159), .B1(G58), .B2(new_n811), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n860), .A2(G143), .B1(new_n217), .B2(new_n830), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n317), .B1(G137), .B2(new_n788), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1059), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n784), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1047), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1019), .A2(new_n838), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1044), .A2(new_n1072), .ZN(G387));
  OR2_X1    g0873(.A1(new_n231), .A2(new_n484), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n695), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1074), .A2(new_n841), .B1(new_n1075), .B2(new_n844), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n695), .B(new_n484), .C1(new_n304), .C2(new_n417), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT50), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n361), .B2(new_n202), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n255), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1076), .A2(new_n1081), .B1(G107), .B2(new_n207), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n779), .B1(new_n1082), .B2(new_n839), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n684), .B2(new_n850), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n798), .A2(G311), .B1(new_n808), .B2(G303), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT104), .B(G322), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1085), .B1(new_n1051), .B2(new_n795), .C1(new_n793), .C2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT105), .Z(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1089), .A2(KEYINPUT48), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(KEYINPUT48), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n856), .A2(new_n474), .B1(new_n735), .B2(new_n810), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(KEYINPUT49), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(KEYINPUT49), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n298), .B1(new_n552), .B2(new_n802), .C1(new_n804), .C2(new_n824), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G159), .A2(new_n860), .B1(new_n808), .B2(G68), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n202), .B2(new_n795), .C1(new_n255), .C2(new_n863), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n298), .B1(new_n788), .B2(G150), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n811), .A2(new_n217), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n1049), .A3(new_n1101), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT103), .Z(new_n1103));
  NOR2_X1   g0903(.A1(new_n856), .A2(new_n364), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1099), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1084), .B1(new_n1106), .B2(new_n783), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1041), .B2(new_n775), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1041), .A2(new_n770), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1040), .A2(new_n768), .A3(new_n769), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n693), .B(KEYINPUT106), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(G393));
  OAI21_X1  g0913(.A(new_n1109), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1042), .A2(new_n1114), .A3(new_n1111), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n825), .A2(new_n795), .B1(new_n793), .B2(new_n1051), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT107), .Z(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT52), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n856), .A2(new_n552), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n317), .B1(new_n804), .B2(new_n1086), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n803), .B1(new_n808), .B2(G294), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n474), .B2(new_n810), .C1(new_n570), .C2(new_n863), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n392), .A2(new_n793), .B1(new_n795), .B2(new_n805), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT51), .Z(new_n1125));
  NOR2_X1   g0925(.A1(new_n856), .A2(new_n417), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n294), .B1(new_n512), .B2(new_n802), .C1(new_n804), .C2(new_n862), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n808), .A2(new_n361), .B1(G68), .B2(new_n811), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n202), .B2(new_n863), .ZN(new_n1129));
  NOR4_X1   g0929(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n783), .B1(new_n1123), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n241), .A2(new_n842), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n839), .B1(new_n465), .B2(new_n207), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n776), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n1010), .B2(new_n838), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n1035), .B2(new_n775), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1115), .A2(new_n1136), .ZN(G390));
  OAI211_X1 g0937(.A(new_n879), .B(G330), .C1(new_n758), .C2(new_n765), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT109), .B1(new_n1139), .B2(new_n916), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n901), .A2(new_n916), .A3(G330), .A4(new_n879), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT109), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1138), .A2(new_n1142), .A3(new_n915), .A4(new_n912), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n901), .A2(new_n879), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n915), .B(new_n912), .C1(new_n1145), .C2(new_n962), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n878), .A2(new_n459), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n726), .A2(new_n672), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n979), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n1139), .B2(new_n916), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1144), .A2(new_n980), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n901), .A2(G330), .A3(new_n461), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(new_n639), .A3(new_n990), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n974), .B1(new_n971), .B2(new_n972), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1148), .A2(new_n979), .B1(new_n912), .B2(new_n915), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT108), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1149), .A2(new_n916), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT108), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1158), .A2(new_n951), .A3(new_n1159), .A4(new_n974), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n986), .A2(new_n975), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n973), .A2(new_n976), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1141), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1139), .A2(new_n916), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1161), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1154), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1157), .A2(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1170), .B2(new_n1141), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1144), .A2(new_n980), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1153), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1169), .A2(new_n1177), .A3(new_n1111), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1161), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(new_n1165), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1163), .A2(new_n836), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G107), .A2(new_n798), .B1(new_n860), .B2(G283), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n465), .B2(new_n807), .C1(new_n552), .C2(new_n795), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n811), .A2(G87), .B1(new_n830), .B2(G68), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1184), .B(new_n317), .C1(new_n735), .C2(new_n804), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1183), .A2(new_n1126), .A3(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n798), .A2(G137), .B1(G50), .B2(new_n830), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT54), .B(G143), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n807), .B2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G128), .A2(new_n860), .B1(new_n832), .B2(G132), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n810), .A2(new_n392), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT53), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n317), .B1(G125), .B2(new_n788), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1189), .B(new_n1194), .C1(G159), .C2(new_n820), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n783), .B1(new_n1186), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n779), .B1(new_n854), .B2(new_n255), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1181), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT110), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT110), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1180), .A2(new_n775), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1178), .A2(new_n1201), .ZN(G378));
  NAND2_X1  g1002(.A1(new_n397), .A2(new_n919), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n414), .A2(KEYINPUT115), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT115), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n638), .A2(new_n1205), .A3(new_n400), .ZN(new_n1206));
  XOR2_X1   g1006(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1204), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1203), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1207), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1203), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1204), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n836), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n776), .B1(new_n855), .B2(G50), .ZN(new_n1219));
  INV_X1    g1019(.A(G132), .ZN(new_n1220));
  INV_X1    g1020(.A(G137), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n863), .A2(new_n1220), .B1(new_n1221), .B2(new_n807), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT113), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1188), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n860), .A2(G125), .B1(new_n811), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n832), .A2(G128), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n856), .C2(new_n392), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1223), .A2(new_n1227), .ZN(new_n1228));
  XOR2_X1   g1028(.A(KEYINPUT114), .B(KEYINPUT59), .Z(new_n1229));
  OR2_X1    g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n830), .A2(G159), .ZN(new_n1232));
  AOI211_X1 g1032(.A(G33), .B(G41), .C1(new_n788), .C2(G124), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n294), .A2(G41), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G283), .B2(new_n788), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1236), .B(new_n1101), .C1(new_n303), .C2(new_n802), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT111), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G97), .A2(new_n798), .B1(new_n860), .B2(G116), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n462), .B2(new_n795), .C1(new_n364), .C2(new_n807), .ZN(new_n1240));
  OR3_X1    g1040(.A1(new_n1238), .A2(new_n1240), .A3(new_n1060), .ZN(new_n1241));
  XOR2_X1   g1041(.A(KEYINPUT112), .B(KEYINPUT58), .Z(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1235), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1234), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1219), .B1(new_n1246), .B2(new_n783), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1218), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1217), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n936), .A2(new_n937), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n901), .A2(new_n916), .A3(new_n879), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT40), .B1(new_n971), .B2(new_n972), .ZN(new_n1252));
  OAI21_X1  g1052(.A(G330), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1249), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n938), .A2(new_n1217), .A3(new_n957), .A4(G330), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n989), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n977), .A2(new_n987), .A3(new_n984), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n1255), .A3(new_n1254), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1248), .B1(new_n1260), .B2(new_n774), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1111), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1258), .A2(new_n1255), .A3(new_n1254), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1254), .A2(new_n1255), .B1(new_n985), .B2(new_n988), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT57), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1175), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1262), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1153), .B1(new_n1180), .B2(new_n1154), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1265), .B1(new_n1269), .B2(new_n1260), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1261), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(G375));
  INV_X1    g1072(.A(KEYINPUT116), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1151), .B2(new_n774), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1174), .A2(KEYINPUT116), .A3(new_n775), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n776), .B1(new_n855), .B2(G68), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n1220), .A2(new_n793), .B1(new_n795), .B2(new_n1221), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n798), .B2(new_n1224), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n807), .A2(new_n392), .B1(new_n810), .B2(new_n805), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n298), .B1(new_n788), .B2(G128), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n303), .B2(new_n802), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1278), .B(new_n1282), .C1(new_n202), .C2(new_n856), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n798), .A2(G116), .B1(new_n808), .B2(G107), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n860), .A2(G294), .B1(G97), .B2(new_n811), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n823), .B1(G303), .B2(new_n788), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n832), .A2(G283), .B1(G77), .B2(new_n830), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1284), .A2(new_n1285), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1283), .B1(new_n1104), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1276), .B1(new_n1289), .B2(new_n783), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n916), .B2(new_n837), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1274), .A2(new_n1275), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1026), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1176), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(G381));
  INV_X1    g1096(.A(G387), .ZN(new_n1297));
  INV_X1    g1097(.A(G390), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1108), .A2(new_n1112), .A3(new_n852), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1297), .A2(new_n891), .A3(new_n1298), .A4(new_n1300), .ZN(new_n1301));
  OR4_X1    g1101(.A1(G378), .A2(new_n1301), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1102(.A(G378), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n670), .A2(G213), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1271), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G407), .A2(G213), .A3(new_n1306), .ZN(G409));
  INV_X1    g1107(.A(KEYINPUT120), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n852), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1309));
  OR3_X1    g1109(.A1(new_n1300), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1308), .B1(new_n1300), .B2(new_n1309), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT121), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1312), .B(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G390), .A2(KEYINPUT122), .ZN(new_n1315));
  OR2_X1    g1115(.A1(G390), .A2(KEYINPUT122), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1297), .B2(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1297), .A2(new_n1316), .A3(new_n1315), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1314), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  AND2_X1   g1119(.A1(G387), .A2(KEYINPUT123), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1312), .B1(new_n1320), .B2(new_n1298), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1298), .B2(new_n1320), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1319), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT60), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1293), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1151), .A2(KEYINPUT60), .A3(new_n1153), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1325), .A2(new_n1111), .A3(new_n1176), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1292), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(new_n891), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1327), .A2(new_n1292), .A3(G384), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(G2897), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1304), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1331), .A2(KEYINPUT119), .A3(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT119), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1330), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G384), .B1(new_n1327), .B2(new_n1292), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1333), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1335), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT118), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1331), .A2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT118), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1334), .B(new_n1340), .C1(new_n1344), .C2(new_n1333), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1346), .A2(new_n1267), .A3(new_n1294), .ZN(new_n1347));
  AOI22_X1  g1147(.A1(new_n1346), .A2(new_n775), .B1(new_n1218), .B2(new_n1247), .ZN(new_n1348));
  AOI21_X1  g1148(.A(G378), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(KEYINPUT117), .B1(new_n1271), .B2(G378), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1257), .A2(KEYINPUT57), .A3(new_n1259), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1111), .B1(new_n1269), .B2(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(KEYINPUT57), .B1(new_n1346), .B2(new_n1267), .ZN(new_n1354));
  OAI211_X1 g1154(.A(G378), .B(new_n1348), .C1(new_n1353), .C2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT117), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1350), .B1(new_n1351), .B2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1345), .B1(new_n1304), .B2(new_n1358), .ZN(new_n1359));
  NOR3_X1   g1159(.A1(new_n1323), .A2(KEYINPUT61), .A3(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT124), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1358), .A2(new_n1361), .A3(new_n1304), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1364));
  NAND4_X1  g1164(.A1(new_n1364), .A2(KEYINPUT117), .A3(G378), .A4(new_n1348), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1349), .B1(new_n1363), .B2(new_n1365), .ZN(new_n1366));
  OAI21_X1  g1166(.A(KEYINPUT124), .B1(new_n1366), .B2(new_n1305), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1344), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1362), .A2(new_n1367), .A3(KEYINPUT63), .A4(new_n1368), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1368), .A2(new_n1358), .A3(new_n1304), .ZN(new_n1370));
  INV_X1    g1170(.A(KEYINPUT63), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1360), .A2(new_n1369), .A3(new_n1372), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT125), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1345), .B1(new_n1362), .B2(new_n1367), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1374), .B1(new_n1375), .B2(KEYINPUT61), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1340), .A2(new_n1334), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1377), .B1(new_n1368), .B2(new_n1339), .ZN(new_n1378));
  AOI21_X1  g1178(.A(new_n1361), .B1(new_n1358), .B2(new_n1304), .ZN(new_n1379));
  NOR3_X1   g1179(.A1(new_n1366), .A2(KEYINPUT124), .A3(new_n1305), .ZN(new_n1380));
  OAI21_X1  g1180(.A(new_n1378), .B1(new_n1379), .B2(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(KEYINPUT61), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1381), .A2(KEYINPUT125), .A3(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT62), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1370), .A2(new_n1384), .ZN(new_n1385));
  NAND4_X1  g1185(.A1(new_n1362), .A2(new_n1367), .A3(KEYINPUT62), .A4(new_n1368), .ZN(new_n1386));
  AOI22_X1  g1186(.A1(new_n1376), .A2(new_n1383), .B1(new_n1385), .B2(new_n1386), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT126), .ZN(new_n1388));
  OAI21_X1  g1188(.A(new_n1323), .B1(new_n1387), .B2(new_n1388), .ZN(new_n1389));
  AND2_X1   g1189(.A1(new_n1386), .A2(new_n1385), .ZN(new_n1390));
  AOI211_X1 g1190(.A(KEYINPUT126), .B(new_n1390), .C1(new_n1376), .C2(new_n1383), .ZN(new_n1391));
  OAI21_X1  g1191(.A(new_n1373), .B1(new_n1389), .B2(new_n1391), .ZN(G405));
  NAND2_X1  g1192(.A1(new_n1323), .A2(KEYINPUT127), .ZN(new_n1393));
  OAI22_X1  g1193(.A1(new_n1351), .A2(new_n1357), .B1(G378), .B2(new_n1271), .ZN(new_n1394));
  NOR2_X1   g1194(.A1(new_n1394), .A2(new_n1331), .ZN(new_n1395));
  INV_X1    g1195(.A(new_n1395), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1394), .A2(new_n1344), .ZN(new_n1397));
  NAND3_X1  g1197(.A1(new_n1393), .A2(new_n1396), .A3(new_n1397), .ZN(new_n1398));
  NOR2_X1   g1198(.A1(new_n1323), .A2(KEYINPUT127), .ZN(new_n1399));
  XNOR2_X1  g1199(.A(new_n1398), .B(new_n1399), .ZN(G402));
endmodule


