//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912;
  INV_X1    g000(.A(G211gat), .ZN(new_n202));
  INV_X1    g001(.A(G218gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT22), .ZN(new_n204));
  NAND2_X1  g003(.A1(G211gat), .A2(G218gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(KEYINPUT74), .A3(new_n207), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n207), .A2(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G211gat), .B2(G218gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT28), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  AND2_X1   g016(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(KEYINPUT65), .ZN(new_n226));
  AOI211_X1 g025(.A(new_n221), .B(KEYINPUT66), .C1(new_n220), .C2(KEYINPUT64), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT27), .B(G183gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(new_n217), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT66), .B1(new_n231), .B2(new_n221), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n225), .A2(KEYINPUT65), .A3(new_n224), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n222), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G169gat), .ZN(new_n235));
  INV_X1    g034(.A(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT26), .ZN(new_n238));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n240), .B(new_n241), .C1(new_n238), .C2(new_n237), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n234), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n241), .B(KEYINPUT24), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(G183gat), .B2(G190gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n237), .B(KEYINPUT23), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n239), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n247), .A4(new_n239), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n244), .A2(KEYINPUT75), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT75), .B1(new_n244), .B2(new_n252), .ZN(new_n254));
  INV_X1    g053(.A(G226gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n253), .A2(new_n254), .A3(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n250), .A2(new_n251), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n244), .A2(KEYINPUT67), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n228), .A2(new_n234), .A3(new_n264), .A4(new_n243), .ZN(new_n265));
  AOI211_X1 g064(.A(new_n258), .B(new_n262), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n215), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT76), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n257), .B1(new_n253), .B2(new_n254), .ZN(new_n270));
  INV_X1    g069(.A(new_n215), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n270), .B(new_n271), .C1(new_n260), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n244), .A2(new_n252), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n244), .A2(new_n252), .A3(KEYINPUT75), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(new_n259), .A3(new_n258), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n265), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n257), .A3(new_n252), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(KEYINPUT76), .A3(new_n215), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT77), .B(G64gat), .Z(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT78), .B(G92gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n269), .A2(new_n273), .A3(new_n282), .A4(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT79), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT80), .B1(new_n291), .B2(KEYINPUT30), .ZN(new_n292));
  XOR2_X1   g091(.A(G1gat), .B(G29gat), .Z(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT86), .ZN(new_n294));
  XOR2_X1   g093(.A(KEYINPUT85), .B(KEYINPUT0), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G57gat), .B(G85gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G120gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT70), .B(G113gat), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT1), .ZN(new_n305));
  INV_X1    g104(.A(G134gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G127gat), .ZN(new_n307));
  INV_X1    g106(.A(G127gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G134gat), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n304), .A2(new_n305), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n303), .A2(G113gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n305), .B1(new_n300), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT68), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n306), .B2(G127gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n308), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(new_n307), .A3(new_n316), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n312), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n313), .B1(new_n312), .B2(new_n317), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n310), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G155gat), .ZN(new_n322));
  INV_X1    g121(.A(G155gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(KEYINPUT82), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT82), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G155gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n328), .A3(G162gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n329), .B2(KEYINPUT2), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G148gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT81), .B(G148gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n331), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G141gat), .B(G148gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n325), .B1(new_n336), .B2(KEYINPUT2), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n320), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n320), .A2(new_n338), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(KEYINPUT4), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n335), .A2(new_n346), .A3(new_n337), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n320), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT83), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n345), .A2(KEYINPUT83), .A3(new_n320), .A4(new_n347), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n320), .A2(KEYINPUT71), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT71), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n310), .B(new_n355), .C1(new_n318), .C2(new_n319), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n338), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n341), .B1(new_n357), .B2(KEYINPUT4), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n352), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n353), .B1(new_n352), .B2(new_n358), .ZN(new_n360));
  OAI211_X1 g159(.A(KEYINPUT5), .B(new_n342), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n350), .A2(new_n351), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n343), .A2(KEYINPUT4), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n362), .B(new_n363), .C1(KEYINPUT4), .C2(new_n357), .ZN(new_n364));
  OR3_X1    g163(.A1(new_n364), .A2(KEYINPUT5), .A3(new_n341), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n298), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT6), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n361), .A2(new_n365), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT87), .ZN(new_n369));
  INV_X1    g168(.A(new_n298), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n361), .A2(new_n365), .A3(new_n298), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n366), .A2(new_n369), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n367), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT76), .B1(new_n281), .B2(new_n215), .ZN(new_n377));
  AOI211_X1 g176(.A(new_n268), .B(new_n271), .C1(new_n278), .C2(new_n280), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n273), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n287), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(new_n289), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n379), .A2(new_n290), .A3(new_n273), .A4(new_n288), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n289), .A2(KEYINPUT79), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n382), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n292), .A2(new_n376), .A3(new_n384), .A4(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT31), .B(G50gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT88), .ZN(new_n394));
  INV_X1    g193(.A(new_n338), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n214), .B1(new_n212), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT89), .B1(new_n210), .B2(new_n211), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n259), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n395), .B1(new_n399), .B2(new_n346), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n347), .A2(new_n259), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(new_n215), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n394), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT90), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(G22gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT3), .B1(new_n215), .B2(new_n259), .ZN(new_n408));
  OAI221_X1 g207(.A(new_n393), .B1(new_n401), .B2(new_n215), .C1(new_n395), .C2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n404), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n407), .B1(new_n404), .B2(new_n409), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n392), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n412), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(new_n391), .A3(new_n410), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n413), .A2(new_n415), .A3(KEYINPUT91), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT91), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n390), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n279), .A2(new_n252), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n354), .A2(new_n356), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n272), .A2(new_n354), .A3(new_n356), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT32), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G15gat), .B(G43gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT72), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(G71gat), .ZN(new_n431));
  INV_X1    g230(.A(G99gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n426), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n433), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n425), .B(KEYINPUT32), .C1(new_n427), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n423), .B1(new_n422), .B2(new_n424), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT34), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n438), .B(KEYINPUT34), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(new_n434), .A3(new_n436), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT36), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(KEYINPUT73), .A3(new_n443), .ZN(new_n446));
  OR3_X1    g245(.A1(new_n437), .A2(KEYINPUT73), .A3(new_n440), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n445), .B1(new_n448), .B2(KEYINPUT36), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n419), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT93), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n364), .A2(KEYINPUT92), .A3(new_n341), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT92), .B1(new_n364), .B2(new_n341), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n455), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n453), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT39), .B1(new_n339), .B2(new_n341), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n456), .B(new_n298), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT40), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n368), .A2(new_n370), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n461), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n388), .B1(new_n387), .B2(new_n382), .ZN(new_n466));
  AOI211_X1 g265(.A(KEYINPUT80), .B(KEYINPUT30), .C1(new_n385), .C2(new_n386), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n465), .B1(new_n468), .B2(new_n384), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n413), .A2(new_n415), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n372), .A3(new_n373), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n269), .A2(new_n472), .A3(new_n282), .A4(new_n273), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT38), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n281), .A2(new_n271), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n270), .B1(new_n260), .B2(new_n272), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n475), .B(KEYINPUT37), .C1(new_n271), .C2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n473), .A2(new_n474), .A3(new_n477), .A4(new_n287), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n387), .A2(new_n471), .A3(new_n367), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n380), .A2(KEYINPUT37), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n473), .A2(new_n287), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n470), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n451), .B1(new_n469), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n465), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n292), .A2(new_n384), .A3(new_n389), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n483), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT93), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n450), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n448), .A2(new_n384), .A3(new_n292), .A4(new_n389), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n367), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT35), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n470), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT94), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n444), .A2(new_n470), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT35), .B1(new_n390), .B2(new_n496), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n466), .A2(new_n467), .A3(new_n383), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n499));
  INV_X1    g298(.A(new_n494), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n448), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n495), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT95), .B1(new_n490), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n450), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n469), .A2(new_n451), .A3(new_n483), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT93), .B1(new_n487), .B2(new_n488), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT95), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n495), .A2(new_n497), .A3(new_n501), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT14), .ZN(new_n515));
  NAND2_X1  g314(.A1(G29gat), .A2(G36gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G43gat), .B(G50gat), .Z(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT96), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n518), .A2(new_n519), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n515), .C1(new_n522), .C2(new_n516), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n524), .B2(new_n520), .ZN(new_n525));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526));
  INV_X1    g325(.A(G85gat), .ZN(new_n527));
  INV_X1    g326(.A(G92gat), .ZN(new_n528));
  AOI22_X1  g327(.A1(KEYINPUT8), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530));
  OAI22_X1  g329(.A1(new_n527), .A2(new_n528), .B1(new_n530), .B2(KEYINPUT103), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT103), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G99gat), .B(G106gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT104), .ZN(new_n537));
  XOR2_X1   g336(.A(G190gat), .B(G218gat), .Z(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n525), .A2(new_n536), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT41), .ZN(new_n541));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n544), .A2(KEYINPUT97), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(KEYINPUT97), .ZN(new_n546));
  OAI22_X1  g345(.A1(new_n545), .A2(new_n546), .B1(new_n543), .B2(new_n525), .ZN(new_n547));
  OAI221_X1 g346(.A(new_n540), .B1(new_n541), .B2(new_n542), .C1(new_n547), .C2(new_n536), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n539), .A2(new_n537), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G134gat), .B(G162gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n542), .A2(new_n541), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n548), .A2(new_n549), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n550), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n550), .B2(new_n554), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT16), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(G1gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(G1gat), .B2(new_n559), .ZN(new_n562));
  INV_X1    g361(.A(G8gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G57gat), .B(G64gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT100), .ZN(new_n566));
  NAND2_X1  g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567));
  INV_X1    g366(.A(G71gat), .ZN(new_n568));
  INV_X1    g367(.A(G78gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n567), .B(new_n570), .C1(new_n565), .C2(new_n571), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT21), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n564), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n202), .ZN(new_n578));
  XOR2_X1   g377(.A(G127gat), .B(G155gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n576), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT101), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT102), .B(G183gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n584), .B(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n558), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n536), .A2(KEYINPUT10), .A3(new_n573), .A4(new_n574), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n575), .B(new_n536), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n593), .B2(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT105), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n592), .B2(new_n595), .ZN(new_n599));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G176gat), .B(G204gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n596), .B1(new_n592), .B2(new_n595), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(new_n602), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OAI221_X1 g409(.A(new_n564), .B1(new_n543), .B2(new_n525), .C1(new_n545), .C2(new_n546), .ZN(new_n611));
  INV_X1    g410(.A(new_n564), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n525), .ZN(new_n613));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n525), .B(new_n564), .Z(new_n618));
  XOR2_X1   g417(.A(new_n614), .B(KEYINPUT13), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(new_n616), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n611), .A2(new_n613), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n623), .A2(new_n614), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n624), .A2(KEYINPUT18), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(KEYINPUT98), .ZN(new_n627));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628));
  INV_X1    g427(.A(G197gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT11), .B(G169gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  NAND3_X1  g432(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n622), .B(new_n625), .C1(KEYINPUT98), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n511), .A2(new_n610), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n376), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT106), .B(G1gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1324gat));
  INV_X1    g440(.A(new_n638), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(KEYINPUT107), .A3(new_n486), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n563), .A2(KEYINPUT42), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT107), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n638), .B2(new_n498), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n638), .B2(new_n498), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT16), .B(G8gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n648), .B(new_n650), .C1(KEYINPUT108), .C2(KEYINPUT42), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n650), .A2(KEYINPUT108), .A3(KEYINPUT42), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(G1325gat));
  INV_X1    g452(.A(G15gat), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n638), .A2(new_n654), .A3(new_n449), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n642), .A2(new_n448), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(new_n654), .ZN(G1326gat));
  INV_X1    g456(.A(new_n418), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n638), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  OAI21_X1  g460(.A(new_n558), .B1(new_n490), .B2(new_n502), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n558), .B2(KEYINPUT95), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  OAI221_X1 g464(.A(new_n558), .B1(KEYINPUT95), .B2(new_n663), .C1(new_n490), .C2(new_n502), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n589), .B(KEYINPUT109), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n607), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n667), .A2(new_n637), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n376), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n558), .A2(new_n589), .A3(new_n608), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n503), .A2(new_n510), .A3(new_n637), .A4(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n376), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n673), .B1(new_n677), .B2(new_n512), .ZN(new_n678));
  NOR4_X1   g477(.A1(new_n676), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n376), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n672), .A2(new_n512), .B1(new_n678), .B2(new_n679), .ZN(G1328gat));
  AOI21_X1  g479(.A(new_n513), .B1(new_n670), .B2(new_n486), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n486), .A2(new_n513), .ZN(new_n683));
  OR3_X1    g482(.A1(new_n676), .A2(KEYINPUT46), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT46), .B1(new_n676), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n681), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n681), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(G1329gat));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690));
  INV_X1    g489(.A(new_n448), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(G43gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT112), .ZN(new_n696));
  INV_X1    g495(.A(new_n449), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n667), .A2(new_n637), .A3(new_n697), .A4(new_n669), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n693), .B1(new_n698), .B2(G43gat), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT112), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n700), .B(new_n690), .C1(new_n693), .C2(new_n694), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n696), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n699), .B1(new_n696), .B2(new_n701), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(G1330gat));
  NOR3_X1   g503(.A1(new_n676), .A2(G50gat), .A3(new_n658), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(KEYINPUT48), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n667), .A2(new_n637), .A3(new_n418), .A4(new_n669), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G50gat), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710));
  INV_X1    g509(.A(new_n470), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n667), .A2(new_n637), .A3(new_n711), .A4(new_n669), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  INV_X1    g512(.A(new_n705), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT113), .B1(new_n709), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n706), .A2(new_n708), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n705), .B1(new_n712), .B2(G50gat), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n717), .B(new_n718), .C1(new_n710), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n720), .ZN(G1331gat));
  AOI211_X1 g520(.A(new_n608), .B(new_n637), .C1(new_n507), .C2(new_n509), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n590), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n376), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT114), .B(G57gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1332gat));
  NOR2_X1   g525(.A1(new_n723), .A2(new_n498), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT49), .B(G64gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n727), .B2(new_n730), .ZN(G1333gat));
  OAI21_X1  g530(.A(new_n568), .B1(new_n723), .B2(new_n691), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n722), .A2(G71gat), .A3(new_n590), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n449), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1334gat));
  NOR2_X1   g535(.A1(new_n723), .A2(new_n658), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n569), .ZN(G1335gat));
  INV_X1    g537(.A(KEYINPUT116), .ZN(new_n739));
  INV_X1    g538(.A(new_n589), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n637), .A2(new_n740), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n667), .A2(new_n607), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(G85gat), .A3(new_n671), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n557), .B1(new_n507), .B2(new_n509), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n741), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(KEYINPUT51), .A3(new_n741), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n608), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n671), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n739), .B1(new_n744), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n750), .A2(new_n671), .ZN(new_n753));
  OAI211_X1 g552(.A(KEYINPUT116), .B(new_n743), .C1(new_n753), .C2(G85gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1336gat));
  AOI21_X1  g554(.A(new_n528), .B1(new_n742), .B2(new_n486), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n486), .A2(new_n528), .A3(new_n607), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT117), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n748), .B2(new_n749), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n756), .A2(KEYINPUT52), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT52), .B1(new_n756), .B2(new_n759), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1337gat));
  AOI21_X1  g561(.A(G99gat), .B1(new_n750), .B2(new_n448), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n742), .A2(G99gat), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n697), .ZN(G1338gat));
  INV_X1    g564(.A(G106gat), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n742), .B2(new_n418), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n750), .A2(new_n766), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n711), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n766), .B1(new_n742), .B2(new_n711), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n750), .A2(new_n766), .A3(new_n711), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n770), .ZN(new_n773));
  OAI22_X1  g572(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n773), .ZN(G1339gat));
  INV_X1    g573(.A(new_n668), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n594), .A2(new_n595), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(KEYINPUT54), .A3(new_n596), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n602), .B(new_n777), .C1(new_n598), .C2(KEYINPUT54), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n606), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n779), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n637), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n623), .A2(new_n614), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n618), .A2(new_n619), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n632), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n607), .B(new_n789), .C1(new_n626), .C2(new_n633), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n558), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n782), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n626), .B2(new_n633), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(new_n557), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n775), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n637), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n610), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n658), .A3(new_n448), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n799), .A2(new_n376), .A3(new_n486), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n299), .B1(new_n800), .B2(new_n637), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n486), .A2(new_n376), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n798), .A2(new_n470), .A3(new_n444), .A4(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n803), .A2(new_n302), .A3(new_n796), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n801), .A2(new_n804), .ZN(G1340gat));
  AOI21_X1  g604(.A(new_n303), .B1(new_n800), .B2(new_n607), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n803), .A2(G120gat), .A3(new_n608), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n806), .A2(new_n807), .ZN(G1341gat));
  NAND3_X1  g607(.A1(new_n800), .A2(G127gat), .A3(new_n668), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n308), .B1(new_n803), .B2(new_n589), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT119), .ZN(G1342gat));
  NOR3_X1   g611(.A1(new_n803), .A2(G134gat), .A3(new_n557), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT56), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n800), .A2(new_n558), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n815), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT120), .B1(new_n815), .B2(G134gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(G1343gat));
  NOR2_X1   g617(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n819));
  AND2_X1   g618(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n820));
  INV_X1    g619(.A(new_n794), .ZN(new_n821));
  INV_X1    g620(.A(new_n790), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n781), .B1(new_n634), .B2(new_n636), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n783), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n821), .B1(new_n824), .B2(new_n558), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n825), .A2(new_n589), .B1(new_n610), .B2(new_n796), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT57), .B1(new_n826), .B2(new_n658), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n798), .A2(new_n828), .A3(new_n711), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n802), .A2(new_n449), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT121), .Z(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G141gat), .B1(new_n832), .B2(new_n796), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n798), .A2(new_n711), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n830), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n637), .A2(new_n331), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT122), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI211_X1 g637(.A(new_n819), .B(new_n820), .C1(new_n833), .C2(new_n838), .ZN(new_n839));
  AND4_X1   g638(.A1(KEYINPUT123), .A2(new_n833), .A3(KEYINPUT58), .A4(new_n838), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(G1344gat));
  AOI211_X1 g640(.A(new_n828), .B(new_n470), .C1(new_n795), .C2(new_n797), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n828), .B1(new_n826), .B2(new_n658), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(KEYINPUT124), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n842), .A2(KEYINPUT124), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n607), .B(new_n831), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n847));
  NOR4_X1   g646(.A1(new_n834), .A2(new_n333), .A3(new_n608), .A4(new_n830), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n333), .B1(new_n832), .B2(new_n608), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(G1345gat));
  NAND2_X1  g651(.A1(new_n326), .A2(new_n328), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n832), .A2(new_n853), .A3(new_n775), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n740), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n853), .B2(new_n855), .ZN(G1346gat));
  AOI21_X1  g655(.A(G162gat), .B1(new_n835), .B2(new_n558), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n832), .A2(new_n557), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(G162gat), .ZN(G1347gat));
  AOI21_X1  g658(.A(new_n671), .B1(new_n795), .B2(new_n797), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n498), .A2(new_n496), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT125), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n235), .A3(new_n637), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n498), .A2(new_n671), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n799), .A2(KEYINPUT126), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT126), .B1(new_n799), .B2(new_n866), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(new_n637), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n864), .B1(new_n870), .B2(new_n235), .ZN(G1348gat));
  AOI21_X1  g670(.A(G176gat), .B1(new_n863), .B2(new_n607), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n869), .A2(new_n607), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(G176gat), .ZN(G1349gat));
  NAND3_X1  g673(.A1(new_n867), .A2(new_n668), .A3(new_n868), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G183gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n863), .A2(new_n740), .A3(new_n230), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT60), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n876), .A2(new_n880), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1350gat));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n217), .A3(new_n558), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n558), .A3(new_n868), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(G190gat), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n884), .B2(G190gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(G1351gat));
  AND4_X1   g687(.A1(new_n486), .A2(new_n860), .A3(new_n711), .A4(new_n449), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n629), .A3(new_n637), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n844), .A2(new_n845), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n866), .A2(new_n697), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n891), .A2(new_n796), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(new_n894), .B2(new_n629), .ZN(G1352gat));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT127), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n889), .B1(KEYINPUT127), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n608), .A2(G204gat), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n889), .A2(KEYINPUT127), .A3(new_n896), .A4(new_n899), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n891), .A2(new_n608), .A3(new_n893), .ZN(new_n903));
  INV_X1    g702(.A(G204gat), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(G1353gat));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n202), .A3(new_n740), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n740), .B(new_n892), .C1(new_n844), .C2(new_n845), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n907), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT63), .B1(new_n907), .B2(G211gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(G1354gat));
  NAND3_X1  g709(.A1(new_n889), .A2(new_n203), .A3(new_n558), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n891), .A2(new_n557), .A3(new_n893), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n203), .ZN(G1355gat));
endmodule


