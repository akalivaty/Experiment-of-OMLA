//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  NOR2_X1   g0009(.A1(G97), .A2(G107), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G87), .ZN(G355));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n202), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n213), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n206), .A2(new_n207), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n213), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(G250), .B1(G257), .B2(G264), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n232), .A2(KEYINPUT0), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(KEYINPUT0), .ZN(new_n234));
  NAND4_X1  g0034(.A1(new_n223), .A2(new_n228), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n222), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n215), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT66), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n253), .A2(KEYINPUT66), .A3(G13), .A4(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n225), .B1(new_n213), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n253), .A2(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(G50), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G50), .B2(new_n258), .ZN(new_n265));
  INV_X1    g0065(.A(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n208), .A2(G20), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n226), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n269), .A2(new_n271), .B1(G150), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n266), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G222), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(G223), .A3(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n278), .B(new_n279), .C1(new_n280), .C2(new_n276), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n286), .B1(G226), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n275), .B1(G169), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n292), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G179), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(G190), .ZN(new_n297));
  XOR2_X1   g0097(.A(new_n297), .B(KEYINPUT69), .Z(new_n298));
  NAND2_X1  g0098(.A1(new_n275), .A2(KEYINPUT9), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n265), .A2(KEYINPUT9), .A3(new_n274), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n294), .A2(G200), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n298), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n298), .A2(new_n301), .A3(new_n305), .A4(new_n302), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n296), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT68), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n256), .A2(new_n309), .A3(new_n257), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n311), .A2(G68), .A3(new_n266), .A4(new_n263), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n271), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n313));
  INV_X1    g0113(.A(new_n272), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n207), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n261), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT11), .ZN(new_n317));
  INV_X1    g0117(.A(new_n310), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n309), .B1(new_n256), .B2(new_n257), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT12), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n258), .B2(G68), .ZN(new_n323));
  AND4_X1   g0123(.A1(new_n312), .A2(new_n317), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n328), .A2(new_n215), .A3(new_n277), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n325), .A2(new_n327), .A3(G226), .A4(new_n277), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n282), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n288), .A2(G274), .ZN(new_n334));
  INV_X1    g0134(.A(new_n285), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n290), .A2(G238), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT13), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n333), .B2(new_n336), .ZN(new_n339));
  OAI21_X1  g0139(.A(G200), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n333), .A2(new_n336), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT13), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(G190), .A3(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n324), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n342), .B2(new_n343), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT71), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(G169), .C1(new_n338), .C2(new_n339), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n338), .A2(new_n339), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(KEYINPUT71), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT70), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT14), .B1(new_n347), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n355), .B(G169), .C1(new_n338), .C2(new_n339), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n350), .B(new_n354), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n324), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n345), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n276), .A2(G232), .A3(new_n277), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n276), .A2(G238), .A3(G1698), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n328), .A2(G107), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n282), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n286), .B1(G244), .B2(new_n290), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT67), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n366), .B2(new_n367), .ZN(new_n371));
  OAI21_X1  g0171(.A(G190), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n366), .A2(new_n367), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT67), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(G200), .A3(new_n369), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n311), .A2(G77), .A3(new_n266), .A4(new_n263), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n268), .A2(new_n314), .B1(new_n226), .B2(new_n280), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT15), .B(G87), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n270), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n261), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n320), .A2(new_n280), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n376), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n372), .A2(new_n375), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n374), .A2(new_n369), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n384), .B2(new_n352), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n374), .A2(new_n346), .A3(new_n369), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n307), .A2(new_n361), .A3(new_n383), .A4(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n268), .B1(new_n253), .B2(G20), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n262), .A2(new_n389), .B1(new_n259), .B2(new_n268), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n276), .A2(G226), .A3(G1698), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n276), .A2(G223), .A3(new_n277), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n282), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n335), .A2(new_n288), .A3(G274), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n215), .B2(new_n289), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G190), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n399), .A2(KEYINPUT74), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(KEYINPUT74), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n395), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n397), .B1(new_n394), .B2(new_n282), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(G200), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G58), .A2(G68), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n204), .A2(new_n205), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G20), .ZN(new_n408));
  INV_X1    g0208(.A(G159), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n409), .A2(G20), .A3(G33), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT72), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(KEYINPUT72), .A3(new_n411), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT7), .B1(new_n328), .B2(new_n226), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n417), .B(G20), .C1(new_n325), .C2(new_n327), .ZN(new_n418));
  OAI21_X1  g0218(.A(G68), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n415), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n261), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT72), .B1(new_n408), .B2(new_n411), .ZN(new_n422));
  AOI211_X1 g0222(.A(new_n413), .B(new_n410), .C1(new_n407), .C2(G20), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT16), .B1(new_n424), .B2(new_n419), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n390), .B(new_n405), .C1(new_n421), .C2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT17), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n390), .B1(new_n421), .B2(new_n425), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n395), .A2(new_n352), .A3(new_n398), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G169), .B2(new_n404), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT18), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT73), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n428), .A2(KEYINPUT18), .A3(new_n431), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n428), .A2(new_n431), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n427), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n388), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n288), .A2(G274), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G1), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(G270), .A3(new_n288), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT80), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n328), .A2(G303), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n325), .A2(new_n327), .A3(G264), .A4(G1698), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n325), .A2(new_n327), .A3(G257), .A4(new_n277), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT79), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT79), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n453), .A2(new_n458), .A3(new_n454), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n452), .B1(new_n460), .B2(new_n282), .ZN(new_n461));
  AOI211_X1 g0261(.A(KEYINPUT80), .B(new_n288), .C1(new_n457), .C2(new_n459), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n451), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n226), .C1(G33), .C2(new_n216), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(G20), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(new_n261), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n320), .A2(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n464), .B1(new_n253), .B2(G33), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n266), .B(new_n473), .C1(new_n318), .C2(new_n319), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n346), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT21), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n463), .A2(new_n478), .A3(new_n475), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT81), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n461), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n470), .A2(new_n471), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(new_n474), .C1(G116), .C2(new_n311), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n449), .A2(G179), .A3(new_n450), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n480), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n484), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n472), .B2(new_n474), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(KEYINPUT81), .C1(new_n462), .C2(new_n461), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n477), .A2(new_n479), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n463), .A2(G200), .ZN(new_n491));
  INV_X1    g0291(.A(new_n483), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n491), .B(new_n492), .C1(new_n402), .C2(new_n463), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n325), .A2(new_n327), .A3(new_n226), .A4(G87), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n495), .B(KEYINPUT22), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT83), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT23), .B1(new_n226), .B2(G107), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT23), .ZN(new_n500));
  INV_X1    g0300(.A(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n501), .A3(G20), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n499), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT82), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT82), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n499), .A2(new_n502), .A3(new_n503), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT83), .B2(KEYINPUT24), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n261), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n258), .A2(G107), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n514), .B(KEYINPUT25), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n253), .A2(G33), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n258), .A2(new_n266), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G107), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT84), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n448), .A2(new_n288), .ZN(new_n522));
  INV_X1    g0322(.A(G264), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n448), .A2(KEYINPUT84), .A3(G264), .A4(new_n288), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n276), .A2(G257), .A3(G1698), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n276), .A2(G250), .A3(new_n277), .ZN(new_n528));
  INV_X1    g0328(.A(G294), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n527), .B(new_n528), .C1(new_n260), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n282), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n526), .A2(new_n531), .A3(G190), .A4(new_n449), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n526), .A2(new_n531), .A3(new_n449), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G200), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n513), .A2(new_n520), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT76), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT6), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G97), .A2(G107), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n540), .B2(new_n210), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT75), .ZN(new_n542));
  MUX2_X1   g0342(.A(new_n542), .B(G97), .S(KEYINPUT6), .Z(new_n543));
  NAND2_X1  g0343(.A1(new_n211), .A2(new_n539), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n536), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n538), .B1(new_n537), .B2(G97), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(new_n211), .A3(new_n539), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n536), .B1(new_n548), .B2(new_n541), .ZN(new_n549));
  OAI21_X1  g0349(.A(G20), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n417), .B1(new_n276), .B2(G20), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n326), .A2(G33), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n553));
  OAI211_X1 g0353(.A(KEYINPUT7), .B(new_n226), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(G107), .B1(G77), .B2(new_n272), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n261), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n325), .A2(new_n327), .A3(G244), .A4(new_n277), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT77), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n276), .A2(G244), .A3(new_n277), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n562), .A2(new_n465), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n282), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n448), .A2(G257), .A3(new_n288), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n449), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G200), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n258), .A2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n517), .B2(G97), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n567), .A2(G190), .A3(new_n569), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n558), .A2(new_n571), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n346), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(new_n352), .A3(new_n569), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n266), .B1(new_n550), .B2(new_n556), .ZN(new_n578));
  INV_X1    g0378(.A(new_n573), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n535), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n276), .A2(new_n226), .A3(G68), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n226), .B1(new_n331), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(G87), .B2(new_n211), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n270), .B2(new_n216), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n261), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n308), .A2(new_n310), .A3(new_n378), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n258), .A2(new_n266), .A3(G87), .A4(new_n516), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n288), .A2(G274), .A3(new_n445), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n253), .A2(G45), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n288), .A2(G250), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n325), .A2(new_n327), .A3(G238), .A4(new_n277), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n325), .A2(new_n327), .A3(G244), .A4(G1698), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n598), .C1(new_n260), .C2(new_n464), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(new_n282), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G190), .ZN(new_n601));
  INV_X1    g0401(.A(G200), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n592), .B(new_n601), .C1(new_n602), .C2(new_n600), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n352), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT78), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n600), .A2(G169), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n600), .A2(KEYINPUT78), .A3(new_n352), .ZN(new_n608));
  INV_X1    g0408(.A(new_n378), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n517), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n588), .A3(new_n589), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n512), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n509), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n519), .B1(new_n614), .B2(new_n261), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n533), .A2(new_n346), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(G179), .B2(new_n533), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n603), .B(new_n612), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  NOR4_X1   g0418(.A1(new_n442), .A2(new_n494), .A3(new_n581), .A4(new_n618), .ZN(G372));
  INV_X1    g0419(.A(new_n390), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n203), .B1(new_n551), .B2(new_n554), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT16), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n266), .B1(new_n424), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n622), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n620), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n437), .B1(new_n627), .B2(new_n430), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n434), .ZN(new_n629));
  INV_X1    g0429(.A(new_n345), .ZN(new_n630));
  INV_X1    g0430(.A(new_n387), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n359), .A2(new_n360), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT17), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n426), .B(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n629), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n304), .A2(new_n306), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n296), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n486), .A2(new_n489), .ZN(new_n640));
  INV_X1    g0440(.A(new_n617), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n513), .A2(new_n520), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n478), .B1(new_n463), .B2(new_n475), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n463), .A2(new_n478), .A3(new_n475), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n640), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT85), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n592), .B(new_n647), .C1(new_n602), .C2(new_n600), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n600), .A2(new_n602), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT85), .B1(new_n649), .B2(new_n591), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n601), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n581), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n607), .A2(new_n611), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n604), .ZN(new_n656));
  INV_X1    g0456(.A(new_n580), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n656), .A3(new_n651), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n603), .A4(new_n612), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n654), .A2(new_n656), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n639), .B1(new_n442), .B2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(new_n490), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n253), .A2(new_n226), .A3(G13), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n492), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n494), .B2(new_n674), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n535), .B1(new_n615), .B2(new_n673), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n643), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n641), .A2(new_n642), .A3(new_n673), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n490), .A2(new_n672), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n685), .B(KEYINPUT86), .Z(G399));
  NOR2_X1   g0486(.A1(new_n230), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n211), .A2(G87), .A3(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n224), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n688), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  AND4_X1   g0493(.A1(new_n484), .A2(new_n526), .A3(new_n531), .A4(new_n600), .ZN(new_n694));
  INV_X1    g0494(.A(new_n570), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n694), .B(new_n695), .C1(new_n462), .C2(new_n461), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n600), .A2(G179), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n570), .A2(new_n533), .A3(new_n698), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n696), .A2(new_n697), .B1(new_n463), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT87), .B1(new_n696), .B2(new_n697), .ZN(new_n701));
  INV_X1    g0501(.A(new_n481), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT87), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n484), .A2(new_n526), .A3(new_n531), .A4(new_n600), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n570), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(KEYINPUT30), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n700), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n672), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n618), .A2(new_n581), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n490), .A3(new_n493), .A4(new_n673), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT88), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT88), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(G330), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n646), .A2(new_n653), .B1(new_n604), .B2(new_n655), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n672), .B1(new_n720), .B2(new_n662), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n603), .A2(new_n612), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n724), .A2(new_n580), .A3(KEYINPUT26), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(KEYINPUT26), .B2(new_n658), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n672), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n723), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n719), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n693), .B1(new_n729), .B2(G1), .ZN(G364));
  INV_X1    g0530(.A(G13), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n731), .A2(new_n444), .A3(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n253), .B1(new_n732), .B2(KEYINPUT89), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(KEYINPUT89), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n687), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n677), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n676), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n735), .B(KEYINPUT90), .ZN(new_n738));
  INV_X1    g0538(.A(G355), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n276), .A2(new_n229), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n739), .A2(new_n740), .B1(G116), .B2(new_n229), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n248), .A2(new_n444), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n230), .A2(new_n276), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n224), .B2(new_n444), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n741), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n225), .B1(G20), .B2(new_n346), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n738), .B1(new_n746), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n402), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n226), .A2(new_n352), .A3(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n399), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n226), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n756), .A2(new_n757), .B1(new_n529), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n755), .A2(new_n399), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(G311), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n602), .A2(G179), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(G20), .A3(G190), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n276), .B1(new_n766), .B2(G303), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n226), .A2(G190), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(new_n352), .A3(new_n602), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(new_n768), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G329), .A2(new_n770), .B1(new_n772), .B2(G283), .ZN(new_n773));
  NAND3_X1  g0573(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT91), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G190), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n775), .A2(new_n402), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(G326), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n763), .A2(new_n767), .A3(new_n773), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n770), .A2(G159), .ZN(new_n781));
  XOR2_X1   g0581(.A(KEYINPUT92), .B(KEYINPUT32), .Z(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n782), .B1(new_n759), .B2(new_n216), .ZN(new_n783));
  INV_X1    g0583(.A(G87), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n765), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n276), .B1(new_n771), .B2(new_n501), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n756), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n788), .A2(G58), .B1(new_n781), .B2(new_n782), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n787), .B(new_n789), .C1(new_n280), .C2(new_n761), .ZN(new_n790));
  INV_X1    g0590(.A(new_n778), .ZN(new_n791));
  INV_X1    g0591(.A(new_n776), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n207), .A2(new_n791), .B1(new_n792), .B2(new_n203), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n780), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT93), .ZN(new_n795));
  INV_X1    g0595(.A(new_n750), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n794), .B2(KEYINPUT93), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n753), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n749), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n676), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n737), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT94), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n796), .A2(new_n748), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n738), .B1(G77), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT95), .Z(new_n806));
  AOI21_X1  g0606(.A(new_n276), .B1(new_n770), .B2(G311), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n761), .A2(new_n464), .B1(new_n759), .B2(new_n216), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n788), .B2(G294), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n766), .A2(G107), .B1(new_n772), .B2(G87), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n776), .A2(G283), .B1(new_n778), .B2(G303), .ZN(new_n811));
  AND4_X1   g0611(.A1(new_n807), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n788), .A2(G143), .B1(G159), .B2(new_n762), .ZN(new_n813));
  INV_X1    g0613(.A(G150), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n792), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G137), .B2(new_n778), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT34), .Z(new_n817));
  OAI21_X1  g0617(.A(new_n276), .B1(new_n765), .B2(new_n207), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n772), .A2(G68), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n820), .B2(new_n769), .ZN(new_n821));
  INV_X1    g0621(.A(new_n759), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n818), .B(new_n821), .C1(G58), .C2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n812), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT96), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n385), .A2(new_n386), .A3(new_n673), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n382), .A2(new_n673), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n383), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n825), .B(new_n826), .C1(new_n631), .C2(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n383), .A2(new_n827), .B1(new_n385), .B2(new_n386), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n385), .A2(new_n386), .A3(new_n673), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT96), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n806), .B1(new_n824), .B2(new_n796), .C1(new_n833), .C2(new_n748), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT97), .B1(new_n721), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n721), .A2(new_n833), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n835), .B(new_n836), .Z(new_n837));
  OAI22_X1  g0637(.A1(new_n837), .A2(new_n719), .B1(new_n687), .B2(new_n734), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n837), .A2(new_n719), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n834), .B1(new_n838), .B2(new_n839), .ZN(G384));
  AOI21_X1  g0640(.A(new_n253), .B1(G13), .B2(new_n226), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT40), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n426), .B1(new_n627), .B2(new_n430), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n627), .A2(new_n670), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n670), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n428), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT37), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n436), .A2(new_n847), .A3(new_n848), .A4(new_n426), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n422), .A2(new_n423), .A3(new_n621), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n261), .B(new_n420), .C1(new_n852), .C2(KEYINPUT16), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n437), .B(new_n430), .C1(new_n853), .C2(new_n390), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n628), .B1(new_n854), .B2(KEYINPUT73), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n438), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n847), .B1(new_n856), .B2(new_n427), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n851), .B1(new_n857), .B2(KEYINPUT99), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT99), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n636), .B1(new_n855), .B2(new_n438), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n860), .B2(new_n847), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n440), .A2(KEYINPUT99), .A3(new_n844), .ZN(new_n863));
  AND4_X1   g0663(.A1(KEYINPUT38), .A2(new_n861), .A3(new_n863), .A4(new_n850), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n360), .A2(new_n672), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n633), .A2(new_n630), .A3(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n360), .B(new_n672), .C1(new_n345), .C2(new_n359), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n867), .A2(new_n868), .B1(new_n829), .B2(new_n832), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n714), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT102), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT102), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n714), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n842), .B1(new_n865), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n714), .A2(new_n869), .A3(KEYINPUT40), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n847), .B1(new_n427), .B2(new_n629), .ZN(new_n877));
  INV_X1    g0677(.A(new_n843), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(KEYINPUT100), .A3(new_n848), .A4(new_n847), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT100), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n849), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(new_n881), .A3(new_n845), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n877), .B1(new_n882), .B2(KEYINPUT101), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT101), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n879), .A2(new_n881), .A3(new_n884), .A4(new_n845), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n876), .B1(new_n864), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n875), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n441), .A2(new_n714), .ZN(new_n889));
  OAI21_X1  g0689(.A(G330), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT103), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n892), .B(new_n893), .C1(new_n888), .C2(new_n889), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n864), .B2(new_n886), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n861), .A2(new_n863), .A3(new_n850), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n861), .A2(new_n863), .A3(KEYINPUT38), .A4(new_n850), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n633), .A2(new_n672), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n897), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n629), .A2(new_n846), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n900), .A2(new_n901), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n831), .B1(new_n721), .B2(new_n833), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n867), .A2(new_n868), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n905), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n728), .A2(new_n441), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n639), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n912), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n841), .B1(new_n895), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n895), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n546), .A2(new_n549), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT98), .Z(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT35), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(KEYINPUT35), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(G116), .A4(new_n227), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT36), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n224), .A2(G77), .A3(new_n406), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(G50), .B2(new_n203), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(G1), .A3(new_n731), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n917), .A2(new_n924), .A3(new_n927), .ZN(G367));
  NAND2_X1  g0728(.A1(new_n244), .A2(new_n743), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n751), .C1(new_n229), .C2(new_n378), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n738), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n591), .A2(new_n672), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n651), .A2(new_n656), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n656), .B2(new_n932), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n756), .A2(new_n814), .B1(new_n203), .B2(new_n759), .ZN(new_n935));
  AOI22_X1  g0735(.A1(G58), .A2(new_n766), .B1(new_n770), .B2(G137), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(new_n276), .C1(new_n280), .C2(new_n771), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n935), .B(new_n937), .C1(G143), .C2(new_n778), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT107), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n792), .A2(new_n409), .B1(new_n207), .B2(new_n761), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT108), .Z(new_n943));
  NAND3_X1  g0743(.A1(new_n766), .A2(KEYINPUT46), .A3(G116), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT46), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n765), .B2(new_n464), .ZN(new_n946));
  INV_X1    g0746(.A(G283), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n944), .B(new_n946), .C1(new_n947), .C2(new_n761), .ZN(new_n948));
  INV_X1    g0748(.A(G303), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n756), .A2(new_n949), .B1(new_n501), .B2(new_n759), .ZN(new_n950));
  INV_X1    g0750(.A(G317), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n328), .B1(new_n771), .B2(new_n216), .C1(new_n951), .C2(new_n769), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n948), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n776), .A2(G294), .B1(new_n778), .B2(G311), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n943), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT47), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n931), .B1(new_n799), .B2(new_n934), .C1(new_n956), .C2(new_n796), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n734), .B(KEYINPUT106), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n657), .A2(new_n672), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n672), .B1(new_n578), .B2(new_n579), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n575), .A2(new_n580), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n684), .B2(new_n680), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT44), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n684), .A2(new_n680), .A3(new_n962), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n682), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n964), .A2(new_n682), .A3(new_n967), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n970), .A2(new_n971), .B1(KEYINPUT105), .B2(new_n968), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(KEYINPUT105), .A3(new_n682), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n681), .B(new_n683), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n677), .B(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n729), .A3(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n729), .ZN(new_n978));
  XOR2_X1   g0778(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n979));
  XNOR2_X1  g0779(.A(new_n687), .B(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n958), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n681), .A2(new_n683), .A3(new_n962), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n580), .B1(new_n961), .B2(new_n643), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n983), .A2(KEYINPUT42), .B1(new_n673), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n984), .A2(new_n986), .B1(KEYINPUT43), .B2(new_n934), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n987), .B(new_n988), .Z(new_n989));
  INV_X1    g0789(.A(new_n962), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n682), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n989), .B(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n957), .B1(new_n982), .B2(new_n993), .ZN(G387));
  NAND2_X1  g0794(.A1(new_n975), .A2(new_n958), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT109), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n689), .A2(new_n740), .B1(G107), .B2(new_n229), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n241), .A2(new_n444), .ZN(new_n998));
  INV_X1    g0798(.A(new_n689), .ZN(new_n999));
  AOI211_X1 g0799(.A(G45), .B(new_n999), .C1(G68), .C2(G77), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n268), .A2(G50), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n744), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n997), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n738), .B1(new_n1004), .B2(new_n752), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n822), .A2(new_n609), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n203), .B2(new_n761), .C1(new_n756), .C2(new_n207), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n276), .B1(new_n771), .B2(new_n216), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n765), .A2(new_n280), .B1(new_n769), .B2(new_n814), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n409), .B2(new_n791), .C1(new_n268), .C2(new_n792), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n276), .B1(new_n770), .B2(G326), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n759), .A2(new_n947), .B1(new_n765), .B2(new_n529), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n788), .A2(G317), .B1(G303), .B2(new_n762), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n776), .A2(G311), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n757), .C2(new_n791), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1012), .B1(new_n464), .B2(new_n771), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1011), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1005), .B1(new_n1023), .B2(new_n750), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n681), .B2(new_n799), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT110), .Z(new_n1026));
  NOR2_X1   g0826(.A1(new_n729), .A2(new_n975), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n729), .A2(new_n975), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n687), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n996), .B(new_n1026), .C1(new_n1027), .C2(new_n1029), .ZN(G393));
  NAND2_X1  g0830(.A1(new_n970), .A2(new_n971), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n688), .B1(new_n1031), .B2(new_n1028), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n977), .A2(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n751), .B1(new_n216), .B2(new_n229), .C1(new_n251), .C2(new_n744), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n738), .A2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n788), .A2(G311), .B1(G317), .B2(new_n778), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n792), .A2(new_n949), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n276), .B1(new_n772), .B2(G107), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n947), .B2(new_n765), .C1(new_n757), .C2(new_n769), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n761), .A2(new_n529), .B1(new_n759), .B2(new_n464), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT111), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT111), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n759), .A2(new_n280), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G68), .A2(new_n766), .B1(new_n770), .B2(G143), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n276), .C1(new_n784), .C2(new_n771), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1045), .B(new_n1047), .C1(new_n269), .C2(new_n762), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n791), .A2(new_n814), .B1(new_n409), .B2(new_n756), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT51), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(new_n207), .C2(new_n792), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1043), .A2(new_n1044), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1035), .B1(new_n1052), .B2(new_n750), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n799), .B2(new_n962), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n958), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n1031), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1033), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(G390));
  NAND3_X1  g0858(.A1(new_n663), .A2(new_n673), .A3(new_n833), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n826), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n903), .B1(new_n1060), .B2(new_n908), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n901), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n845), .B1(new_n880), .B2(new_n849), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n849), .A2(new_n880), .ZN(new_n1065));
  OAI21_X1  g0865(.A(KEYINPUT101), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n877), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n885), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n899), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT39), .B1(new_n1069), .B2(new_n901), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1062), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n901), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n654), .A2(new_n656), .A3(new_n726), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n673), .A3(new_n833), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n826), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT112), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n908), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n867), .A2(KEYINPUT112), .A3(new_n868), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n903), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1072), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n716), .A2(new_n718), .A3(new_n833), .A4(new_n908), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1071), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n833), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n715), .A2(new_n1085), .A3(new_n909), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1061), .B1(new_n897), .B2(new_n902), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1072), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1084), .A2(new_n1089), .A3(new_n958), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n748), .B1(new_n897), .B2(new_n902), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n792), .A2(new_n501), .B1(new_n216), .B2(new_n761), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1092), .A2(KEYINPUT115), .B1(G283), .B2(new_n778), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(KEYINPUT115), .B2(new_n1092), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT116), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n819), .B1(new_n529), .B2(new_n769), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1096), .A2(new_n276), .A3(new_n785), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1045), .B1(new_n788), .B2(G116), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(G125), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n276), .B1(new_n771), .B2(new_n207), .C1(new_n1100), .C2(new_n769), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n765), .A2(new_n814), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT54), .B(G143), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1103), .B1(new_n409), .B2(new_n759), .C1(new_n761), .C2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1101), .B(new_n1105), .C1(G137), .C2(new_n776), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n788), .A2(G132), .B1(G128), .B2(new_n778), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT114), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n796), .B1(new_n1099), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n738), .B1(new_n269), .B2(new_n804), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n1091), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1090), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1079), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1085), .B2(new_n715), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1075), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1083), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n716), .A2(new_n718), .A3(new_n833), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1086), .B1(new_n1120), .B2(new_n909), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1121), .B2(new_n907), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n442), .A2(new_n715), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n914), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1115), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1084), .A2(new_n1089), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1127));
  AND4_X1   g0927(.A1(KEYINPUT113), .A2(new_n1126), .A3(new_n687), .A4(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n688), .B1(new_n1115), .B2(new_n1125), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT113), .B1(new_n1129), .B2(new_n1127), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1114), .B1(new_n1128), .B2(new_n1130), .ZN(G378));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1127), .A2(new_n1124), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n873), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n872), .B1(new_n714), .B2(new_n869), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT40), .B1(new_n1136), .B2(new_n906), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n887), .A2(G330), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n307), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n275), .A2(new_n846), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT117), .Z(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n307), .A2(new_n1140), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1142), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n307), .A2(new_n1140), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1144), .B1(new_n1148), .B2(new_n1141), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1137), .A2(new_n1138), .A3(new_n1150), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1152));
  INV_X1    g0952(.A(G330), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n1072), .B2(new_n876), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1152), .B1(new_n875), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n912), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1150), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n875), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n904), .A4(new_n911), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1132), .B1(new_n1133), .B2(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1127), .A2(new_n1124), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(KEYINPUT57), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n687), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1156), .A2(new_n958), .A3(new_n1159), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n735), .B1(G50), .B2(new_n804), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(G33), .A2(G41), .ZN(new_n1168));
  INV_X1    g0968(.A(G41), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G50), .B(new_n1168), .C1(new_n328), .C2(new_n1169), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n761), .A2(new_n378), .B1(new_n759), .B2(new_n203), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n788), .B2(G107), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n776), .A2(G97), .B1(new_n778), .B2(G116), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G41), .B(new_n276), .C1(new_n766), .C2(G77), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G283), .A2(new_n770), .B1(new_n772), .B2(G58), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1170), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n759), .A2(new_n814), .B1(new_n765), .B2(new_n1104), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n762), .A2(G137), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G128), .C2(new_n788), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n1100), .B2(new_n791), .C1(new_n820), .C2(new_n792), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1168), .B1(new_n771), .B2(new_n409), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G124), .B2(new_n770), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1178), .B1(new_n1177), .B2(new_n1176), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1167), .B1(new_n1188), .B2(new_n750), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n1150), .B2(new_n748), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT118), .Z(new_n1191));
  NAND2_X1  g0991(.A1(new_n1166), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1165), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(G375));
  OR2_X1    g0995(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(new_n981), .A3(new_n1125), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n788), .A2(G137), .B1(G50), .B2(new_n822), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n814), .B2(new_n761), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G128), .A2(new_n770), .B1(new_n766), .B2(G159), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1200), .B(new_n276), .C1(new_n202), .C2(new_n771), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n820), .A2(new_n791), .B1(new_n792), .B2(new_n1104), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n464), .A2(new_n792), .B1(new_n791), .B2(new_n529), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1006), .B1(new_n501), .B2(new_n761), .C1(new_n756), .C2(new_n947), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n276), .B1(new_n772), .B2(G77), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n216), .B2(new_n765), .C1(new_n949), .C2(new_n769), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n750), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1209), .B(new_n738), .C1(G68), .C2(new_n804), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1116), .B2(new_n747), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1122), .B2(new_n958), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1197), .A2(new_n1212), .ZN(G381));
  NOR3_X1   g1013(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT119), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1057), .B(new_n957), .C1(new_n982), .C2(new_n993), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1129), .A2(new_n1127), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(new_n1113), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1215), .A2(new_n1216), .A3(G381), .A4(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1220), .A2(KEYINPUT120), .A3(new_n1194), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT120), .B1(new_n1220), .B2(new_n1194), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1221), .A2(new_n1222), .ZN(G407));
  NAND3_X1  g1023(.A1(new_n1194), .A2(new_n671), .A3(new_n1218), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(G407), .A2(G213), .A3(new_n1224), .ZN(G409));
  INV_X1    g1025(.A(KEYINPUT61), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1125), .A2(KEYINPUT60), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(new_n1196), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n687), .B1(new_n1227), .B2(new_n1196), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1212), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(G384), .ZN(new_n1231));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(G343), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(G2897), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1231), .B(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1165), .A2(G378), .A3(new_n1193), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT121), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1192), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1166), .A2(KEYINPUT121), .A3(new_n1191), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1162), .A2(new_n981), .A3(new_n1163), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1218), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1233), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1226), .B1(new_n1235), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1236), .A2(new_n1242), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1233), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1231), .A3(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1249), .A2(KEYINPUT63), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G387), .A2(G390), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT122), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1216), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(new_n802), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1251), .A2(new_n1254), .A3(new_n1252), .A4(new_n1216), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1249), .A2(KEYINPUT63), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1245), .A2(new_n1250), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT124), .ZN(new_n1261));
  XOR2_X1   g1061(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n1262));
  AOI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n1243), .C2(new_n1231), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1262), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT124), .B1(new_n1248), .B2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1246), .A2(KEYINPUT62), .A3(new_n1231), .A4(new_n1247), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT125), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1243), .A2(KEYINPUT125), .A3(KEYINPUT62), .A4(new_n1231), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1244), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1258), .B(KEYINPUT126), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1260), .B1(new_n1272), .B2(new_n1273), .ZN(G405));
  OAI21_X1  g1074(.A(new_n1236), .B1(new_n1194), .B2(new_n1219), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(new_n1231), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1258), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1256), .A2(KEYINPUT127), .A3(new_n1257), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1278), .B2(new_n1276), .ZN(G402));
endmodule


