//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1208, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n202), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n212), .B(new_n218), .C1(G107), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n210), .B(new_n227), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n221), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(G33), .A2(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n250), .B1(G232), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G226), .A2(G1698), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n255), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n258), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n256), .B(new_n260), .C1(new_n223), .C2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(KEYINPUT13), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(KEYINPUT69), .A3(G169), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT14), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(G179), .A3(new_n265), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n228), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n274), .A2(new_n202), .B1(new_n229), .B2(G68), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n229), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n272), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT11), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n272), .B1(new_n257), .B2(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT12), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(new_n229), .A3(G1), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n283), .B1(new_n285), .B2(new_n222), .ZN(new_n286));
  INV_X1    g0086(.A(new_n285), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(KEYINPUT12), .A3(G68), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n280), .B1(new_n222), .B2(new_n282), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT70), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n270), .B(new_n290), .C1(new_n268), .C2(new_n267), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n266), .B2(G200), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n266), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g0095(.A(new_n295), .B(KEYINPUT71), .Z(new_n296));
  INV_X1    g0096(.A(KEYINPUT18), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT72), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT3), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(new_n301), .A3(G33), .ZN(new_n302));
  INV_X1    g0102(.A(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G223), .B2(G1698), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n251), .A2(G226), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n306), .A2(new_n307), .B1(new_n303), .B2(new_n214), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n255), .ZN(new_n309));
  INV_X1    g0109(.A(new_n262), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G232), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n260), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G169), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n309), .A2(G179), .A3(new_n260), .A4(new_n311), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT66), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n282), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n318), .B1(new_n285), .B2(new_n317), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT16), .ZN(new_n320));
  AND3_X1   g0120(.A1(KEYINPUT74), .A2(G58), .A3(G68), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT74), .B1(G58), .B2(G68), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n321), .A2(new_n322), .A3(new_n201), .ZN(new_n323));
  INV_X1    g0123(.A(G159), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n323), .A2(new_n229), .B1(new_n324), .B2(new_n274), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n302), .A2(new_n229), .A3(new_n304), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT7), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT7), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n302), .A2(new_n328), .A3(new_n229), .A4(new_n304), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(G68), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT73), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n327), .A2(KEYINPUT73), .A3(G68), .A4(new_n329), .ZN(new_n333));
  AOI211_X1 g0133(.A(new_n320), .B(new_n325), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n328), .B1(new_n250), .B2(G20), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT72), .B(KEYINPUT3), .ZN(new_n336));
  OAI211_X1 g0136(.A(KEYINPUT7), .B(new_n229), .C1(new_n336), .C2(G33), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n298), .A2(new_n303), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n325), .B1(new_n339), .B2(G68), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n272), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n341));
  OAI211_X1 g0141(.A(KEYINPUT75), .B(new_n319), .C1(new_n334), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n332), .A2(new_n333), .ZN(new_n344));
  INV_X1    g0144(.A(new_n325), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(KEYINPUT16), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n341), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT75), .B1(new_n348), .B2(new_n319), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n315), .B1(new_n343), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n297), .B1(new_n350), .B2(KEYINPUT76), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT77), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n350), .B2(KEYINPUT76), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n313), .A2(new_n314), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT75), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n325), .B1(new_n332), .B2(new_n333), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n341), .B1(new_n356), .B2(KEYINPUT16), .ZN(new_n357));
  INV_X1    g0157(.A(new_n319), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n354), .B1(new_n359), .B2(new_n342), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT77), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n351), .B1(new_n353), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n312), .A2(G200), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n348), .A2(new_n319), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n312), .A2(new_n293), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT17), .ZN(new_n368));
  INV_X1    g0168(.A(new_n366), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n369), .A2(new_n348), .A3(new_n319), .A4(new_n364), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT17), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n350), .A2(KEYINPUT76), .A3(new_n352), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT77), .B1(new_n360), .B2(new_n361), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT18), .B1(new_n360), .B2(new_n361), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n363), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n296), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n203), .A2(G20), .ZN(new_n380));
  INV_X1    g0180(.A(G150), .ZN(new_n381));
  OAI221_X1 g0181(.A(new_n380), .B1(new_n381), .B2(new_n274), .C1(new_n317), .C2(new_n276), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n272), .B1(new_n202), .B2(new_n285), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n202), .B2(new_n282), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT9), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G222), .A2(G1698), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n251), .A2(G223), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n250), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n255), .C1(G77), .C2(new_n250), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n389), .B(new_n260), .C1(new_n211), .C2(new_n262), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G200), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n385), .B(new_n391), .C1(new_n293), .C2(new_n390), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT10), .ZN(new_n393));
  INV_X1    g0193(.A(G169), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n384), .B(new_n395), .C1(G179), .C2(new_n390), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n316), .A2(new_n274), .B1(new_n229), .B2(new_n277), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT15), .B(G87), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(new_n276), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n272), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT67), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n281), .A2(G77), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n401), .B(new_n402), .C1(G77), .C2(new_n287), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n250), .A2(G238), .A3(G1698), .ZN(new_n405));
  INV_X1    g0205(.A(G107), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n404), .B(new_n405), .C1(new_n406), .C2(new_n250), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n255), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n310), .A2(G244), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n260), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n394), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n403), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n412), .A2(KEYINPUT68), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n410), .A2(G179), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(KEYINPUT68), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n403), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n410), .A2(G200), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n293), .C2(new_n410), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n393), .A2(new_n396), .A3(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n379), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G41), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(KEYINPUT5), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n257), .A2(G45), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT79), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G41), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT79), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n257), .A4(G45), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n423), .A2(KEYINPUT5), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n426), .A2(new_n430), .A3(G274), .A4(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n255), .ZN(new_n433));
  NOR2_X1   g0233(.A1(G250), .A2(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n251), .A2(G257), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n305), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G294), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n303), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n261), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n426), .A2(new_n431), .A3(new_n430), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n443), .A2(G264), .A3(new_n261), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT87), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  AOI211_X1 g0245(.A(new_n434), .B(new_n436), .C1(new_n302), .C2(new_n304), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n255), .B1(new_n446), .B2(new_n440), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT87), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(G264), .A3(new_n261), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n433), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n433), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n447), .A2(new_n452), .A3(new_n449), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n451), .A2(G200), .B1(new_n453), .B2(G190), .ZN(new_n454));
  INV_X1    g0254(.A(new_n272), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n287), .B(new_n455), .C1(G1), .C2(new_n303), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n456), .A2(new_n406), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n285), .A2(new_n406), .ZN(new_n458));
  XOR2_X1   g0258(.A(new_n458), .B(KEYINPUT25), .Z(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n250), .A2(new_n460), .A3(new_n229), .A4(G87), .ZN(new_n461));
  AOI211_X1 g0261(.A(G20), .B(new_n214), .C1(new_n302), .C2(new_n304), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n303), .A2(new_n216), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n229), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n229), .A2(G107), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT23), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT24), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n463), .A2(KEYINPUT24), .A3(new_n465), .A4(new_n467), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n272), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n454), .A2(new_n457), .A3(new_n459), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n451), .A2(G179), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n453), .A2(G169), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n472), .A2(new_n457), .A3(new_n459), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n261), .A2(G250), .A3(new_n425), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n251), .A2(G244), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n302), .B2(new_n304), .ZN(new_n482));
  NOR2_X1   g0282(.A1(G238), .A2(G1698), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n464), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n480), .B1(new_n487), .B2(new_n255), .ZN(new_n488));
  INV_X1    g0288(.A(G179), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n425), .A2(new_n259), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n488), .A2(KEYINPUT81), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n464), .B1(new_n482), .B2(new_n484), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n491), .B(new_n479), .C1(new_n494), .C2(new_n261), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(G179), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n305), .A2(new_n229), .A3(G68), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  INV_X1    g0298(.A(G97), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n276), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n229), .B1(new_n249), .B2(new_n498), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT82), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NOR3_X1   g0303(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n497), .B(new_n500), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n272), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n398), .A2(new_n285), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n456), .A2(new_n398), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n495), .A2(new_n394), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n492), .A2(new_n496), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n488), .A2(G190), .A3(new_n491), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n495), .A2(G200), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n505), .A2(new_n272), .B1(new_n285), .B2(new_n398), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n456), .A2(new_n214), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n515), .B(KEYINPUT83), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n512), .A2(new_n513), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n473), .A2(new_n478), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(G1698), .B1(new_n302), .B2(new_n304), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT4), .B1(new_n520), .B2(G244), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G283), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n250), .A2(G250), .A3(G1698), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n255), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n443), .A2(G257), .A3(new_n261), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n452), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT80), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n528), .A2(new_n529), .A3(G200), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n528), .B2(G200), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n456), .A2(new_n499), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n339), .A2(G107), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n273), .A2(G77), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n406), .A2(KEYINPUT6), .A3(G97), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n499), .A2(new_n406), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n539), .B2(KEYINPUT6), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G20), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n534), .A2(new_n535), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n533), .B1(new_n542), .B2(new_n272), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n285), .A2(new_n499), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n544), .B(KEYINPUT78), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n526), .A2(G190), .A3(new_n527), .A4(new_n452), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n532), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n543), .A2(new_n546), .B1(new_n394), .B2(new_n528), .ZN(new_n551));
  INV_X1    g0351(.A(new_n528), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n489), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n443), .A2(G270), .A3(new_n261), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT84), .B1(new_n556), .B2(new_n433), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n443), .A2(G270), .A3(new_n261), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT84), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n255), .C2(new_n432), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n305), .A2(G257), .A3(new_n251), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT85), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n250), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G303), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n520), .A2(KEYINPUT85), .A3(G257), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n305), .A2(G264), .A3(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n564), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n255), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n523), .B(new_n229), .C1(G33), .C2(new_n499), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n572), .B(new_n272), .C1(new_n229), .C2(G116), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT20), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT86), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n574), .B2(new_n573), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT86), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n285), .A2(new_n216), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n216), .C2(new_n456), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n571), .A2(G169), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n557), .A2(new_n560), .B1(new_n569), .B2(new_n255), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(G179), .A3(new_n582), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n561), .A2(new_n570), .A3(G190), .ZN(new_n588));
  INV_X1    g0388(.A(G200), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n588), .B(new_n581), .C1(new_n589), .C2(new_n586), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n394), .B1(new_n561), .B2(new_n570), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(KEYINPUT21), .A3(new_n582), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n585), .A2(new_n587), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n519), .A2(new_n555), .A3(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n422), .A2(new_n594), .ZN(G372));
  NAND4_X1  g0395(.A1(new_n478), .A2(new_n587), .A3(new_n592), .A4(new_n585), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT88), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n495), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n489), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n600), .A2(new_n509), .A3(new_n510), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n601), .A2(new_n517), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n473), .A2(new_n550), .A3(new_n554), .A4(new_n602), .ZN(new_n603));
  NOR4_X1   g0403(.A1(new_n586), .A2(new_n584), .A3(new_n394), .A4(new_n581), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT21), .B1(new_n591), .B2(new_n582), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT88), .A3(new_n587), .A4(new_n478), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n598), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n551), .A2(new_n553), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(new_n518), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT26), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n609), .A2(new_n611), .A3(new_n602), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(new_n601), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n422), .A2(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n414), .A2(new_n294), .A3(new_n415), .A4(new_n413), .ZN(new_n616));
  INV_X1    g0416(.A(new_n291), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n373), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n315), .B1(new_n357), .B2(new_n358), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(new_n297), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n393), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n615), .A2(new_n396), .A3(new_n622), .ZN(G369));
  NAND2_X1  g0423(.A1(new_n606), .A2(new_n587), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n284), .A2(G20), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n257), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G343), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n581), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n593), .B2(new_n633), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G330), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n473), .A2(new_n478), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n477), .A2(new_n631), .ZN(new_n639));
  INV_X1    g0439(.A(new_n478), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n638), .A2(new_n639), .B1(new_n640), .B2(new_n631), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n631), .B1(new_n606), .B2(new_n587), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n638), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n640), .B2(new_n632), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(G399));
  INV_X1    g0449(.A(new_n207), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(G41), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G1), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n504), .A2(new_n216), .ZN(new_n654));
  OAI22_X1  g0454(.A1(new_n653), .A2(new_n654), .B1(new_n231), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT29), .B1(new_n614), .B2(new_n632), .ZN(new_n657));
  INV_X1    g0457(.A(new_n601), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n611), .B1(new_n609), .B2(new_n602), .ZN(new_n659));
  AOI211_X1 g0459(.A(new_n658), .B(new_n659), .C1(new_n611), .C2(new_n610), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n603), .A2(new_n596), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n631), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n657), .B1(KEYINPUT29), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n586), .A2(new_n552), .A3(G179), .A4(new_n599), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT30), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n445), .A2(new_n450), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OR3_X1    g0467(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n586), .A2(new_n451), .A3(new_n599), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n489), .A3(new_n528), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n665), .B1(new_n664), .B2(new_n667), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n631), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT31), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g0475(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n631), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT90), .B1(new_n594), .B2(new_n632), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n532), .A2(new_n549), .B1(new_n551), .B2(new_n553), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(new_n478), .A3(new_n473), .A4(new_n518), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT90), .ZN(new_n681));
  NOR4_X1   g0481(.A1(new_n680), .A2(new_n681), .A3(new_n593), .A4(new_n631), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n675), .B(new_n677), .C1(new_n678), .C2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n663), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n656), .B1(new_n685), .B2(G1), .ZN(G364));
  INV_X1    g0486(.A(G45), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n232), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n305), .A2(new_n650), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n688), .B(new_n689), .C1(new_n247), .C2(new_n687), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n250), .A2(G355), .A3(new_n207), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n690), .B(new_n691), .C1(G116), .C2(new_n207), .ZN(new_n692));
  NOR2_X1   g0492(.A1(G13), .A2(G33), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G20), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n228), .B1(G20), .B2(new_n394), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n229), .A2(G190), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(G179), .A3(new_n589), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n250), .B1(new_n701), .B2(G311), .ZN(new_n702));
  NOR2_X1   g0502(.A1(G179), .A2(G200), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n229), .B1(new_n703), .B2(G190), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n589), .A2(G179), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT92), .ZN(new_n707));
  INV_X1    g0507(.A(G283), .ZN(new_n708));
  OAI221_X1 g0508(.A(new_n702), .B1(new_n439), .B2(new_n704), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XOR2_X1   g0509(.A(KEYINPUT33), .B(G317), .Z(new_n710));
  NOR2_X1   g0510(.A1(new_n489), .A2(new_n589), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n699), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n229), .A2(new_n293), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n705), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT94), .ZN(new_n716));
  INV_X1    g0516(.A(G303), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n699), .A2(new_n703), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n713), .B(new_n718), .C1(G329), .C2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G322), .ZN(new_n726));
  INV_X1    g0526(.A(new_n714), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n727), .A2(new_n489), .A3(G200), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n725), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n714), .A2(new_n711), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n709), .B(new_n730), .C1(G326), .C2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n565), .B1(new_n732), .B2(G50), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n700), .A2(KEYINPUT91), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n700), .A2(KEYINPUT91), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n734), .B1(new_n214), .B2(new_n715), .C1(new_n737), .C2(new_n277), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n707), .A2(new_n406), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n720), .A2(G159), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(KEYINPUT32), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n712), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n740), .A2(KEYINPUT32), .B1(G68), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n704), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(KEYINPUT93), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(KEYINPUT93), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n742), .B(new_n744), .C1(new_n499), .C2(new_n748), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n738), .B(new_n749), .C1(G58), .C2(new_n728), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n733), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT96), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n698), .B1(new_n752), .B2(new_n696), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n653), .B1(G45), .B2(new_n625), .ZN(new_n754));
  INV_X1    g0554(.A(new_n695), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n753), .B(new_n754), .C1(new_n635), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n637), .A2(new_n754), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G330), .B2(new_n635), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(G396));
  NAND2_X1  g0560(.A1(new_n614), .A2(new_n632), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n403), .A2(new_n631), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n416), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n420), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n764), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n614), .A2(new_n766), .A3(new_n632), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n684), .ZN(new_n769));
  INV_X1    g0569(.A(new_n754), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(KEYINPUT99), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(KEYINPUT99), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(new_n684), .C2(new_n768), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n764), .A2(new_n693), .ZN(new_n775));
  INV_X1    g0575(.A(G132), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n723), .A2(new_n776), .B1(new_n716), .B2(new_n202), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT98), .B(G143), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n728), .A2(new_n778), .B1(new_n743), .B2(G150), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n732), .A2(G137), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(new_n737), .C2(new_n324), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT34), .Z(new_n782));
  INV_X1    g0582(.A(new_n305), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n707), .A2(new_n222), .ZN(new_n784));
  OR3_X1    g0584(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n777), .B(new_n785), .C1(G58), .C2(new_n745), .ZN(new_n786));
  INV_X1    g0586(.A(new_n748), .ZN(new_n787));
  INV_X1    g0587(.A(new_n716), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n787), .A2(G97), .B1(new_n788), .B2(G107), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n216), .B2(new_n737), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n729), .A2(new_n439), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n707), .A2(new_n214), .B1(new_n708), .B2(new_n712), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n565), .B1(new_n717), .B2(new_n731), .C1(new_n723), .C2(new_n793), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n696), .B1(new_n786), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n696), .A2(new_n693), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT97), .Z(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n277), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n775), .A2(new_n754), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n774), .A2(new_n801), .ZN(G384));
  NAND3_X1  g0602(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n631), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(KEYINPUT102), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT102), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n672), .A2(new_n805), .A3(KEYINPUT31), .A4(new_n631), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n676), .B1(new_n672), .B2(new_n631), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(new_n678), .C2(new_n682), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n422), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT103), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n629), .B1(new_n359), .B2(new_n342), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n368), .A2(KEYINPUT100), .A3(new_n372), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n620), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT100), .B1(new_n368), .B2(new_n372), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n360), .A2(new_n813), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n367), .A2(KEYINPUT37), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n370), .A2(new_n619), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT37), .B1(new_n821), .B2(new_n813), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT38), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n334), .A2(new_n455), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n356), .A2(KEYINPUT16), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n358), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n629), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n315), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n370), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT37), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n820), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n827), .A2(new_n629), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n378), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n824), .B1(new_n834), .B2(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n290), .A2(new_n631), .ZN(new_n836));
  INV_X1    g0636(.A(new_n270), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n290), .B1(new_n267), .B2(new_n268), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n294), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n836), .B1(new_n291), .B2(new_n294), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n810), .A2(new_n843), .A3(new_n766), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT40), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n835), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n473), .A2(new_n478), .A3(new_n518), .ZN(new_n847));
  INV_X1    g0647(.A(new_n593), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n847), .A2(new_n848), .A3(new_n679), .A4(new_n632), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n681), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n519), .A2(new_n555), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n851), .A2(KEYINPUT90), .A3(new_n848), .A4(new_n632), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n808), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n764), .B(new_n842), .C1(new_n853), .C2(new_n807), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n378), .A2(new_n833), .ZN(new_n855));
  INV_X1    g0655(.A(new_n832), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT38), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n858), .B(new_n832), .C1(new_n378), .C2(new_n833), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n854), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n846), .B1(new_n845), .B2(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n812), .B(new_n861), .Z(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(G330), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n622), .A2(new_n396), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n422), .B2(new_n663), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n863), .B(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n291), .A2(new_n631), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n859), .B2(new_n824), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n855), .A2(new_n856), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n858), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n855), .A2(KEYINPUT38), .A3(new_n856), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n867), .B(new_n869), .C1(new_n873), .C2(new_n868), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n620), .A2(new_n828), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n416), .A2(new_n631), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n842), .B1(new_n767), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n875), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n874), .A2(new_n879), .A3(KEYINPUT101), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT101), .B1(new_n874), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n866), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n257), .B2(new_n625), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n216), .B1(new_n540), .B2(KEYINPUT35), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n885), .B(new_n230), .C1(KEYINPUT35), .C2(new_n540), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT36), .ZN(new_n887));
  NOR4_X1   g0687(.A1(new_n321), .A2(new_n322), .A3(new_n231), .A4(new_n277), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n222), .A2(G50), .ZN(new_n889));
  OAI211_X1 g0689(.A(G1), .B(new_n284), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n884), .A2(new_n887), .A3(new_n890), .ZN(G367));
  NAND2_X1  g0691(.A1(new_n516), .A2(new_n514), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n631), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n602), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n601), .B2(new_n893), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT43), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n895), .B(KEYINPUT104), .Z(new_n897));
  INV_X1    g0697(.A(KEYINPUT43), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n632), .B1(new_n543), .B2(new_n546), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n555), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n902), .B(new_n903), .C1(new_n554), .C2(new_n632), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT106), .Z(new_n905));
  OR2_X1    g0705(.A1(new_n905), .A2(new_n478), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n631), .B1(new_n906), .B2(new_n554), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n904), .A2(new_n647), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n896), .B(new_n899), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n907), .A2(new_n909), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n899), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n905), .A2(new_n645), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n912), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n257), .B1(new_n625), .B2(G45), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n636), .A2(new_n643), .A3(new_n641), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n645), .A2(new_n646), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n904), .B2(new_n648), .ZN(new_n922));
  NOR2_X1   g0722(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT109), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n904), .A2(new_n648), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n645), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n685), .B(new_n920), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n685), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n651), .B(KEYINPUT41), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n917), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n895), .A2(new_n755), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n748), .A2(new_n222), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G137), .B2(new_n720), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n732), .A2(new_n778), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n937), .B(new_n938), .C1(new_n277), .C2(new_n706), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G150), .B2(new_n728), .ZN(new_n940));
  INV_X1    g0740(.A(new_n737), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(G50), .ZN(new_n942));
  INV_X1    g0742(.A(new_n715), .ZN(new_n943));
  AOI22_X1  g0743(.A1(G58), .A2(new_n943), .B1(new_n743), .B2(G159), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n940), .A2(new_n250), .A3(new_n942), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT46), .B1(new_n716), .B2(new_n216), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n216), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n941), .A2(G283), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n745), .A2(G107), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n948), .A2(new_n783), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(G311), .B2(new_n732), .ZN(new_n952));
  INV_X1    g0752(.A(new_n706), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G294), .A2(new_n743), .B1(new_n953), .B2(G97), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n952), .B(new_n954), .C1(new_n717), .C2(new_n729), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n720), .A2(G317), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n945), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT47), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n696), .ZN(new_n959));
  INV_X1    g0759(.A(new_n689), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n697), .B1(new_n207), .B2(new_n398), .C1(new_n960), .C2(new_n240), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT110), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n959), .A2(new_n754), .A3(new_n962), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n915), .A2(new_n934), .B1(new_n935), .B2(new_n963), .ZN(G387));
  NAND2_X1  g0764(.A1(new_n685), .A2(new_n920), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n919), .B1(new_n663), .B2(new_n684), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n651), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n748), .A2(new_n398), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n317), .A2(new_n712), .B1(new_n222), .B2(new_n700), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n499), .B2(new_n707), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n715), .A2(new_n277), .B1(new_n719), .B2(new_n381), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n971), .A2(new_n783), .A3(new_n972), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n202), .B2(new_n729), .C1(new_n324), .C2(new_n731), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n728), .A2(G317), .B1(G311), .B2(new_n743), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n726), .B2(new_n731), .C1(new_n737), .C2(new_n717), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT48), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n708), .B2(new_n704), .C1(new_n439), .C2(new_n715), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT49), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n720), .A2(G326), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n783), .B(new_n980), .C1(new_n216), .C2(new_n706), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n974), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n696), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n689), .B1(new_n237), .B2(new_n687), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n654), .A2(new_n207), .A3(new_n250), .ZN(new_n985));
  AOI211_X1 g0785(.A(G45), .B(new_n654), .C1(G68), .C2(G77), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n316), .A2(G50), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT50), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n207), .A2(G107), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n697), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n770), .B1(new_n641), .B2(new_n695), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n983), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n967), .B(new_n993), .C1(new_n916), .C2(new_n919), .ZN(G393));
  XNOR2_X1  g0794(.A(new_n929), .B(new_n645), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n965), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(new_n651), .A3(new_n931), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n770), .B1(new_n905), .B2(new_n695), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n783), .B1(new_n720), .B2(new_n778), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n728), .A2(G159), .B1(new_n732), .B2(G150), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(KEYINPUT51), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n748), .A2(new_n277), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n737), .A2(new_n316), .B1(new_n222), .B2(new_n715), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n707), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G87), .A2(new_n1006), .B1(new_n1001), .B2(KEYINPUT51), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1002), .B(new_n1008), .C1(G50), .C2(new_n743), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT52), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n728), .A2(G311), .B1(new_n732), .B2(G317), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n739), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n717), .B2(new_n712), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n565), .B1(new_n439), .B2(new_n700), .C1(new_n1012), .C2(new_n1010), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n719), .A2(new_n726), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n715), .A2(new_n708), .B1(new_n704), .B2(new_n216), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n696), .B1(new_n1009), .B2(new_n1018), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n697), .B1(new_n499), .B2(new_n207), .C1(new_n960), .C2(new_n244), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n999), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n998), .B(new_n1021), .C1(new_n916), .C2(new_n996), .ZN(G390));
  NAND4_X1  g0822(.A1(new_n379), .A2(G330), .A3(new_n421), .A4(new_n810), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT113), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n865), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT114), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n683), .A2(G330), .A3(new_n766), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n842), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n810), .A2(new_n843), .A3(G330), .A4(new_n766), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n767), .A2(new_n877), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1027), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n767), .A2(new_n877), .ZN(new_n1034));
  AOI211_X1 g0834(.A(KEYINPUT114), .B(new_n1034), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n810), .A2(G330), .A3(new_n766), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n842), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n876), .B1(new_n662), .B2(new_n766), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n842), .C2(new_n1028), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1026), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1028), .A2(new_n842), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT112), .B2(new_n1037), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n867), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n1039), .B2(new_n842), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(new_n835), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n824), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT39), .B1(new_n872), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n857), .A2(new_n859), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1049), .B1(KEYINPUT39), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1032), .A2(new_n843), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT111), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n1053), .A3(new_n1044), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT111), .B1(new_n878), .B2(new_n867), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1043), .B(new_n1047), .C1(new_n1051), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1053), .B1(new_n1052), .B2(new_n1044), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n878), .A2(KEYINPUT111), .A3(new_n867), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n869), .B1(new_n873), .B2(new_n868), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1046), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n854), .A2(KEYINPUT112), .A3(G330), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1041), .B(new_n1057), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1057), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1026), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1040), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1064), .A2(new_n651), .A3(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1057), .B(new_n917), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n770), .B1(new_n799), .B2(new_n317), .ZN(new_n1072));
  XOR2_X1   g0872(.A(KEYINPUT54), .B(G143), .Z(new_n1073));
  AOI22_X1  g0873(.A1(new_n941), .A2(new_n1073), .B1(G137), .B2(new_n743), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n324), .B2(new_n748), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT115), .Z(new_n1076));
  NOR2_X1   g0876(.A1(new_n715), .A2(new_n381), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT53), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n250), .B1(new_n706), .B2(new_n202), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n724), .B2(G125), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT116), .Z(new_n1082));
  OAI22_X1  g0882(.A1(new_n729), .A2(new_n776), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G128), .B2(new_n732), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1076), .A2(new_n1079), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n737), .A2(new_n499), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1086), .B(new_n1003), .C1(G87), .C2(new_n788), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n729), .A2(new_n216), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n712), .A2(new_n406), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n565), .B1(new_n731), .B2(new_n708), .ZN(new_n1090));
  NOR4_X1   g0890(.A1(new_n784), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1087), .B(new_n1091), .C1(new_n439), .C2(new_n723), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1085), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n696), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1072), .B(new_n1094), .C1(new_n1051), .C2(new_n694), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1070), .A2(new_n1071), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(G378));
  OAI211_X1 g0897(.A(new_n1057), .B(new_n1067), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1066), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n854), .B(KEYINPUT40), .C1(new_n859), .C2(new_n824), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n844), .B1(new_n871), .B2(new_n872), .ZN(new_n1101));
  OAI211_X1 g0901(.A(G330), .B(new_n1100), .C1(new_n1101), .C2(KEYINPUT40), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n393), .A2(new_n396), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n384), .A2(new_n828), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1103), .B(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1106), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1103), .B1(new_n384), .B2(new_n828), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1104), .B1(new_n393), .B2(new_n396), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1102), .A2(KEYINPUT119), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT119), .B1(new_n1102), .B2(new_n1113), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT120), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n861), .A2(new_n1117), .A3(G330), .A4(new_n1112), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n860), .A2(new_n845), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1119), .A2(G330), .A3(new_n1100), .A4(new_n1112), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1116), .A2(new_n1122), .A3(new_n882), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n881), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n874), .A2(KEYINPUT101), .A3(new_n879), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1102), .A2(new_n1113), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT119), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1102), .A2(KEYINPUT119), .A3(new_n1113), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1120), .B(new_n1117), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1126), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1099), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT57), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n652), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(KEYINPUT57), .B(new_n1099), .C1(new_n1123), .C2(new_n1133), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT121), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1098), .A2(new_n1066), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n882), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1131), .A2(new_n1132), .A3(new_n1126), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT121), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT57), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1136), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n917), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n770), .B1(new_n1113), .B2(new_n693), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n706), .A2(new_n220), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n731), .A2(new_n216), .B1(new_n715), .B2(new_n277), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n936), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n708), .B2(new_n723), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n305), .B(new_n1152), .C1(G107), .C2(new_n728), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n398), .A2(new_n700), .B1(new_n712), .B2(new_n499), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT117), .Z(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n423), .A3(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT58), .Z(new_n1157));
  AOI22_X1  g0957(.A1(G137), .A2(new_n701), .B1(new_n943), .B2(new_n1073), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n729), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n748), .A2(new_n381), .B1(new_n776), .B2(new_n712), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(G125), .C2(new_n732), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1163));
  AOI21_X1  g0963(.A(G33), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n720), .B2(G124), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n324), .C2(new_n706), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(new_n336), .B2(G33), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1166), .A2(new_n1167), .B1(G50), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n696), .B1(new_n1157), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1148), .B(new_n1170), .C1(G50), .C2(new_n798), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1147), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1145), .A2(new_n1173), .ZN(G375));
  OAI22_X1  g0974(.A1(new_n843), .A2(new_n694), .B1(G68), .B2(new_n798), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n716), .A2(new_n499), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1176), .B(new_n968), .C1(G77), .C2(new_n1006), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n565), .B1(new_n729), .B2(new_n708), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n737), .A2(new_n406), .B1(new_n216), .B2(new_n712), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(G303), .C2(new_n724), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1177), .B(new_n1180), .C1(new_n439), .C2(new_n731), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT122), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n748), .A2(new_n202), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n743), .A2(new_n1073), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n305), .B(new_n1184), .C1(new_n723), .C2(new_n1159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1149), .B(new_n1185), .C1(G159), .C2(new_n788), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n728), .A2(G137), .B1(new_n732), .B2(G132), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n381), .C2(new_n700), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1182), .B1(new_n1183), .B2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n770), .B(new_n1175), .C1(new_n696), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1067), .B2(new_n917), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1036), .A2(new_n1026), .A3(new_n1040), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n933), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1191), .B1(new_n1193), .B2(new_n1041), .ZN(G381));
  OR2_X1    g0994(.A1(G387), .A2(G390), .ZN(new_n1195));
  OR3_X1    g0995(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1195), .A2(G384), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT123), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(G375), .A2(G378), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT124), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1201), .A2(KEYINPUT124), .A3(new_n1202), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1205), .A2(new_n1206), .ZN(G407));
  NAND2_X1  g1007(.A1(new_n1200), .A2(new_n630), .ZN(new_n1208));
  OAI211_X1 g1008(.A(G213), .B(new_n1208), .C1(new_n1205), .C2(new_n1206), .ZN(G409));
  NAND2_X1  g1009(.A1(new_n1142), .A2(new_n933), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1096), .A2(new_n1210), .A3(new_n1147), .A4(new_n1171), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n630), .A2(G213), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT60), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1192), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1192), .A2(new_n1214), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n651), .A4(new_n1068), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1217), .A2(G384), .A3(new_n1191), .ZN(new_n1218));
  AOI21_X1  g1018(.A(G384), .B1(new_n1217), .B2(new_n1191), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AND4_X1   g1020(.A1(new_n1143), .A2(new_n1146), .A3(KEYINPUT57), .A4(new_n1099), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1143), .B1(new_n1142), .B2(KEYINPUT57), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1172), .B1(new_n1223), .B2(new_n1136), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1213), .B(new_n1220), .C1(new_n1224), .C2(new_n1096), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT125), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT63), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(G393), .B(new_n759), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G387), .A2(G390), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1195), .A2(KEYINPUT126), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT126), .B1(new_n1195), .B2(new_n1230), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1229), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1232), .A2(new_n1229), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n630), .A2(G213), .A3(G2897), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1217), .A2(new_n1191), .ZN(new_n1239));
  INV_X1    g1039(.A(G384), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1217), .A2(G384), .A3(new_n1191), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n1236), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1238), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1096), .B1(new_n1145), .B2(new_n1173), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT63), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1225), .A2(KEYINPUT125), .A3(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1227), .A2(new_n1235), .A3(new_n1249), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1225), .A2(KEYINPUT62), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1245), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT62), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(new_n1255), .A3(new_n1213), .A4(new_n1220), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1247), .A2(KEYINPUT127), .A3(new_n1248), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT127), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1252), .B1(new_n1260), .B2(new_n1235), .ZN(G405));
  NAND2_X1  g1061(.A1(new_n1224), .A2(new_n1096), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1254), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(new_n1220), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1220), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1235), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1264), .A2(new_n1233), .A3(new_n1234), .A4(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(G402));
endmodule


