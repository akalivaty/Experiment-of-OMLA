//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT64), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT66), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n462), .B2(new_n464), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n472), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n461), .B1(new_n462), .B2(new_n464), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT67), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n461), .A2(G114), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n492), .A2(new_n487), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n486), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n472), .A2(new_n496), .A3(G138), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n461), .C1(new_n466), .C2(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT68), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n465), .A2(new_n468), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n495), .B1(new_n500), .B2(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT69), .Z(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(new_n507), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n511), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(new_n509), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(G89), .B1(new_n505), .B2(new_n506), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n513), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT70), .ZN(new_n530));
  INV_X1    g105(.A(G77), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI221_X1 g107(.A(KEYINPUT70), .B1(new_n531), .B2(new_n508), .C1(new_n513), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n530), .A2(G651), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT72), .B(G90), .Z(new_n537));
  AOI22_X1  g112(.A1(new_n514), .A2(new_n537), .B1(new_n509), .B2(G52), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n534), .A2(new_n535), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND2_X1  g117(.A1(new_n514), .A2(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(new_n522), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n516), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT74), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n513), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n514), .B2(G91), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n509), .B2(G53), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n509), .A2(new_n560), .A3(G53), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n565), .A2(new_n561), .A3(new_n562), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  OAI21_X1  g145(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT75), .Z(new_n572));
  AOI22_X1  g147(.A1(new_n514), .A2(G87), .B1(new_n509), .B2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n512), .A2(new_n576), .A3(G61), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n576), .B1(new_n512), .B2(G61), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n575), .B(G651), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n512), .A2(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT76), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n585), .A2(new_n577), .A3(new_n579), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n575), .B1(new_n586), .B2(G651), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n514), .A2(G86), .B1(new_n509), .B2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n514), .A2(G85), .B1(new_n509), .B2(G47), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n516), .B2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(new_n514), .A2(G92), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT10), .Z(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n513), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n509), .B2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G284));
  OAI21_X1  g178(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n567), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n567), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(new_n600), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT79), .B(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(G860), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n609), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n465), .A2(new_n468), .ZN(new_n616));
  NOR3_X1   g191(.A1(new_n616), .A2(new_n474), .A3(G2105), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT82), .B(G2100), .Z(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n472), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n480), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n461), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n623), .A2(new_n624), .A3(new_n630), .ZN(G156));
  XOR2_X1   g206(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n632));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2430), .Z(new_n635));
  AOI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n634), .B2(new_n635), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n637), .B(new_n641), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(G14), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n643), .ZN(G401));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  NOR2_X1   g224(.A1(G2072), .A2(G2078), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n442), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n649), .A2(new_n651), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n651), .B(KEYINPUT17), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n656), .B(new_n653), .C1(new_n649), .C2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n649), .A3(new_n652), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n664), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n665), .B2(new_n670), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n667), .A2(new_n669), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n675), .A2(new_n670), .A3(new_n664), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n673), .B(new_n676), .C1(new_n664), .C2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G6), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n588), .A2(new_n589), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT32), .B(G1981), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT86), .B(G16), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(G166), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(G22), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1971), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n687), .A2(new_n688), .ZN(new_n696));
  MUX2_X1   g271(.A(G23), .B(G288), .S(G16), .Z(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT33), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n689), .A2(new_n695), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(KEYINPUT88), .A3(KEYINPUT34), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n480), .A2(G119), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n472), .A2(G131), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n461), .A2(G107), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n707), .B(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G25), .B(new_n711), .S(G29), .Z(new_n712));
  XOR2_X1   g287(.A(KEYINPUT35), .B(G1991), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n690), .A2(G24), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT87), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G290), .B2(new_n691), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G1986), .Z(new_n719));
  NOR3_X1   g294(.A1(new_n706), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n721));
  AND3_X1   g296(.A1(new_n705), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n721), .B1(new_n705), .B2(new_n720), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  OAI22_X1  g300(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n705), .A2(new_n720), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n724), .A2(new_n725), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n705), .A2(new_n720), .A3(new_n721), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n608), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G4), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1348), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n549), .A2(new_n691), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G19), .B2(new_n691), .ZN(new_n738));
  INV_X1    g313(.A(G1341), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n684), .A2(G21), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G168), .B2(new_n684), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT31), .B(G11), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT94), .B(G28), .Z(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT30), .B2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n745), .B(new_n748), .C1(new_n629), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n738), .B2(new_n739), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n736), .A2(new_n740), .A3(new_n744), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n749), .A2(G35), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT96), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n749), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT29), .B(G2090), .Z(new_n756));
  XOR2_X1   g331(.A(new_n755), .B(new_n756), .Z(new_n757));
  XOR2_X1   g332(.A(KEYINPUT27), .B(G1996), .Z(new_n758));
  AOI22_X1  g333(.A1(new_n472), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n480), .A2(G129), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n763), .A2(KEYINPUT93), .A3(new_n749), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n749), .ZN(new_n765));
  OAI21_X1  g340(.A(KEYINPUT93), .B1(G29), .B2(G32), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n757), .B1(new_n758), .B2(new_n767), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n768), .B1(new_n758), .B2(new_n767), .C1(new_n734), .C2(new_n735), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n749), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n749), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2078), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n752), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n749), .A2(G33), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT25), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n465), .A2(new_n468), .A3(G127), .ZN(new_n778));
  NAND2_X1  g353(.A1(G115), .A2(G2104), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n461), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n777), .B(new_n780), .C1(G139), .C2(new_n472), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(new_n749), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2072), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT24), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n749), .B1(new_n784), .B2(G34), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n784), .B2(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G160), .B2(G29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n783), .B1(G2084), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n749), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT28), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n480), .A2(G128), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT91), .Z(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n793));
  INV_X1    g368(.A(G116), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G2105), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G140), .B2(new_n472), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n797), .A2(KEYINPUT92), .A3(G29), .ZN(new_n798));
  AOI21_X1  g373(.A(KEYINPUT92), .B1(new_n797), .B2(G29), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n790), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n684), .A2(G5), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G171), .B2(new_n684), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n801), .B1(G1961), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n788), .B(new_n804), .C1(G1961), .C2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n690), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT23), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n567), .B2(new_n684), .ZN(new_n809));
  INV_X1    g384(.A(G1956), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n787), .A2(G2084), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT95), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n812), .A2(KEYINPUT95), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n774), .A2(new_n805), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(KEYINPUT98), .B1(new_n732), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT98), .ZN(new_n818));
  INV_X1    g393(.A(new_n816), .ZN(new_n819));
  AOI211_X1 g394(.A(new_n818), .B(new_n819), .C1(new_n726), .C2(new_n731), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n817), .A2(new_n820), .ZN(G311));
  NAND2_X1  g396(.A1(new_n732), .A2(new_n816), .ZN(G150));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n513), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n516), .B1(new_n825), .B2(KEYINPUT99), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(KEYINPUT99), .B2(new_n825), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n514), .A2(G93), .B1(new_n509), .B2(G55), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n608), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n829), .B1(new_n548), .B2(new_n545), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n549), .A2(new_n827), .A3(new_n828), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n834), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT100), .Z(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n838), .B2(new_n839), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n832), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT102), .ZN(G145));
  OAI21_X1  g420(.A(KEYINPUT4), .B1(new_n498), .B2(KEYINPUT68), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n496), .B1(new_n472), .B2(G138), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n503), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n495), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n493), .B1(new_n492), .B2(new_n487), .ZN(new_n851));
  OR2_X1    g426(.A1(G102), .A2(G2105), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n852), .A2(new_n490), .A3(KEYINPUT67), .A4(G2104), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(KEYINPUT103), .A3(new_n486), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n848), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n763), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n781), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n797), .B(KEYINPUT104), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n480), .A2(G130), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n461), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(G142), .B2(new_n472), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(new_n711), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n619), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT105), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n860), .A2(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n860), .A2(new_n867), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G160), .B(new_n629), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G162), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n868), .A2(new_n876), .ZN(new_n880));
  AOI21_X1  g455(.A(G37), .B1(new_n880), .B2(new_n870), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT40), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n877), .A2(new_n878), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT106), .B1(new_n874), .B2(new_n876), .ZN(new_n884));
  OAI211_X1 g459(.A(KEYINPUT40), .B(new_n881), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n882), .A2(new_n886), .ZN(G395));
  XNOR2_X1  g462(.A(G305), .B(G166), .ZN(new_n888));
  XOR2_X1   g463(.A(G288), .B(G290), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n890), .B(KEYINPUT108), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n608), .A2(new_n567), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n600), .A2(G299), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT41), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(KEYINPUT107), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(KEYINPUT107), .B2(new_n900), .ZN(new_n902));
  INV_X1    g477(.A(new_n837), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n612), .ZN(new_n904));
  MUX2_X1   g479(.A(new_n897), .B(new_n902), .S(new_n904), .Z(new_n905));
  XOR2_X1   g480(.A(new_n894), .B(new_n905), .Z(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(G868), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n829), .A2(new_n601), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(G295));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n910), .A3(new_n908), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n894), .B(new_n905), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(new_n601), .ZN(new_n913));
  INV_X1    g488(.A(new_n908), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT109), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n915), .ZN(G331));
  XNOR2_X1  g491(.A(G301), .B(G168), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n903), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(new_n897), .ZN(new_n920));
  XNOR2_X1  g495(.A(G301), .B(G286), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n837), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(KEYINPUT110), .A3(new_n837), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n919), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n923), .B1(new_n927), .B2(new_n902), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(new_n893), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  INV_X1    g507(.A(new_n893), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n928), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT43), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n925), .A2(new_n926), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n918), .A2(new_n922), .B1(new_n900), .B2(new_n898), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n937), .A2(new_n920), .B1(new_n938), .B2(KEYINPUT111), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n938), .A2(KEYINPUT111), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n893), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n934), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT44), .B1(new_n936), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n930), .B2(new_n934), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n934), .A2(new_n941), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n946), .B2(KEYINPUT43), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n944), .B1(new_n948), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n856), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(G160), .A2(G40), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n953), .A2(KEYINPUT112), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT112), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G2067), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n797), .B(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n763), .B(G1996), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n711), .B(new_n713), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT113), .B1(G290), .B2(G1986), .ZN(new_n965));
  NAND2_X1  g540(.A1(G290), .A2(G1986), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n957), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT117), .ZN(new_n969));
  OAI21_X1  g544(.A(G8), .B1(new_n511), .B2(new_n518), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n970), .B(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n954), .B1(new_n951), .B2(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(G2090), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  INV_X1    g551(.A(new_n495), .ZN(new_n977));
  AOI21_X1  g552(.A(G1384), .B1(new_n848), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR4_X1   g555(.A1(G164), .A2(KEYINPUT116), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n974), .B(new_n975), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n856), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n983));
  INV_X1    g558(.A(G40), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n471), .A2(new_n984), .A3(new_n477), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n952), .B1(G164), .B2(G1384), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1971), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n969), .B(new_n973), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n982), .B2(new_n989), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT117), .B1(new_n993), .B2(new_n972), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n985), .B1(new_n978), .B2(new_n979), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n856), .A2(new_n979), .A3(new_n950), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n856), .A2(KEYINPUT114), .A3(new_n979), .A4(new_n950), .ZN(new_n1000));
  AOI211_X1 g575(.A(G2090), .B(new_n996), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n989), .ZN(new_n1002));
  OAI211_X1 g577(.A(G8), .B(new_n972), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(G288), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n856), .A2(new_n985), .A3(new_n950), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n572), .A2(G1976), .A3(new_n573), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(G8), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(G8), .A3(new_n1007), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT52), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1012), .B(new_n589), .C1(new_n583), .C2(new_n587), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n586), .A2(G651), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n589), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G1981), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(KEYINPUT49), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1013), .A2(KEYINPUT115), .A3(new_n1016), .A4(KEYINPUT49), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT49), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1006), .A2(G8), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1011), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1003), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n996), .B1(new_n999), .B2(new_n1000), .ZN(new_n1029));
  INV_X1    g604(.A(G2084), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n954), .B1(KEYINPUT45), .B2(new_n978), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n953), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1029), .A2(new_n1030), .B1(new_n743), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n991), .B1(new_n1033), .B2(G168), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n999), .A2(new_n1000), .ZN(new_n1035));
  INV_X1    g610(.A(new_n996), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1030), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1032), .A2(new_n743), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G286), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1028), .B1(new_n1034), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(G168), .A3(new_n1038), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1042), .A2(new_n1028), .A3(G8), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n995), .B(new_n1027), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n987), .B2(G2078), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2078), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1031), .A2(new_n953), .A3(KEYINPUT53), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n1029), .B2(G1961), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT122), .B(new_n1049), .C1(new_n1029), .C2(G1961), .ZN(new_n1053));
  AOI211_X1 g628(.A(G171), .B(new_n1047), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1048), .A2(KEYINPUT53), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n954), .B2(KEYINPUT124), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1055), .A2(new_n953), .A3(new_n1057), .A4(new_n983), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1046), .A2(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n854), .A2(KEYINPUT103), .A3(new_n486), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT103), .B1(new_n854), .B2(new_n486), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1384), .B1(new_n1062), .B2(new_n848), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT114), .B1(new_n1063), .B2(new_n979), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1000), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1036), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT123), .B1(new_n1029), .B2(G1961), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1059), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT54), .B1(new_n1071), .B2(G301), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1054), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1044), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(G301), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1047), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(G301), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1077), .A2(KEYINPUT125), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT125), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1074), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1348), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n856), .A2(new_n985), .A3(new_n950), .A4(new_n958), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1084), .B(KEYINPUT118), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1088), .B(KEYINPUT119), .C1(new_n1029), .C2(G1348), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n608), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n974), .B1(new_n980), .B2(new_n981), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n810), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT56), .B(G2072), .Z(new_n1093));
  OR2_X1    g668(.A1(new_n987), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n567), .B(KEYINPUT57), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1090), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1092), .A2(new_n1096), .A3(new_n1094), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1101), .B(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n1006), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n987), .B2(G1996), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n549), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT59), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1098), .A2(new_n1110), .A3(new_n1100), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1066), .A2(new_n735), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT119), .B1(new_n1115), .B2(new_n1088), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1083), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT60), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n600), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n608), .B1(new_n1122), .B2(KEYINPUT121), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1120), .A2(new_n1123), .B1(KEYINPUT121), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1121), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1109), .B(new_n1114), .C1(new_n1124), .C2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1081), .B1(new_n1104), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1025), .A2(G8), .A3(G168), .A4(new_n1039), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n989), .B1(new_n1066), .B2(G2090), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n972), .B1(new_n1131), .B2(G8), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT63), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1025), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G288), .A2(G1976), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1135), .A2(new_n1136), .B1(new_n1012), .B2(new_n686), .ZN(new_n1137));
  OAI221_X1 g712(.A(new_n1133), .B1(new_n1003), .B2(new_n1134), .C1(new_n1023), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1039), .A2(G8), .A3(G168), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(KEYINPUT63), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1076), .A2(G301), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1043), .B1(new_n1144), .B2(KEYINPUT51), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1142), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1042), .A2(G8), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1033), .A2(G168), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT51), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1034), .A2(new_n1028), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT62), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1141), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1026), .B1(new_n994), .B2(new_n992), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1139), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n968), .B1(new_n1129), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G1996), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n957), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT46), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n957), .B1(new_n763), .B2(new_n960), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1160), .A2(KEYINPUT126), .A3(new_n1161), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT47), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1164), .A2(KEYINPUT47), .A3(new_n1165), .ZN(new_n1169));
  INV_X1    g744(.A(new_n957), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n711), .A2(new_n714), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n962), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n792), .A2(new_n958), .A3(new_n796), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1170), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1170), .A2(G1986), .A3(G290), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1175), .A2(KEYINPUT48), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1175), .A2(KEYINPUT48), .B1(new_n957), .B2(new_n964), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1168), .A2(new_n1169), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1157), .A2(KEYINPUT127), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n1182));
  INV_X1    g757(.A(new_n968), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1151), .B(new_n1154), .C1(new_n1054), .C2(new_n1072), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1077), .A2(KEYINPUT125), .A3(new_n1078), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1184), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1109), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1122), .A2(KEYINPUT121), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n600), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1122), .A2(KEYINPUT121), .A3(new_n608), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1190), .B1(new_n1194), .B2(new_n1126), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1189), .B1(new_n1195), .B2(new_n1103), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1076), .A2(G301), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1151), .B2(KEYINPUT62), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1145), .A2(new_n1143), .ZN(new_n1199));
  OAI22_X1  g774(.A1(new_n1198), .A2(new_n1199), .B1(KEYINPUT63), .B2(new_n1140), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1138), .B1(new_n1200), .B2(new_n1154), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1183), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1182), .B1(new_n1202), .B2(new_n1179), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1181), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g779(.A1(new_n879), .A2(new_n881), .ZN(new_n1206));
  INV_X1    g780(.A(G319), .ZN(new_n1207));
  NOR4_X1   g781(.A1(G229), .A2(new_n1207), .A3(G401), .A4(G227), .ZN(new_n1208));
  NAND3_X1  g782(.A1(new_n1206), .A2(new_n947), .A3(new_n1208), .ZN(G225));
  INV_X1    g783(.A(G225), .ZN(G308));
endmodule


