//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n550, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n575,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(new_n459), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n471), .A2(new_n459), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  OR2_X1    g054(.A1(G102), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G114), .C2(new_n459), .ZN(new_n481));
  OAI211_X1 g056(.A(G126), .B(G2105), .C1(new_n469), .C2(new_n470), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n459), .C1(new_n469), .C2(new_n470), .ZN(new_n485));
  AND2_X1   g060(.A1(KEYINPUT67), .A2(KEYINPUT4), .ZN(new_n486));
  NOR2_X1   g061(.A1(KEYINPUT67), .A2(KEYINPUT4), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n484), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT67), .B(KEYINPUT4), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n459), .A2(G138), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n461), .A2(new_n490), .A3(KEYINPUT68), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n485), .A2(KEYINPUT66), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n461), .A2(new_n495), .A3(new_n491), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT4), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n483), .B1(new_n493), .B2(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT69), .A2(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(KEYINPUT69), .A2(KEYINPUT6), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  AND3_X1   g088(.A1(KEYINPUT69), .A2(KEYINPUT6), .A3(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT6), .B1(KEYINPUT69), .B2(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n512), .A2(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n506), .A2(new_n520), .ZN(G166));
  AOI22_X1  g096(.A1(new_n509), .A2(new_n510), .B1(new_n501), .B2(new_n502), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n500), .B1(new_n509), .B2(new_n510), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n523), .A2(new_n525), .A3(new_n527), .A4(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n516), .A2(new_n517), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n524), .A2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n522), .A2(G90), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n532), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n524), .A2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n522), .A2(G81), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g124(.A(KEYINPUT70), .B(KEYINPUT8), .Z(new_n550));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  OAI21_X1  g128(.A(G65), .B1(new_n516), .B2(new_n517), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G651), .B1(new_n522), .B2(G91), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT71), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n511), .A2(KEYINPUT9), .A3(G543), .A4(new_n560), .ZN(new_n561));
  OAI211_X1 g136(.A(G543), .B(new_n560), .C1(new_n514), .C2(new_n515), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n557), .A2(new_n558), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n501), .B2(new_n502), .ZN(new_n567));
  INV_X1    g142(.A(new_n555), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n511), .A2(G91), .A3(new_n503), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n569), .A2(new_n564), .A3(new_n561), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT72), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  OR2_X1    g149(.A1(new_n506), .A2(new_n520), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT73), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g152(.A1(G166), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(G303));
  NAND2_X1  g154(.A1(new_n522), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n524), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G288));
  INV_X1    g159(.A(G48), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n512), .A2(new_n585), .B1(new_n518), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n503), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n505), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(KEYINPUT74), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n590), .B1(new_n532), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n594), .A2(KEYINPUT74), .A3(G651), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n588), .B1(new_n592), .B2(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n532), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT75), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n601), .B(new_n597), .C1(new_n532), .C2(new_n598), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(G651), .A3(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n522), .A2(G85), .B1(new_n524), .B2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NOR2_X1   g181(.A1(G301), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n522), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n518), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n511), .A2(G54), .A3(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n532), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G79), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(new_n500), .ZN(new_n617));
  OAI21_X1  g192(.A(G651), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n612), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n607), .B1(new_n623), .B2(new_n606), .ZN(G284));
  AOI21_X1  g199(.A(new_n607), .B1(new_n623), .B2(new_n606), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n573), .B2(G868), .ZN(G297));
  XNOR2_X1  g202(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n623), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n472), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n474), .A2(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n459), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  INV_X1    g218(.A(G2100), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n640), .A2(new_n645), .A3(new_n646), .ZN(G156));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT79), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT80), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n673), .A2(new_n667), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT81), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n668), .B(KEYINPUT17), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n675), .B1(new_n667), .B2(new_n676), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n672), .B(new_n677), .C1(new_n678), .C2(new_n669), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n684), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n689), .B(new_n691), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n686), .A2(new_n687), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(new_n697));
  XOR2_X1   g272(.A(G1981), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT83), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n697), .B(new_n701), .ZN(G229));
  NAND2_X1  g277(.A1(G160), .A2(G29), .ZN(new_n703));
  INV_X1    g278(.A(G34), .ZN(new_n704));
  AOI21_X1  g279(.A(G29), .B1(new_n704), .B2(KEYINPUT24), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(KEYINPUT24), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2084), .ZN(new_n708));
  INV_X1    g283(.A(G1961), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NOR2_X1   g285(.A1(G171), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G5), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G33), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n715));
  NAND3_X1  g290(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n472), .A2(G139), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(new_n459), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n719), .B1(KEYINPUT89), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(KEYINPUT89), .B2(new_n721), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n714), .B1(new_n723), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2072), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n708), .B1(new_n709), .B2(new_n712), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n713), .A2(G27), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G164), .B2(new_n713), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G2078), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n713), .A2(G32), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n474), .A2(G129), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT90), .Z(new_n737));
  INV_X1    g312(.A(G141), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n462), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n730), .B1(new_n741), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT93), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n729), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n726), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n744), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n728), .A2(G2078), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n724), .A2(new_n725), .ZN(new_n749));
  AND3_X1   g324(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G11), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n713), .B1(new_n753), .B2(G28), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(KEYINPUT95), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(G28), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n754), .B2(KEYINPUT95), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n752), .B1(new_n755), .B2(new_n757), .C1(new_n639), .C2(new_n713), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT96), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n713), .A2(G35), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n713), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT29), .B(G2090), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n712), .A2(new_n709), .ZN(new_n764));
  NOR2_X1   g339(.A1(G16), .A2(G19), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n547), .B2(G16), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G1341), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n759), .A2(new_n763), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n713), .A2(G26), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT86), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n472), .A2(G140), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n474), .A2(G128), .ZN(new_n773));
  OR2_X1    g348(.A1(G104), .A2(G2105), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n771), .B1(new_n777), .B2(new_n713), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT87), .B(G2067), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n710), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n710), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n780), .B(new_n784), .C1(G1341), .C2(new_n766), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n768), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n710), .A2(G20), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT23), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n573), .B2(new_n710), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1956), .Z(new_n790));
  NAND4_X1  g365(.A1(new_n746), .A2(new_n750), .A3(new_n786), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n710), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n623), .B2(new_n710), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1348), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n710), .A2(G23), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n583), .B2(new_n710), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n710), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n710), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n710), .A2(G6), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n594), .A2(G651), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n591), .A2(KEYINPUT74), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n587), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n807), .B1(new_n812), .B2(new_n710), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT84), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT32), .B(G1981), .Z(new_n815));
  AOI21_X1  g390(.A(new_n806), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n713), .A2(G25), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n472), .A2(G131), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n474), .A2(G119), .ZN(new_n822));
  OR2_X1    g397(.A1(G95), .A2(G2105), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n823), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n820), .B1(new_n826), .B2(new_n713), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G1991), .Z(new_n828));
  XOR2_X1   g403(.A(new_n827), .B(new_n828), .Z(new_n829));
  MUX2_X1   g404(.A(G24), .B(G290), .S(G16), .Z(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(G1986), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(G1986), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n818), .A2(new_n819), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT85), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT36), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(KEYINPUT36), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n818), .A2(new_n837), .A3(new_n819), .A4(new_n833), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n796), .B1(new_n836), .B2(new_n838), .ZN(G311));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n838), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(new_n795), .ZN(new_n842));
  AOI211_X1 g417(.A(KEYINPUT97), .B(new_n796), .C1(new_n836), .C2(new_n838), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(G150));
  NAND2_X1  g419(.A1(new_n623), .A2(G559), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  INV_X1    g424(.A(G67), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n532), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G651), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT99), .B(G93), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n522), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n524), .A2(G55), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n546), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n546), .A2(new_n856), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n848), .B(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(G860), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n861), .A2(KEYINPUT100), .A3(KEYINPUT39), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n864));
  INV_X1    g439(.A(new_n860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n848), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n862), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n856), .A2(G860), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT101), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(G145));
  NAND2_X1  g448(.A1(new_n493), .A2(new_n497), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT103), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT103), .B1(new_n481), .B2(new_n482), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n776), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n826), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n472), .A2(G142), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n474), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n459), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n642), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n879), .B(new_n825), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n723), .A2(new_n740), .ZN(new_n892));
  INV_X1    g467(.A(new_n741), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(new_n723), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n887), .A2(new_n890), .A3(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G160), .B(KEYINPUT102), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n478), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n639), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g481(.A(new_n631), .B(new_n865), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n617), .B1(new_n503), .B2(G66), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n613), .B1(new_n908), .B2(new_n505), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n611), .B2(new_n608), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n565), .A3(new_n572), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n910), .A2(new_n565), .A3(new_n572), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(KEYINPUT105), .A3(new_n914), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n919), .B1(new_n573), .B2(new_n619), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT107), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n917), .A2(new_n923), .A3(new_n918), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n573), .A2(new_n619), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n573), .A2(new_n927), .A3(new_n619), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n915), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n919), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n922), .A2(new_n924), .A3(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n907), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n912), .A2(KEYINPUT105), .A3(new_n914), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT105), .B1(new_n912), .B2(new_n914), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n907), .A2(new_n925), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n583), .A2(new_n603), .A3(new_n604), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n583), .B1(new_n603), .B2(new_n604), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT108), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(G290), .A2(G288), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(G305), .A2(new_n575), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n812), .A2(G166), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n940), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n947), .A2(new_n942), .A3(new_n941), .A4(new_n937), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT110), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n948), .A3(KEYINPUT109), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n950), .B2(KEYINPUT109), .ZN(new_n952));
  MUX2_X1   g527(.A(new_n950), .B(new_n952), .S(KEYINPUT42), .Z(new_n953));
  AND3_X1   g528(.A1(new_n932), .A2(new_n936), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n932), .B2(new_n936), .ZN(new_n955));
  OAI21_X1  g530(.A(G868), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n856), .A2(new_n606), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(G295));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n957), .ZN(G331));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  AND2_X1   g535(.A1(G301), .A2(G286), .ZN(new_n961));
  NOR2_X1   g536(.A1(G301), .A2(G286), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n858), .A2(new_n859), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G171), .A2(G168), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n542), .A2(G651), .B1(new_n522), .B2(G81), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n851), .A2(G651), .B1(G55), .B2(new_n524), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n965), .A2(new_n966), .A3(new_n544), .A4(new_n854), .ZN(new_n967));
  NAND2_X1  g542(.A1(G301), .A2(G286), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n964), .A2(new_n857), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n931), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n963), .A2(KEYINPUT111), .A3(new_n969), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n860), .A2(new_n974), .A3(new_n968), .A4(new_n964), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n925), .B2(new_n935), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n949), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n951), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n972), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n929), .A2(KEYINPUT41), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n917), .A2(new_n925), .A3(new_n918), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n976), .B(new_n984), .C1(new_n985), .C2(KEYINPUT41), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n970), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(G37), .B1(new_n988), .B2(new_n981), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n977), .B1(new_n931), .B2(new_n971), .ZN(new_n993));
  AOI21_X1  g568(.A(G37), .B1(new_n993), .B2(new_n982), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n921), .A2(KEYINPUT107), .B1(new_n919), .B2(new_n929), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n970), .B1(new_n995), .B2(new_n924), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n981), .B1(new_n996), .B2(new_n977), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n992), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n960), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n960), .B1(new_n990), .B2(KEYINPUT43), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n997), .A2(new_n983), .A3(new_n992), .A4(new_n904), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT112), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI211_X1 g577(.A(new_n977), .B(new_n981), .C1(new_n931), .C2(new_n971), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n935), .A2(new_n919), .A3(new_n925), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n973), .A2(new_n975), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(KEYINPUT41), .B2(new_n929), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1004), .A2(new_n1006), .B1(new_n985), .B2(new_n970), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n904), .B1(new_n1007), .B2(new_n982), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT43), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  AND4_X1   g584(.A1(KEYINPUT112), .A2(new_n1001), .A3(new_n1009), .A4(KEYINPUT44), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n999), .B1(new_n1002), .B2(new_n1010), .ZN(G397));
  INV_X1    g586(.A(G91), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n518), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n505), .B1(new_n554), .B2(new_n555), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT117), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n564), .A2(new_n561), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n569), .A2(new_n1017), .A3(new_n570), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1016), .A2(KEYINPUT57), .A3(new_n557), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT115), .B(G1956), .Z(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G40), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n464), .A2(new_n467), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G164), .A2(G1384), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT4), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n485), .B2(KEYINPUT66), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n489), .A2(new_n492), .B1(new_n1037), .B2(new_n496), .ZN(new_n1038));
  INV_X1    g613(.A(new_n876), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT103), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1035), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT50), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1028), .B1(new_n1034), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(G164), .B2(G1384), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT45), .B(new_n1035), .C1(new_n1038), .C2(new_n1041), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(new_n1030), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT56), .B(G2072), .Z(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1026), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT118), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1384), .B1(new_n874), .B2(new_n877), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1031), .B1(new_n1056), .B2(KEYINPUT45), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1049), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1046), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1035), .B1(new_n1038), .B2(new_n483), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1030), .B1(new_n1060), .B2(KEYINPUT50), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1056), .A2(new_n1033), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1027), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1055), .A2(new_n1059), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1051), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT61), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1030), .B(new_n1035), .C1(new_n1038), .C2(new_n1041), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(G2067), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1033), .B(new_n1035), .C1(new_n1038), .C2(new_n1041), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1030), .ZN(new_n1072));
  INV_X1    g647(.A(G1348), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT60), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n621), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n619), .B(KEYINPUT76), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(KEYINPUT60), .A3(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1074), .A2(KEYINPUT60), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1051), .A2(new_n1064), .A3(KEYINPUT61), .ZN(new_n1081));
  INV_X1    g656(.A(G1996), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1057), .A2(new_n1082), .A3(new_n1046), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1084), .B(G1341), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1068), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT59), .B1(new_n1087), .B2(new_n547), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n1089));
  AOI211_X1 g664(.A(new_n1089), .B(new_n546), .C1(new_n1083), .C2(new_n1086), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1067), .A2(new_n1080), .A3(new_n1081), .A4(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT119), .B1(new_n1074), .B2(new_n621), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1031), .B1(new_n1056), .B2(new_n1033), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1348), .B1(new_n1095), .B2(new_n1070), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1094), .B(new_n1077), .C1(new_n1096), .C2(new_n1069), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1051), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1064), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT120), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1101), .A3(new_n1064), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1092), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1030), .B1(new_n1056), .B2(KEYINPUT45), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(G2078), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1047), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1104), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1031), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1110), .A2(KEYINPUT123), .A3(new_n1047), .A4(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G2078), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1046), .A2(new_n1047), .A3(new_n1113), .A4(new_n1030), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1114), .A2(new_n1106), .B1(new_n1072), .B2(new_n709), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G171), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1045), .A2(G1384), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1038), .B2(new_n483), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1110), .A2(new_n1119), .A3(new_n1107), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1115), .A2(G301), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(KEYINPUT54), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT124), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1117), .A2(new_n1124), .A3(KEYINPUT54), .A4(new_n1121), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n1127));
  INV_X1    g702(.A(G2084), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1070), .A2(new_n1071), .A3(new_n1128), .A4(new_n1030), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1095), .A2(KEYINPUT113), .A3(new_n1128), .A4(new_n1070), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1030), .B(new_n1119), .C1(new_n1056), .C2(KEYINPUT45), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n783), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G8), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1127), .B1(new_n1136), .B2(KEYINPUT122), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(G286), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1131), .A2(new_n1132), .A3(G168), .A4(new_n1134), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(G8), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1135), .B2(G8), .ZN(new_n1143));
  OAI211_X1 g718(.A(G8), .B(new_n1139), .C1(new_n1143), .C2(new_n1127), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n576), .A2(G8), .A3(new_n578), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT55), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n576), .A2(KEYINPUT55), .A3(G8), .A4(new_n578), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1072), .A2(G2090), .ZN(new_n1151));
  AOI21_X1  g726(.A(G1971), .B1(new_n1057), .B2(new_n1046), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1150), .B(G8), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(G1981), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1154), .B(new_n588), .C1(new_n592), .C2(new_n595), .ZN(new_n1155));
  OAI21_X1  g730(.A(G1981), .B1(new_n587), .B2(new_n591), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT49), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1155), .A2(KEYINPUT49), .A3(new_n1156), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1159), .A2(G8), .A3(new_n1068), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(G1976), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT52), .B1(G288), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n583), .A2(G1976), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1068), .A2(new_n1163), .A3(G8), .A4(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1068), .A2(G8), .A3(new_n1164), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT52), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1161), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1048), .A2(new_n803), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1034), .A2(new_n1043), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1169), .B1(new_n1170), .B2(G2090), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1171), .A2(G8), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1153), .B(new_n1168), .C1(new_n1172), .C2(new_n1150), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(G171), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(G171), .B2(new_n1116), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1103), .A2(new_n1126), .A3(new_n1145), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1168), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1068), .A2(G8), .ZN(new_n1181));
  NOR2_X1   g756(.A1(G288), .A2(G1976), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1161), .A2(new_n1182), .B1(new_n1154), .B2(new_n812), .ZN(new_n1183));
  OAI22_X1  g758(.A1(new_n1180), .A2(new_n1153), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1135), .A2(G8), .A3(G168), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT114), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT114), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1135), .A2(new_n1187), .A3(G8), .A4(G168), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1168), .A2(new_n1153), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1150), .B1(new_n1171), .B2(G8), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1169), .B1(G2090), .B2(new_n1072), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1196), .A2(G8), .ZN(new_n1197));
  OAI21_X1  g772(.A(KEYINPUT63), .B1(new_n1197), .B2(new_n1150), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n1190), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1189), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1184), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1141), .A2(new_n1202), .A3(new_n1144), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1202), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n1206));
  OAI211_X1 g781(.A(new_n1203), .B(new_n1204), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  AOI211_X1 g782(.A(KEYINPUT125), .B(new_n1202), .C1(new_n1141), .C2(new_n1144), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1179), .B(new_n1201), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1056), .A2(new_n1031), .A3(KEYINPUT45), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n893), .A2(new_n1082), .ZN(new_n1211));
  OR2_X1    g786(.A1(new_n776), .A2(G2067), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n776), .A2(G2067), .ZN(new_n1213));
  AND2_X1   g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n740), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1215), .A2(G1996), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1211), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  OR2_X1    g792(.A1(new_n826), .A2(new_n828), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n826), .A2(new_n828), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(G290), .B(G1986), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1210), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1209), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g798(.A(new_n1214), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1210), .B1(new_n1224), .B2(new_n1215), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1210), .A2(new_n1082), .ZN(new_n1226));
  AND2_X1   g801(.A1(new_n1226), .A2(KEYINPUT46), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1226), .A2(KEYINPUT46), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1225), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  XOR2_X1   g804(.A(new_n1229), .B(KEYINPUT47), .Z(new_n1230));
  NOR2_X1   g805(.A1(G290), .A2(G1986), .ZN(new_n1231));
  AOI21_X1  g806(.A(KEYINPUT48), .B1(new_n1210), .B2(new_n1231), .ZN(new_n1232));
  AND3_X1   g807(.A1(new_n1210), .A2(KEYINPUT48), .A3(new_n1231), .ZN(new_n1233));
  AOI211_X1 g808(.A(new_n1232), .B(new_n1233), .C1(new_n1220), .C2(new_n1210), .ZN(new_n1234));
  INV_X1    g809(.A(new_n1217), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1212), .B1(new_n1235), .B2(new_n1219), .ZN(new_n1236));
  AOI211_X1 g811(.A(new_n1230), .B(new_n1234), .C1(new_n1210), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1223), .A2(new_n1237), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g813(.A1(new_n991), .A2(new_n998), .ZN(new_n1240));
  INV_X1    g814(.A(G319), .ZN(new_n1241));
  NOR2_X1   g815(.A1(G227), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g816(.A1(new_n665), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g817(.A1(new_n1243), .A2(KEYINPUT126), .ZN(new_n1244));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1245));
  NAND3_X1  g819(.A1(new_n665), .A2(new_n1245), .A3(new_n1242), .ZN(new_n1246));
  AOI21_X1  g820(.A(G229), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g821(.A1(new_n905), .A2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g822(.A1(new_n1240), .A2(new_n1248), .ZN(G308));
  OR2_X1    g823(.A1(new_n1240), .A2(new_n1248), .ZN(G225));
endmodule


