//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n212), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n203), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n209), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n222), .B1(new_n202), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(G87), .B2(G250), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  AND2_X1   g0027(.A1(KEYINPUT67), .A2(G77), .ZN(new_n228));
  NOR2_X1   g0028(.A1(KEYINPUT67), .A2(G77), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n225), .B(new_n226), .C1(new_n227), .C2(new_n230), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n206), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OR2_X1    g0034(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n236));
  AND3_X1   g0036(.A1(new_n221), .A2(new_n235), .A3(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  AOI21_X1  g0053(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G226), .ZN(new_n259));
  INV_X1    g0059(.A(new_n257), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G274), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n259), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT69), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n269), .B1(new_n230), .B2(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n214), .A2(new_n261), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n264), .A2(new_n265), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n266), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT71), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n216), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT71), .B1(G20), .B2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT70), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OR3_X1    g0088(.A1(new_n287), .A2(new_n201), .A3(KEYINPUT8), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n216), .A2(G33), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n278), .B1(new_n279), .B2(new_n285), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n211), .A2(new_n213), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G1), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(G13), .A3(G20), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n211), .A2(new_n213), .A3(new_n297), .A4(new_n293), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G50), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n296), .B2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n297), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n299), .A2(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n277), .A2(G200), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n266), .A2(new_n275), .A3(new_n276), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G190), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n306), .B(new_n308), .C1(new_n305), .C2(new_n304), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(new_n304), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n277), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G179), .B2(new_n277), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n290), .B1(new_n296), .B2(G20), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(new_n299), .B1(new_n302), .B2(new_n290), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G58), .A2(G68), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n216), .B1(new_n203), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n283), .ZN(new_n320));
  NOR3_X1   g0120(.A1(KEYINPUT71), .A2(G20), .A3(G33), .ZN(new_n321));
  OAI21_X1  g0121(.A(G159), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT80), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n284), .A2(KEYINPUT80), .A3(G159), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n319), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT79), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT7), .B1(new_n267), .B2(G20), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT7), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT3), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n329), .B(new_n216), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n327), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(G33), .ZN(new_n336));
  AOI21_X1  g0136(.A(G20), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n327), .A2(new_n329), .ZN(new_n338));
  OAI21_X1  g0138(.A(G68), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n326), .B(KEYINPUT16), .C1(new_n334), .C2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT82), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n342));
  INV_X1    g0142(.A(new_n319), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT80), .B1(new_n284), .B2(G159), .ZN(new_n344));
  INV_X1    g0144(.A(G159), .ZN(new_n345));
  AOI211_X1 g0145(.A(new_n323), .B(new_n345), .C1(new_n282), .C2(new_n283), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n343), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n328), .A2(G68), .A3(new_n333), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n341), .B(new_n342), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n340), .A2(new_n349), .A3(new_n294), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n328), .A2(new_n333), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n343), .B1(new_n344), .B2(new_n346), .C1(new_n351), .C2(new_n202), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n341), .B1(new_n352), .B2(new_n342), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n317), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n267), .A2(G223), .A3(new_n268), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G87), .ZN(new_n356));
  INV_X1    g0156(.A(G226), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n355), .B(new_n356), .C1(new_n270), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n274), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n263), .A2(new_n260), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(G232), .B2(new_n258), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G179), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n312), .B2(new_n362), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n354), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT18), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n354), .A2(new_n367), .A3(new_n364), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n342), .B1(new_n347), .B2(new_n348), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT82), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n370), .A2(new_n349), .A3(new_n340), .A4(new_n294), .ZN(new_n371));
  INV_X1    g0171(.A(G190), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n359), .A2(new_n372), .A3(new_n361), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n362), .B2(G200), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n317), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT17), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n371), .A2(KEYINPUT17), .A3(new_n317), .A4(new_n374), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n366), .A2(new_n368), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n267), .A2(G232), .A3(new_n268), .ZN(new_n380));
  AND2_X1   g0180(.A1(KEYINPUT72), .A2(G107), .ZN(new_n381));
  NOR2_X1   g0181(.A1(KEYINPUT72), .A2(G107), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI221_X1 g0183(.A(new_n380), .B1(new_n267), .B2(new_n383), .C1(new_n270), .C2(new_n223), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n274), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n360), .B1(G244), .B2(new_n258), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(G179), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n388), .B(KEYINPUT74), .ZN(new_n389));
  INV_X1    g0189(.A(new_n294), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n286), .B1(new_n284), .B2(KEYINPUT73), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(KEYINPUT73), .B2(new_n284), .ZN(new_n392));
  INV_X1    g0192(.A(new_n230), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n281), .A2(G20), .ZN(new_n396));
  AOI22_X1  g0196(.A1(G20), .A2(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n390), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n296), .A2(G20), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G77), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n298), .A2(new_n400), .B1(new_n393), .B2(new_n297), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n312), .B2(new_n387), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n389), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n387), .A2(G200), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(new_n402), .C1(new_n372), .C2(new_n387), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT77), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT12), .B1(new_n297), .B2(G68), .ZN(new_n409));
  INV_X1    g0209(.A(G13), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(G1), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT12), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(G20), .A4(new_n202), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n399), .A2(G68), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n298), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT76), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n414), .B(KEYINPUT76), .C1(new_n298), .C2(new_n415), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n300), .B1(new_n282), .B2(new_n283), .ZN(new_n421));
  INV_X1    g0221(.A(G77), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n291), .A2(new_n422), .B1(new_n216), .B2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n294), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT11), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(KEYINPUT11), .B(new_n294), .C1(new_n421), .C2(new_n423), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n408), .B1(new_n419), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n426), .A2(new_n427), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n430), .A2(KEYINPUT77), .A3(new_n418), .A4(new_n420), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n335), .A2(new_n336), .A3(G232), .A4(G1698), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n335), .A2(new_n336), .A3(G226), .A4(new_n268), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT75), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT75), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n433), .A2(new_n434), .A3(new_n438), .A4(new_n435), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n274), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT13), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n360), .B1(G238), .B2(new_n258), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n444));
  OAI21_X1  g0244(.A(G200), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n442), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT13), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(G190), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n432), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT78), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n432), .A2(new_n445), .A3(new_n449), .A4(KEYINPUT78), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n432), .ZN(new_n455));
  OAI21_X1  g0255(.A(G169), .B1(new_n443), .B2(new_n444), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n447), .A2(new_n448), .ZN(new_n457));
  INV_X1    g0257(.A(G179), .ZN(new_n458));
  OAI22_X1  g0258(.A1(new_n456), .A2(KEYINPUT14), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT14), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n457), .B2(G169), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n455), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  NOR4_X1   g0263(.A1(new_n315), .A2(new_n379), .A3(new_n407), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT84), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT83), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n422), .B1(new_n282), .B2(new_n283), .ZN(new_n467));
  XNOR2_X1  g0267(.A(G97), .B(G107), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT6), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n469), .A2(new_n471), .A3(G107), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n467), .B1(new_n474), .B2(G20), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT72), .B(G107), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n328), .A2(new_n333), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n390), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n297), .A2(G97), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n281), .A2(G1), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n298), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n481), .B2(G97), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n466), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n477), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n472), .B1(new_n469), .B2(new_n468), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n486), .A2(new_n216), .B1(new_n422), .B2(new_n285), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n294), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(KEYINPUT83), .A3(new_n482), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT5), .B(G41), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n256), .A2(G1), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G257), .A3(new_n262), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n491), .A2(G274), .A3(new_n262), .A4(new_n492), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n335), .A2(new_n336), .A3(G244), .A4(new_n268), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .A4(new_n268), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n267), .A2(G250), .A3(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n496), .B1(new_n274), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G190), .ZN(new_n505));
  INV_X1    g0305(.A(G200), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(new_n504), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n465), .B1(new_n490), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n274), .ZN(new_n509));
  INV_X1    g0309(.A(new_n496), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(G190), .B2(new_n504), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(KEYINPUT84), .A3(new_n484), .A4(new_n489), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G169), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n504), .A2(G179), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n515), .A2(new_n516), .B1(new_n488), .B2(new_n482), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n267), .A2(new_n216), .A3(G87), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT22), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT22), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n267), .A2(new_n521), .A3(new_n216), .A4(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT23), .B1(new_n476), .B2(new_n216), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT91), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT23), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n216), .A2(G107), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n526), .A2(new_n527), .B1(new_n396), .B2(G116), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n524), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n525), .B1(new_n524), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(KEYINPUT24), .B(new_n523), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n294), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n411), .A2(new_n527), .ZN(new_n536));
  XOR2_X1   g0336(.A(new_n536), .B(KEYINPUT25), .Z(new_n537));
  INV_X1    g0337(.A(new_n481), .ZN(new_n538));
  INV_X1    g0338(.A(G107), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT92), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n537), .B(KEYINPUT92), .C1(new_n539), .C2(new_n538), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n254), .B1(new_n492), .B2(new_n491), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G264), .ZN(new_n546));
  MUX2_X1   g0346(.A(G250), .B(G257), .S(G1698), .Z(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n267), .B1(G33), .B2(G294), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n495), .C1(new_n548), .C2(new_n273), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G190), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(G200), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n535), .A2(new_n544), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  AND4_X1   g0353(.A1(new_n508), .A2(new_n513), .A3(new_n518), .A4(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G87), .A2(G97), .ZN(new_n555));
  NAND3_X1  g0355(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n383), .A2(new_n555), .B1(new_n216), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n335), .A2(new_n336), .A3(new_n216), .A4(G68), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT19), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n291), .B2(new_n471), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n294), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n481), .A2(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n394), .A2(new_n302), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT86), .ZN(new_n566));
  INV_X1    g0366(.A(G250), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n296), .B2(G45), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n262), .A3(KEYINPUT85), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n262), .A2(G274), .A3(new_n492), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT85), .B1(new_n568), .B2(new_n262), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n262), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT85), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n570), .A4(new_n569), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n267), .A2(G238), .A3(new_n268), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G33), .A2(G116), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n270), .C2(new_n227), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n573), .A2(new_n577), .B1(new_n580), .B2(new_n274), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n565), .B1(new_n581), .B2(new_n506), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT87), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n565), .B(KEYINPUT87), .C1(new_n581), .C2(new_n506), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n573), .A2(new_n577), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(new_n274), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(G190), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n458), .A3(new_n587), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n562), .B(new_n564), .C1(new_n538), .C2(new_n394), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(G169), .C2(new_n581), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT21), .ZN(new_n596));
  AOI21_X1  g0396(.A(G20), .B1(G33), .B2(G283), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n281), .A2(G97), .ZN(new_n598));
  INV_X1    g0398(.A(G116), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n597), .A2(new_n598), .B1(G20), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n294), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n294), .A3(KEYINPUT20), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(KEYINPUT90), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n297), .A2(new_n599), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n481), .B2(new_n599), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT90), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n601), .A2(new_n608), .A3(new_n602), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n605), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n335), .A2(new_n336), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n268), .ZN(new_n613));
  XNOR2_X1  g0413(.A(KEYINPUT89), .B(G303), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(G264), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n335), .A2(new_n336), .A3(G257), .A4(new_n268), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT88), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n267), .A2(KEYINPUT88), .A3(G257), .A4(new_n268), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n273), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n545), .A2(G270), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n495), .ZN(new_n623));
  OAI21_X1  g0423(.A(G169), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n596), .B1(new_n611), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n623), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n615), .A2(new_n620), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n273), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(KEYINPUT21), .A3(G169), .A4(new_n610), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n621), .A2(new_n458), .A3(new_n623), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n610), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n625), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n549), .A2(new_n312), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(G179), .B2(new_n549), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n535), .B2(new_n544), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n621), .A2(new_n623), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G190), .ZN(new_n637));
  OAI21_X1  g0437(.A(G200), .B1(new_n621), .B2(new_n623), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n637), .A2(new_n611), .A3(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n632), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n464), .A2(new_n554), .A3(new_n595), .A4(new_n640), .ZN(G372));
  AND2_X1   g0441(.A1(new_n366), .A2(new_n368), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n450), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n462), .B1(new_n644), .B2(new_n404), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n377), .A2(new_n378), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n310), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n314), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n464), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT93), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n588), .B(new_n565), .C1(new_n506), .C2(new_n581), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n593), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n593), .A2(new_n653), .A3(new_n652), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n484), .A2(new_n489), .B1(new_n515), .B2(new_n516), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n517), .B(new_n593), .C1(new_n584), .C2(new_n589), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT26), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n660), .A2(new_n593), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n632), .ZN(new_n664));
  INV_X1    g0464(.A(new_n635), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n554), .A2(new_n666), .A3(new_n657), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT94), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n593), .A2(new_n653), .A3(new_n652), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n669), .A2(new_n654), .B1(new_n632), .B2(new_n635), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n508), .A2(new_n513), .A3(new_n518), .A4(new_n553), .ZN(new_n671));
  OR3_X1    g0471(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT94), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n663), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n650), .B1(new_n651), .B2(new_n673), .ZN(G369));
  NAND2_X1  g0474(.A1(new_n411), .A2(new_n216), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n610), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n632), .B(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G330), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n682), .A2(new_n683), .A3(new_n639), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n535), .A2(new_n544), .ZN(new_n685));
  INV_X1    g0485(.A(new_n680), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n553), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n665), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n635), .A2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n664), .A2(new_n680), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n688), .A2(new_n693), .B1(new_n635), .B2(new_n686), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n207), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G1), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n383), .A2(new_n599), .A3(new_n555), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(new_n218), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  NAND4_X1  g0502(.A1(new_n554), .A2(new_n595), .A3(new_n640), .A4(new_n686), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n548), .A2(new_n273), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(G264), .B2(new_n545), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n581), .A2(new_n706), .A3(new_n504), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n626), .B(G179), .C1(new_n627), .C2(new_n273), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT95), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n707), .A2(new_n708), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT30), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT95), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n713), .B(new_n704), .C1(new_n707), .C2(new_n708), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n636), .A2(new_n581), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(new_n458), .A3(new_n514), .A4(new_n549), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n710), .A2(new_n712), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n680), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n712), .A2(new_n709), .A3(new_n716), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n703), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT98), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n593), .B1(new_n670), .B2(new_n671), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT96), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n661), .A2(new_n728), .A3(new_n658), .ZN(new_n729));
  OAI211_X1 g0529(.A(KEYINPUT26), .B(new_n659), .C1(new_n669), .C2(new_n654), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n728), .B1(new_n661), .B2(new_n658), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n727), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT97), .B1(new_n734), .B2(new_n680), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n729), .A2(new_n730), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n667), .B(new_n593), .C1(new_n736), .C2(new_n732), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT97), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n738), .A3(new_n686), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n726), .B1(new_n740), .B2(KEYINPUT29), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  AOI211_X1 g0542(.A(KEYINPUT98), .B(new_n742), .C1(new_n735), .C2(new_n739), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n668), .A2(new_n672), .ZN(new_n745));
  INV_X1    g0545(.A(new_n663), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n680), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n742), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n725), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n702), .B1(new_n751), .B2(new_n296), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT99), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n682), .A2(new_n639), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G330), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n410), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n296), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n697), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n684), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT100), .Z(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n682), .B2(new_n639), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n215), .B1(G20), .B2(new_n312), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT101), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n696), .A2(new_n612), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G355), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G116), .B2(new_n207), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n249), .A2(new_n256), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n267), .B(new_n696), .C1(new_n219), .C2(new_n256), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n760), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n458), .A2(G200), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(G20), .A3(new_n372), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n779), .A2(G20), .A3(G190), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n230), .A2(new_n780), .B1(new_n781), .B2(new_n201), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n216), .A2(new_n458), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n372), .A2(new_n506), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n216), .A2(G179), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n372), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G50), .A2(new_n786), .B1(new_n789), .B2(G107), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n783), .A2(new_n372), .A3(G200), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n790), .B(new_n267), .C1(new_n202), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n784), .A2(new_n787), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n782), .B(new_n792), .C1(G87), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G179), .A2(G200), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT102), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n797), .A2(new_n216), .A3(G190), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G159), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT32), .Z(new_n800));
  OAI21_X1  g0600(.A(G20), .B1(new_n797), .B2(new_n372), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G97), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n795), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT103), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n791), .B1(new_n805), .B2(KEYINPUT103), .ZN(new_n807));
  INV_X1    g0607(.A(new_n781), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n806), .A2(new_n807), .B1(G322), .B2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT104), .Z(new_n810));
  INV_X1    g0610(.A(G326), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n785), .A2(new_n811), .B1(new_n793), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G283), .B2(new_n789), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n798), .A2(G329), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n801), .A2(G294), .ZN(new_n816));
  INV_X1    g0616(.A(new_n780), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n267), .B1(new_n817), .B2(G311), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n803), .B1(new_n810), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n778), .B1(new_n820), .B2(new_n768), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n756), .A2(new_n761), .B1(new_n767), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  INV_X1    g0623(.A(new_n404), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n402), .A2(new_n686), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n407), .B2(new_n825), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n748), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n673), .A2(new_n680), .A3(new_n828), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n760), .B1(new_n832), .B2(new_n724), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n724), .B2(new_n832), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n769), .A2(new_n763), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n760), .B1(new_n835), .B2(G77), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n808), .A2(G143), .B1(new_n817), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n837), .B1(new_n838), .B2(new_n785), .C1(new_n279), .C2(new_n791), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT105), .Z(new_n840));
  OR2_X1    g0640(.A1(new_n840), .A2(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(KEYINPUT34), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n612), .B1(new_n789), .B2(G68), .ZN(new_n843));
  INV_X1    g0643(.A(new_n798), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n843), .B1(new_n300), .B2(new_n793), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G58), .B2(new_n801), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n841), .A2(new_n842), .A3(new_n847), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n785), .A2(new_n812), .B1(new_n780), .B2(new_n599), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n267), .B(new_n849), .C1(G107), .C2(new_n794), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n798), .A2(G311), .ZN(new_n851));
  INV_X1    g0651(.A(G283), .ZN(new_n852));
  INV_X1    g0652(.A(G87), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n791), .A2(new_n852), .B1(new_n788), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G294), .B2(new_n808), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n850), .A2(new_n802), .A3(new_n851), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n836), .B1(new_n857), .B2(new_n768), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n827), .B2(new_n763), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n834), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  OR2_X1    g0661(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n862), .A2(G116), .A3(new_n217), .A4(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT36), .Z(new_n865));
  NAND3_X1  g0665(.A1(new_n219), .A2(new_n393), .A3(new_n318), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n300), .A2(G68), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n296), .B(G13), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n456), .A2(KEYINPUT14), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n457), .A2(new_n460), .A3(G169), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n870), .B(new_n871), .C1(new_n458), .C2(new_n457), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n455), .A3(new_n686), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT110), .ZN(new_n875));
  INV_X1    g0675(.A(new_n317), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n339), .B1(new_n351), .B2(KEYINPUT79), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n342), .B1(new_n877), .B2(new_n347), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n294), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT108), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n326), .B1(new_n334), .B2(new_n339), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n879), .A2(new_n880), .B1(KEYINPUT16), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n878), .A2(KEYINPUT108), .A3(new_n294), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n876), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n678), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n379), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT109), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n379), .A2(KEYINPUT109), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n375), .B1(new_n885), .B2(new_n678), .ZN(new_n892));
  INV_X1    g0692(.A(new_n364), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n678), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n354), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n365), .A2(new_n897), .A3(new_n375), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n891), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n379), .A2(KEYINPUT109), .A3(new_n886), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT109), .B1(new_n379), .B2(new_n886), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n900), .B(KEYINPUT38), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT39), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n897), .B1(new_n642), .B2(new_n646), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n898), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n908), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n904), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n875), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n908), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n907), .B1(new_n916), .B2(new_n904), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n904), .A2(new_n907), .A3(new_n912), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT110), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n874), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n824), .A2(new_n686), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT106), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n747), .B2(new_n827), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n455), .A2(new_n680), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n459), .A2(new_n461), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n925), .B1(new_n454), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n450), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n872), .B2(new_n455), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT107), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n462), .A2(new_n450), .A3(new_n925), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT107), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n872), .B1(new_n452), .B2(new_n453), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n931), .B(new_n932), .C1(new_n933), .C2(new_n925), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n924), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n916), .A2(new_n904), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n936), .A2(new_n937), .B1(new_n643), .B2(new_n678), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n920), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n651), .B1(new_n748), .B2(new_n742), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n741), .B2(new_n743), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(new_n650), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n939), .B(new_n942), .Z(new_n943));
  NAND2_X1  g0743(.A1(new_n904), .A2(new_n912), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n703), .A2(new_n720), .A3(new_n945), .ZN(new_n946));
  AND4_X1   g0746(.A1(new_n827), .A2(new_n930), .A3(new_n946), .A4(new_n934), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT40), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n937), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n464), .A2(new_n946), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n683), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n943), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n296), .B2(new_n757), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n943), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n869), .B1(new_n957), .B2(new_n958), .ZN(G367));
  XOR2_X1   g0759(.A(new_n690), .B(new_n693), .Z(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n684), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n750), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n490), .A2(new_n680), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n508), .A2(new_n513), .A3(new_n518), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n659), .A2(new_n680), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n694), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT45), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n694), .A2(new_n966), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT44), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n971), .A2(new_n692), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n692), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT112), .B1(new_n962), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT112), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n750), .A2(new_n974), .A3(new_n977), .A4(new_n961), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n751), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n697), .B(KEYINPUT41), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n758), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n966), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n692), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT111), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n565), .A2(new_n686), .ZN(new_n985));
  MUX2_X1   g0785(.A(new_n657), .B(new_n594), .S(new_n985), .Z(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n984), .B(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n691), .A2(new_n693), .A3(new_n966), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT42), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n966), .A2(new_n635), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n680), .B1(new_n992), .B2(new_n518), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n989), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n988), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n981), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n696), .A2(new_n267), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n245), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n207), .B2(new_n394), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n760), .B1(new_n771), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT114), .B(G317), .Z(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT46), .B1(new_n794), .B2(G116), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n844), .A2(new_n1001), .B1(KEYINPUT113), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(KEYINPUT113), .B2(new_n1002), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n794), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n614), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n612), .C1(new_n1006), .C2(new_n781), .ZN(new_n1007));
  INV_X1    g0807(.A(G294), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n791), .A2(new_n1008), .B1(new_n780), .B2(new_n852), .ZN(new_n1009));
  INV_X1    g0809(.A(G311), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n1010), .A2(new_n785), .B1(new_n788), .B2(new_n471), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1007), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n801), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1004), .B(new_n1012), .C1(new_n383), .C2(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n844), .A2(new_n838), .B1(new_n201), .B2(new_n793), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT115), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G143), .A2(new_n786), .B1(new_n808), .B2(G150), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G50), .A2(new_n817), .B1(new_n789), .B2(new_n393), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n791), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n612), .B(new_n1020), .C1(G159), .C2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1017), .B(new_n1022), .C1(new_n202), .C2(new_n1013), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1014), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT47), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1000), .B1(new_n1026), .B2(new_n768), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n765), .B2(new_n986), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n996), .A2(new_n1028), .ZN(G387));
  NAND2_X1  g0829(.A1(new_n242), .A2(G45), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1030), .A2(new_n997), .B1(new_n700), .B2(new_n772), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n286), .A2(G50), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT50), .Z(new_n1033));
  OAI21_X1  g0833(.A(new_n256), .B1(new_n202), .B2(new_n422), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1033), .A2(new_n700), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n539), .B2(new_n696), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n760), .B1(new_n1037), .B2(new_n771), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n691), .A2(new_n765), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n290), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G150), .A2(new_n798), .B1(new_n1040), .B2(new_n1021), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n801), .A2(new_n395), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n612), .B1(new_n789), .B2(G97), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n785), .A2(new_n345), .B1(new_n793), .B2(new_n230), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n781), .A2(new_n300), .B1(new_n780), .B2(new_n202), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n267), .B1(new_n789), .B2(G116), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1001), .A2(new_n781), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1006), .A2(new_n780), .B1(new_n791), .B2(new_n1010), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G322), .C2(new_n786), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1051), .A2(KEYINPUT48), .B1(G283), .B2(new_n801), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(KEYINPUT48), .B2(new_n1051), .C1(new_n1008), .C2(new_n793), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1048), .B1(new_n811), .B2(new_n844), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1047), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1038), .B(new_n1039), .C1(new_n768), .C2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n961), .B2(new_n759), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n962), .A2(KEYINPUT116), .A3(new_n697), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n750), .B2(new_n961), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT116), .B1(new_n962), .B2(new_n697), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(G393));
  NAND2_X1  g0863(.A1(new_n982), .A2(new_n766), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n252), .A2(new_n997), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n471), .B2(new_n207), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n760), .B1(new_n771), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n267), .B1(new_n788), .B2(new_n853), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n794), .A2(G68), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n300), .B2(new_n791), .C1(new_n286), .C2(new_n780), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(G143), .C2(new_n798), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n801), .A2(G77), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n785), .A2(new_n279), .B1(new_n781), .B2(new_n345), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G317), .A2(new_n786), .B1(new_n808), .B2(G311), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT52), .Z(new_n1078));
  OAI22_X1  g0878(.A1(new_n1006), .A2(new_n791), .B1(new_n780), .B2(new_n1008), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n267), .B(new_n1079), .C1(G107), .C2(new_n789), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n599), .C2(new_n1013), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n798), .A2(G322), .B1(G283), .B2(new_n794), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT118), .Z(new_n1083));
  OAI21_X1  g0883(.A(new_n1076), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1068), .B1(new_n1084), .B2(new_n768), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1065), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n975), .B2(new_n758), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n976), .A2(new_n978), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n698), .B1(new_n962), .B2(new_n975), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G390));
  INV_X1    g0891(.A(new_n739), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n738), .B1(new_n737), .B2(new_n686), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n827), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n725), .A2(new_n827), .A3(new_n930), .A4(new_n934), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n946), .A2(G330), .A3(new_n827), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n935), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n922), .A4(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n725), .A2(new_n827), .B1(new_n930), .B2(new_n934), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1096), .A2(new_n935), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1099), .A2(new_n1100), .B1(new_n830), .B2(new_n923), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n464), .A2(G330), .A3(new_n946), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1102), .A2(new_n941), .A3(new_n650), .A4(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n906), .A2(new_n875), .A3(new_n913), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT110), .B1(new_n917), .B2(new_n918), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n873), .B1(new_n924), .B2(new_n935), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n923), .B1(new_n740), .B2(new_n827), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n873), .B(new_n944), .C1(new_n1109), .C2(new_n935), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1108), .A2(new_n1110), .A3(new_n1095), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1100), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1104), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1100), .ZN(new_n1116));
  AND4_X1   g0916(.A1(new_n650), .A2(new_n1102), .A3(new_n941), .A4(new_n1103), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1108), .A2(new_n1110), .A3(new_n1095), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1114), .A2(new_n1119), .A3(new_n697), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n759), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1105), .A2(new_n1106), .A3(new_n762), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n760), .B1(new_n835), .B2(new_n1040), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n788), .A2(new_n202), .B1(new_n781), .B2(new_n599), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n267), .B(new_n1125), .C1(G87), .C2(new_n794), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n798), .A2(G294), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n791), .A2(new_n383), .B1(new_n780), .B2(new_n471), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G283), .B2(new_n786), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1126), .A2(new_n1073), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G128), .A2(new_n786), .B1(new_n808), .B2(G132), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT119), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n345), .B2(new_n1013), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n793), .A2(new_n279), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n798), .A2(G125), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT54), .B(G143), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n612), .B1(new_n817), .B2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G137), .A2(new_n1021), .B1(new_n789), .B2(G50), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1135), .A2(new_n1136), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1130), .B1(new_n1133), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1124), .B1(new_n1142), .B2(new_n768), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1123), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1120), .A2(new_n1122), .A3(new_n1144), .ZN(G378));
  AND2_X1   g0945(.A1(new_n942), .A2(new_n1103), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1119), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n311), .A2(new_n678), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n315), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n315), .A2(new_n1149), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OR3_X1    g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT40), .B1(new_n916), .B2(new_n904), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n947), .A2(new_n1158), .B1(new_n948), .B2(KEYINPUT40), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1159), .B2(new_n683), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n952), .A2(G330), .A3(new_n1156), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n939), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n920), .A2(new_n1160), .A3(new_n938), .A4(new_n1161), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1148), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n698), .B1(new_n1147), .B2(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1119), .A2(new_n1146), .B1(new_n1164), .B2(new_n1163), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(KEYINPUT57), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1157), .A2(new_n762), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n760), .B1(new_n835), .B2(G50), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n267), .A2(G41), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G50), .B(new_n1172), .C1(new_n281), .C2(new_n255), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n791), .A2(new_n471), .B1(new_n781), .B2(new_n539), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G116), .A2(new_n786), .B1(new_n789), .B2(G58), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n394), .B2(new_n780), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1174), .B(new_n1176), .C1(G68), .C2(new_n801), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1172), .B1(new_n230), .B2(new_n793), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT120), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n798), .A2(G283), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1177), .B(new_n1180), .C1(new_n1179), .C2(new_n1178), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT58), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1173), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n798), .A2(G124), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G33), .B(G41), .C1(new_n789), .C2(G159), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G125), .A2(new_n786), .B1(new_n808), .B2(G128), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT122), .B1(new_n793), .B2(new_n1137), .ZN(new_n1187));
  OR3_X1    g0987(.A1(new_n793), .A2(new_n1137), .A3(KEYINPUT122), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n791), .A2(new_n845), .B1(new_n780), .B2(new_n838), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT121), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1189), .B(new_n1191), .C1(G150), .C2(new_n801), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT59), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1184), .B(new_n1185), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1183), .B1(new_n1182), .B2(new_n1181), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1171), .B1(new_n1196), .B2(new_n768), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1169), .A2(new_n759), .B1(new_n1170), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1168), .A2(new_n1198), .ZN(G375));
  NAND2_X1  g0999(.A1(new_n942), .A2(new_n1103), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1102), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n980), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n1203), .A3(new_n1104), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n935), .A2(new_n762), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n760), .B1(new_n835), .B2(G68), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n791), .A2(new_n599), .B1(new_n788), .B2(new_n422), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n267), .B(new_n1207), .C1(G294), .C2(new_n786), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n798), .A2(G303), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n383), .A2(new_n780), .B1(new_n793), .B2(new_n471), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G283), .B2(new_n808), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1042), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n791), .A2(new_n1137), .B1(new_n785), .B2(new_n845), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G150), .B2(new_n817), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n798), .A2(G128), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n612), .B1(new_n789), .B2(G58), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G137), .A2(new_n808), .B1(new_n794), .B2(G159), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1013), .A2(new_n300), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1212), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1220), .A2(KEYINPUT123), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n769), .B1(new_n1220), .B2(KEYINPUT123), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1206), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1102), .A2(new_n759), .B1(new_n1205), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1204), .A2(new_n1224), .ZN(G381));
  NAND3_X1  g1025(.A1(new_n1204), .A2(new_n860), .A3(new_n1224), .ZN(new_n1226));
  OR3_X1    g1026(.A1(G390), .A2(new_n1226), .A3(G378), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n822), .B(new_n1059), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1227), .A2(G387), .A3(G375), .A4(new_n1228), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT124), .Z(G407));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(G343), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT125), .Z(new_n1234));
  NAND4_X1  g1034(.A1(new_n1168), .A2(new_n1231), .A3(new_n1198), .A4(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(G213), .A3(new_n1235), .ZN(G409));
  AOI21_X1  g1036(.A(new_n1200), .B1(new_n1121), .B2(new_n1117), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n920), .A2(new_n1160), .A3(new_n938), .A4(new_n1161), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n920), .A2(new_n938), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n697), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1147), .B2(new_n1169), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G378), .B(new_n1198), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT126), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT126), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1168), .A2(new_n1245), .A3(G378), .A4(new_n1198), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1167), .A2(new_n1203), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1198), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1231), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1233), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1104), .A2(KEYINPUT60), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1202), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1200), .A2(KEYINPUT60), .A3(new_n1201), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n697), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1224), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n860), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(G384), .A3(new_n1224), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1251), .A2(new_n1252), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1258), .A2(new_n1259), .B1(G2897), .B2(new_n1234), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1233), .A2(G2897), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1260), .A2(new_n1267), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1265), .A2(new_n1233), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1234), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(KEYINPUT63), .A3(new_n1261), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G387), .A2(new_n1090), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G393), .A2(G396), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1228), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n996), .A2(new_n1028), .A3(G390), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1272), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G390), .B1(new_n996), .B2(new_n1028), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1028), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1279), .B(new_n1090), .C1(new_n981), .C2(new_n995), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1274), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1277), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1264), .A2(new_n1269), .A3(new_n1271), .A4(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1268), .A2(new_n1266), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1282), .B1(new_n1270), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1262), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1270), .A2(KEYINPUT62), .A3(new_n1261), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1284), .B1(new_n1290), .B2(new_n1292), .ZN(G405));
  NAND2_X1  g1093(.A1(new_n1261), .A2(KEYINPUT127), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1244), .A2(new_n1246), .B1(new_n1231), .B2(G375), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1294), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1298), .A2(new_n1302), .ZN(G402));
endmodule


