//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n202), .B1(new_n208), .B2(KEYINPUT70), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(KEYINPUT70), .B2(new_n208), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(KEYINPUT71), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n203), .A2(new_n202), .A3(new_n207), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(KEYINPUT71), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G226gat), .ZN(new_n216));
  INV_X1    g015(.A(G233gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OR2_X1    g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n225));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n224), .A2(new_n225), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n225), .B2(new_n224), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n229), .A2(KEYINPUT66), .ZN(new_n231));
  AOI21_X1  g030(.A(G190gat), .B1(new_n231), .B2(KEYINPUT27), .ZN(new_n232));
  OR3_X1    g031(.A1(new_n229), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT28), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT27), .B(G183gat), .Z(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n235), .A2(new_n236), .A3(G190gat), .ZN(new_n237));
  OAI221_X1 g036(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n234), .C2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(new_n229), .B2(new_n230), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n240), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n220), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n239), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n250), .A2(new_n220), .A3(new_n247), .A4(new_n246), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n245), .A2(new_n249), .B1(new_n251), .B2(KEYINPUT25), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n238), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n238), .A2(KEYINPUT72), .A3(new_n252), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n219), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n253), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n218), .A2(KEYINPUT29), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n215), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n218), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n255), .A2(new_n256), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n214), .B(new_n263), .C1(new_n264), .C2(new_n260), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT37), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT83), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT83), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n265), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(KEYINPUT37), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n267), .B1(new_n262), .B2(new_n265), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT85), .ZN(new_n274));
  XOR2_X1   g073(.A(G8gat), .B(G36gat), .Z(new_n275));
  XNOR2_X1  g074(.A(G64gat), .B(G92gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  OR3_X1    g076(.A1(new_n273), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n274), .B1(new_n273), .B2(new_n277), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n272), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT38), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n282));
  XOR2_X1   g081(.A(G113gat), .B(G120gat), .Z(new_n283));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G134gat), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT68), .B1(new_n289), .B2(G127gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n285), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT2), .ZN(new_n295));
  INV_X1    g094(.A(G141gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(G148gat), .ZN(new_n297));
  INV_X1    g096(.A(G148gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(G141gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  INV_X1    g101(.A(G162gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n296), .B2(G148gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n298), .A2(KEYINPUT74), .A3(G141gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n307), .B(new_n308), .C1(G141gat), .C2(new_n298), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n301), .B1(new_n304), .B2(KEYINPUT2), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT4), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n315), .B(KEYINPUT76), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n305), .A2(new_n311), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n293), .B(new_n319), .C1(new_n322), .C2(new_n318), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n314), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n313), .B1(new_n322), .B2(new_n294), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n316), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(KEYINPUT77), .A3(new_n316), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n324), .A2(new_n329), .A3(KEYINPUT5), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G1gat), .B(G29gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT0), .ZN(new_n334));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n282), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n337), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT82), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n336), .B1(new_n325), .B2(new_n331), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT82), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(KEYINPUT6), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT84), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n277), .A2(KEYINPUT38), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n264), .A2(new_n260), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n218), .B2(new_n258), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n267), .B1(new_n350), .B2(new_n215), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n214), .B1(new_n257), .B2(new_n261), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n353), .A2(new_n272), .B1(new_n277), .B2(new_n266), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n281), .A2(new_n345), .A3(new_n347), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n314), .A2(new_n323), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n316), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n336), .B1(new_n357), .B2(KEYINPUT39), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT40), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT39), .B1(new_n326), .B2(new_n316), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n360), .B1(new_n356), .B2(new_n316), .ZN(new_n361));
  OR3_X1    g160(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n358), .B2(new_n361), .ZN(new_n363));
  AND4_X1   g162(.A1(new_n341), .A2(new_n344), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n262), .A2(new_n265), .A3(KEYINPUT30), .A4(new_n277), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n277), .B1(new_n262), .B2(new_n265), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n266), .A2(new_n277), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G22gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n374), .B(KEYINPUT78), .Z(new_n375));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n312), .B2(new_n318), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n211), .B2(new_n213), .ZN(new_n377));
  INV_X1    g176(.A(new_n202), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n208), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n212), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n312), .B1(new_n382), .B2(new_n318), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n375), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n319), .A2(new_n381), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n376), .A2(KEYINPUT79), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n214), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(G228gat), .A3(G233gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n211), .A2(new_n381), .A3(new_n213), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n322), .B1(new_n391), .B2(new_n318), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n373), .B(new_n384), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT31), .B(G50gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT81), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n384), .B1(new_n390), .B2(new_n392), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G22gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n393), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n405), .A3(new_n398), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n400), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n395), .B2(new_n398), .ZN(new_n408));
  INV_X1    g207(.A(new_n398), .ZN(new_n409));
  AOI211_X1 g208(.A(KEYINPUT81), .B(new_n409), .C1(new_n393), .C2(new_n394), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n403), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n364), .A2(new_n372), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n355), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n258), .A2(new_n293), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n253), .A2(new_n294), .ZN(new_n418));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT64), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n416), .B1(new_n421), .B2(KEYINPUT32), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n416), .A2(KEYINPUT69), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n416), .A2(KEYINPUT69), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(KEYINPUT33), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(KEYINPUT32), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n417), .A2(new_n418), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n419), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n420), .A2(KEYINPUT34), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n432), .A2(KEYINPUT34), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n425), .A2(new_n434), .A3(new_n429), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT36), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT36), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n436), .A2(new_n440), .A3(new_n437), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n407), .A2(new_n411), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n346), .B1(new_n338), .B2(new_n342), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(new_n367), .A3(new_n371), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n442), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n438), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT35), .B1(new_n449), .B2(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n347), .A2(new_n345), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT35), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n438), .B1(new_n407), .B2(new_n411), .ZN(new_n453));
  INV_X1    g252(.A(new_n372), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n413), .A2(new_n447), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT15), .ZN(new_n457));
  OR2_X1    g256(.A1(G43gat), .A2(G50gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(G43gat), .A2(G50gat), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G29gat), .ZN(new_n461));
  INV_X1    g260(.A(G36gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT14), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT14), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(G29gat), .B2(G36gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT86), .ZN(new_n466));
  NAND2_X1  g265(.A1(G29gat), .A2(G36gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT86), .B1(new_n463), .B2(new_n465), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n460), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(new_n465), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n457), .A3(new_n459), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n471), .A2(new_n473), .A3(new_n467), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(G1gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT16), .ZN(new_n478));
  INV_X1    g277(.A(G15gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G22gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n373), .A2(G15gat), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(G1gat), .B1(new_n480), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g282(.A(G8gat), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n485));
  INV_X1    g284(.A(G8gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(new_n486), .C1(G1gat), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT89), .B1(new_n476), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n466), .A3(new_n467), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n474), .A2(new_n465), .A3(new_n463), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n461), .A2(new_n462), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n460), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n493), .A2(new_n460), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n484), .A2(new_n488), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n476), .A2(new_n489), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n490), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n503), .B(KEYINPUT13), .Z(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT90), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  INV_X1    g307(.A(new_n503), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n470), .A2(KEYINPUT17), .A3(new_n475), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n511));
  OAI211_X1 g310(.A(new_n510), .B(new_n499), .C1(new_n497), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n476), .B2(new_n489), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n511), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n476), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n517), .A2(new_n513), .A3(new_n499), .A4(new_n510), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n509), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n506), .A2(new_n508), .B1(new_n519), .B2(KEYINPUT18), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(KEYINPUT18), .ZN(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G197gat), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT11), .B(G169gat), .Z(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT12), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n526), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT91), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n521), .B1(new_n520), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n506), .A2(new_n508), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n519), .A2(KEYINPUT18), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n532), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n529), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT92), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n537), .B(new_n529), .C1(new_n531), .C2(new_n534), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n528), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n456), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n445), .ZN(new_n541));
  AND2_X1   g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G57gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G64gat), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G57gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G71gat), .B(G78gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n546), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G127gat), .B(G155gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n560), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n499), .B1(new_n557), .B2(new_n556), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n565), .A2(new_n570), .A3(new_n566), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT7), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(G85gat), .A3(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n579), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n583), .B1(new_n579), .B2(new_n586), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n517), .A2(new_n510), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n579), .A2(new_n586), .ZN(new_n591));
  INV_X1    g390(.A(new_n583), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n579), .A2(new_n583), .A3(new_n586), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n476), .A2(new_n595), .B1(KEYINPUT41), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G190gat), .B(G218gat), .Z(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT94), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OR3_X1    g405(.A1(new_n600), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n600), .B2(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n574), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G120gat), .B(G148gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n589), .A2(new_n616), .A3(new_n556), .ZN(new_n617));
  INV_X1    g416(.A(new_n582), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(KEYINPUT96), .A3(new_n580), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n619), .A2(new_n579), .A3(new_n586), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(new_n579), .B2(new_n586), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n620), .A2(new_n556), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n547), .A2(new_n555), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n595), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n589), .A2(KEYINPUT95), .A3(new_n556), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n617), .B1(new_n627), .B2(new_n616), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT97), .Z(new_n630));
  NOR2_X1   g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n627), .A2(new_n629), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n615), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OR3_X1    g432(.A1(new_n620), .A2(new_n556), .A3(new_n621), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT95), .B1(new_n589), .B2(new_n556), .ZN(new_n635));
  AND4_X1   g434(.A1(KEYINPUT95), .A2(new_n556), .A3(new_n593), .A4(new_n594), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n634), .B(new_n616), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n617), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n629), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n640), .B(new_n614), .C1(new_n629), .C2(new_n627), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n611), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n540), .A2(new_n541), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g444(.A1(new_n540), .A2(new_n372), .A3(new_n643), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT16), .B(G8gat), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n648), .A2(KEYINPUT98), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n646), .A2(G8gat), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n648), .B1(new_n654), .B2(new_n649), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n650), .B1(new_n653), .B2(new_n655), .ZN(G1325gat));
  INV_X1    g455(.A(new_n540), .ZN(new_n657));
  INV_X1    g456(.A(new_n643), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n442), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n660), .A2(new_n479), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n479), .B1(new_n660), .B2(new_n438), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(G1326gat));
  NAND2_X1  g465(.A1(new_n659), .A2(new_n444), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n574), .A2(new_n642), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n610), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n540), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n541), .A2(new_n461), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT100), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n676));
  INV_X1    g475(.A(new_n674), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n540), .A2(new_n676), .A3(new_n672), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n456), .B2(new_n610), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n413), .A2(new_n447), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n450), .A2(new_n455), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(KEYINPUT44), .A3(new_n609), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n539), .A2(new_n671), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n541), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G29gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n675), .A2(KEYINPUT45), .A3(new_n678), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n681), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n681), .A2(KEYINPUT101), .A3(new_n691), .A4(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n673), .A2(G36gat), .A3(new_n454), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n688), .A2(new_n372), .A3(new_n689), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n462), .B2(new_n700), .ZN(G1329gat));
  NAND3_X1  g500(.A1(new_n688), .A2(new_n442), .A3(new_n689), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G43gat), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n673), .A2(G43gat), .A3(new_n438), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1330gat));
  NAND4_X1  g506(.A1(new_n683), .A2(new_n687), .A3(new_n444), .A4(new_n689), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT102), .B1(new_n708), .B2(G50gat), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n673), .A2(G50gat), .A3(new_n443), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(G50gat), .B2(new_n708), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n711), .B(new_n713), .ZN(G1331gat));
  INV_X1    g513(.A(new_n539), .ZN(new_n715));
  INV_X1    g514(.A(new_n642), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n715), .A2(new_n611), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n686), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n445), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT103), .B(G57gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1332gat));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n454), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  AND2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n722), .B2(new_n723), .ZN(G1333gat));
  NOR3_X1   g525(.A1(new_n718), .A2(G71gat), .A3(new_n438), .ZN(new_n727));
  INV_X1    g526(.A(new_n718), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n442), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(G71gat), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n444), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  INV_X1    g532(.A(new_n574), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n539), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT104), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n716), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n688), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n445), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n456), .A2(new_n610), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n738), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n686), .A2(new_n609), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n739), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT105), .B(KEYINPUT51), .Z(new_n749));
  OAI21_X1  g548(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n642), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n541), .A2(new_n584), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n742), .B1(new_n754), .B2(new_n755), .ZN(G1336gat));
  NOR3_X1   g555(.A1(new_n454), .A2(G92gat), .A3(new_n716), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n747), .A2(new_n739), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n758), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n743), .B2(new_n738), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n757), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n683), .A2(new_n687), .A3(new_n372), .A4(new_n740), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(KEYINPUT107), .A3(G92gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT107), .B1(new_n763), .B2(G92gat), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT52), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n688), .A2(KEYINPUT109), .A3(new_n372), .A4(new_n740), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n585), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(new_n750), .B2(new_n757), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n767), .B1(new_n774), .B2(new_n775), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n741), .B2(new_n661), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n438), .A2(G99gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n754), .B2(new_n778), .ZN(G1338gat));
  OR2_X1    g578(.A1(new_n759), .A2(new_n761), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n443), .A2(G106gat), .A3(new_n716), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT111), .Z(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n688), .A2(new_n444), .A3(new_n740), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n780), .A2(new_n783), .B1(new_n784), .B2(G106gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n784), .A2(G106gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n750), .A2(new_n783), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n786), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n785), .A2(new_n786), .B1(new_n787), .B2(new_n789), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n515), .A2(new_n509), .A3(new_n518), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n504), .B2(new_n502), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n525), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n527), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n642), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n637), .A2(new_n630), .A3(new_n638), .ZN(new_n798));
  INV_X1    g597(.A(new_n629), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n798), .B(KEYINPUT54), .C1(new_n628), .C2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n614), .B1(new_n631), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n640), .A2(KEYINPUT112), .A3(KEYINPUT54), .A4(new_n798), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n802), .A2(new_n804), .A3(new_n805), .A4(KEYINPUT55), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(new_n641), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n808), .B2(new_n810), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n797), .B1(new_n539), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n610), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n532), .A2(new_n533), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n526), .B1(new_n519), .B2(KEYINPUT18), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT114), .B(new_n794), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n609), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT115), .B1(new_n813), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n808), .A2(new_n810), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT113), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n820), .A2(new_n609), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT114), .B1(new_n527), .B2(new_n794), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n826), .A2(new_n829), .A3(new_n830), .A4(new_n807), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n822), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n574), .B1(new_n815), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n643), .A2(new_n539), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n791), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n822), .A2(new_n831), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n610), .B2(new_n814), .ZN(new_n838));
  OAI211_X1 g637(.A(KEYINPUT116), .B(new_n834), .C1(new_n838), .C2(new_n574), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n449), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n372), .A2(new_n445), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n715), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n642), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(G120gat), .ZN(G1341gat));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n574), .B1(new_n849), .B2(G127gat), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(G127gat), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(KEYINPUT118), .Z(new_n853));
  XNOR2_X1  g652(.A(new_n851), .B(new_n853), .ZN(G1342gat));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n841), .A2(new_n541), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n454), .A2(new_n609), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n289), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n855), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT119), .B(KEYINPUT56), .C1(new_n856), .C2(new_n859), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n841), .A2(new_n541), .A3(new_n858), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n860), .A2(new_n861), .B1(G134gat), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(G1343gat));
  NOR2_X1   g666(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n836), .A2(new_n444), .A3(new_n839), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n443), .A2(new_n871), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n807), .A2(new_n823), .ZN(new_n874));
  AOI22_X1  g673(.A1(new_n715), .A2(new_n874), .B1(new_n642), .B2(new_n796), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(new_n609), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n574), .B1(new_n876), .B2(new_n832), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n873), .B1(new_n877), .B2(new_n835), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n842), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n442), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n715), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G141gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n836), .A2(new_n839), .A3(new_n444), .A4(new_n881), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n539), .A2(G141gat), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n869), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n888), .B(new_n868), .C1(new_n882), .C2(G141gat), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(G1344gat));
  NAND2_X1  g691(.A1(new_n881), .A2(new_n642), .ZN(new_n893));
  OR3_X1    g692(.A1(new_n870), .A2(G148gat), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n834), .B(KEYINPUT121), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n875), .A2(new_n609), .B1(new_n813), .B2(new_n821), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n734), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n871), .B1(new_n898), .B2(new_n443), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n836), .A2(new_n839), .A3(new_n873), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n893), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n298), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n895), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n881), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n872), .B2(new_n878), .ZN(new_n907));
  AOI211_X1 g706(.A(KEYINPUT59), .B(new_n298), .C1(new_n907), .C2(new_n642), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n894), .B1(new_n905), .B2(new_n908), .ZN(G1345gat));
  NOR2_X1   g708(.A1(new_n885), .A2(new_n734), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT123), .ZN(new_n911));
  AOI21_X1  g710(.A(G155gat), .B1(new_n910), .B2(KEYINPUT123), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n734), .A2(new_n302), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n911), .A2(new_n912), .B1(new_n907), .B2(new_n913), .ZN(G1346gat));
  AND2_X1   g713(.A1(new_n907), .A2(new_n609), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n858), .A2(new_n303), .A3(new_n541), .A4(new_n661), .ZN(new_n916));
  OAI22_X1  g715(.A1(new_n915), .A2(new_n303), .B1(new_n870), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n454), .A2(new_n541), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n840), .A2(new_n449), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n715), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n642), .ZN(new_n923));
  XOR2_X1   g722(.A(KEYINPUT124), .B(G176gat), .Z(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(G1349gat));
  AND2_X1   g724(.A1(new_n836), .A2(new_n839), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n453), .A3(new_n918), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n229), .B1(new_n927), .B2(new_n734), .ZN(new_n928));
  OR2_X1    g727(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n920), .A2(new_n235), .A3(new_n574), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(G1350gat));
  NAND2_X1  g732(.A1(new_n920), .A2(new_n609), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n230), .B1(new_n935), .B2(KEYINPUT61), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(KEYINPUT126), .A3(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n934), .B(new_n936), .C1(new_n935), .C2(KEYINPUT61), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n939), .B(new_n940), .C1(G190gat), .C2(new_n934), .ZN(G1351gat));
  NAND2_X1  g740(.A1(new_n899), .A2(new_n900), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n919), .A2(new_n442), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(G197gat), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(new_n539), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n919), .A2(new_n443), .A3(new_n442), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n926), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n715), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n946), .A2(new_n950), .ZN(G1352gat));
  NOR3_X1   g750(.A1(new_n948), .A2(G204gat), .A3(new_n716), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT127), .B1(new_n944), .B2(new_n716), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G204gat), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n944), .A2(KEYINPUT127), .A3(new_n716), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1353gat));
  NAND3_X1  g756(.A1(new_n949), .A2(new_n205), .A3(new_n574), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n574), .A3(new_n943), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n944), .B2(new_n610), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n949), .A2(new_n206), .A3(new_n609), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


