

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(n717), .B(KEYINPUT29), .ZN(n718) );
  XNOR2_X1 U556 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U557 ( .A1(G651), .A2(n624), .ZN(n653) );
  NOR2_X1 U558 ( .A1(n541), .A2(n540), .ZN(G160) );
  NOR2_X1 U559 ( .A1(G543), .A2(G651), .ZN(n652) );
  NAND2_X1 U560 ( .A1(n652), .A2(G89), .ZN(n519) );
  XNOR2_X1 U561 ( .A(n519), .B(KEYINPUT4), .ZN(n521) );
  XOR2_X1 U562 ( .A(G543), .B(KEYINPUT0), .Z(n624) );
  INV_X1 U563 ( .A(G651), .ZN(n523) );
  NOR2_X1 U564 ( .A1(n624), .A2(n523), .ZN(n646) );
  NAND2_X1 U565 ( .A1(G76), .A2(n646), .ZN(n520) );
  NAND2_X1 U566 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U567 ( .A(n522), .B(KEYINPUT5), .ZN(n529) );
  NAND2_X1 U568 ( .A1(G51), .A2(n653), .ZN(n526) );
  NOR2_X1 U569 ( .A1(G543), .A2(n523), .ZN(n524) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n524), .Z(n649) );
  NAND2_X1 U571 ( .A1(G63), .A2(n649), .ZN(n525) );
  NAND2_X1 U572 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U573 ( .A(KEYINPUT6), .B(n527), .Z(n528) );
  NAND2_X1 U574 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U575 ( .A(n530), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U576 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U577 ( .A(G2105), .ZN(n532) );
  NOR2_X2 U578 ( .A1(G2104), .A2(n532), .ZN(n874) );
  NAND2_X1 U579 ( .A1(G125), .A2(n874), .ZN(n531) );
  XNOR2_X1 U580 ( .A(n531), .B(KEYINPUT64), .ZN(n535) );
  AND2_X1 U581 ( .A1(n532), .A2(G2104), .ZN(n879) );
  NAND2_X1 U582 ( .A1(G101), .A2(n879), .ZN(n533) );
  XOR2_X1 U583 ( .A(KEYINPUT23), .B(n533), .Z(n534) );
  NAND2_X1 U584 ( .A1(n535), .A2(n534), .ZN(n541) );
  XNOR2_X1 U585 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n537) );
  NOR2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n537), .B(n536), .ZN(n878) );
  NAND2_X1 U588 ( .A1(G137), .A2(n878), .ZN(n539) );
  AND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n875) );
  NAND2_X1 U590 ( .A1(G113), .A2(n875), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U592 ( .A1(G52), .A2(n653), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G64), .A2(n649), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U595 ( .A1(G77), .A2(n646), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G90), .A2(n652), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U599 ( .A1(n548), .A2(n547), .ZN(G171) );
  XOR2_X1 U600 ( .A(G2438), .B(G2454), .Z(n550) );
  XNOR2_X1 U601 ( .A(G2435), .B(G2430), .ZN(n549) );
  XNOR2_X1 U602 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U603 ( .A(n551), .B(G2427), .Z(n553) );
  XNOR2_X1 U604 ( .A(G1341), .B(G1348), .ZN(n552) );
  XNOR2_X1 U605 ( .A(n553), .B(n552), .ZN(n557) );
  XOR2_X1 U606 ( .A(G2443), .B(G2446), .Z(n555) );
  XNOR2_X1 U607 ( .A(KEYINPUT104), .B(G2451), .ZN(n554) );
  XNOR2_X1 U608 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U609 ( .A(n557), .B(n556), .Z(n558) );
  AND2_X1 U610 ( .A1(G14), .A2(n558), .ZN(G401) );
  AND2_X1 U611 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U612 ( .A(G82), .ZN(G220) );
  NAND2_X1 U613 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U614 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U615 ( .A(G223), .ZN(n821) );
  NAND2_X1 U616 ( .A1(n821), .A2(G567), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n560), .B(KEYINPUT11), .ZN(n561) );
  XNOR2_X1 U618 ( .A(KEYINPUT71), .B(n561), .ZN(G234) );
  XOR2_X1 U619 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n563) );
  NAND2_X1 U620 ( .A1(G56), .A2(n649), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n563), .B(n562), .ZN(n569) );
  NAND2_X1 U622 ( .A1(n652), .A2(G81), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G68), .A2(n646), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(n567), .Z(n568) );
  NOR2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U628 ( .A1(n653), .A2(G43), .ZN(n570) );
  NAND2_X1 U629 ( .A1(n571), .A2(n570), .ZN(n977) );
  INV_X1 U630 ( .A(G860), .ZN(n616) );
  OR2_X1 U631 ( .A1(n977), .A2(n616), .ZN(G153) );
  XNOR2_X1 U632 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G868), .A2(G301), .ZN(n572) );
  XNOR2_X1 U634 ( .A(n572), .B(KEYINPUT74), .ZN(n582) );
  INV_X1 U635 ( .A(G868), .ZN(n597) );
  NAND2_X1 U636 ( .A1(G92), .A2(n652), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G66), .A2(n649), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U639 ( .A1(G79), .A2(n646), .ZN(n576) );
  NAND2_X1 U640 ( .A1(G54), .A2(n653), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT75), .B(n577), .Z(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT15), .B(n580), .ZN(n960) );
  NAND2_X1 U645 ( .A1(n597), .A2(n960), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT76), .B(n583), .ZN(G284) );
  NAND2_X1 U648 ( .A1(G78), .A2(n646), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G91), .A2(n652), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U651 ( .A1(G53), .A2(n653), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G65), .A2(n649), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U654 ( .A(KEYINPUT67), .B(n588), .Z(n589) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n961) );
  XOR2_X1 U656 ( .A(n961), .B(KEYINPUT68), .Z(G299) );
  NOR2_X1 U657 ( .A1(G299), .A2(G868), .ZN(n592) );
  NOR2_X1 U658 ( .A1(G286), .A2(n597), .ZN(n591) );
  NOR2_X1 U659 ( .A1(n592), .A2(n591), .ZN(G297) );
  NAND2_X1 U660 ( .A1(G559), .A2(n616), .ZN(n593) );
  XOR2_X1 U661 ( .A(KEYINPUT77), .B(n593), .Z(n594) );
  INV_X1 U662 ( .A(n960), .ZN(n614) );
  NAND2_X1 U663 ( .A1(n594), .A2(n614), .ZN(n595) );
  XNOR2_X1 U664 ( .A(n595), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U665 ( .A1(G868), .A2(n977), .ZN(n596) );
  XNOR2_X1 U666 ( .A(KEYINPUT78), .B(n596), .ZN(n602) );
  NOR2_X1 U667 ( .A1(n960), .A2(n597), .ZN(n598) );
  XNOR2_X1 U668 ( .A(n598), .B(KEYINPUT79), .ZN(n599) );
  NOR2_X1 U669 ( .A1(G559), .A2(n599), .ZN(n600) );
  XNOR2_X1 U670 ( .A(KEYINPUT80), .B(n600), .ZN(n601) );
  NOR2_X1 U671 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G123), .A2(n874), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT18), .B(n603), .Z(n604) );
  XNOR2_X1 U674 ( .A(n604), .B(KEYINPUT81), .ZN(n606) );
  NAND2_X1 U675 ( .A1(G111), .A2(n875), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U677 ( .A1(G135), .A2(n878), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G99), .A2(n879), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n936) );
  XNOR2_X1 U681 ( .A(n936), .B(G2096), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT82), .ZN(n613) );
  INV_X1 U683 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U685 ( .A1(G559), .A2(n614), .ZN(n615) );
  XOR2_X1 U686 ( .A(n977), .B(n615), .Z(n665) );
  NAND2_X1 U687 ( .A1(n616), .A2(n665), .ZN(n623) );
  NAND2_X1 U688 ( .A1(G55), .A2(n653), .ZN(n618) );
  NAND2_X1 U689 ( .A1(G67), .A2(n649), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U691 ( .A1(G80), .A2(n646), .ZN(n620) );
  NAND2_X1 U692 ( .A1(G93), .A2(n652), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n667) );
  XOR2_X1 U695 ( .A(n623), .B(n667), .Z(G145) );
  NAND2_X1 U696 ( .A1(n624), .A2(G87), .ZN(n629) );
  NAND2_X1 U697 ( .A1(G49), .A2(n653), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U700 ( .A1(n649), .A2(n627), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U702 ( .A(KEYINPUT83), .B(n630), .Z(G288) );
  NAND2_X1 U703 ( .A1(G88), .A2(n652), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G50), .A2(n653), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n638) );
  NAND2_X1 U706 ( .A1(G62), .A2(n649), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(KEYINPUT86), .ZN(n636) );
  NAND2_X1 U708 ( .A1(G75), .A2(n646), .ZN(n634) );
  XOR2_X1 U709 ( .A(KEYINPUT87), .B(n634), .Z(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U711 ( .A1(n638), .A2(n637), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G72), .A2(n646), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G85), .A2(n652), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U715 ( .A1(G60), .A2(n649), .ZN(n641) );
  XOR2_X1 U716 ( .A(KEYINPUT66), .B(n641), .Z(n642) );
  NOR2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n653), .A2(G47), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G73), .A2(n646), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(KEYINPUT2), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n648), .B(KEYINPUT84), .ZN(n651) );
  NAND2_X1 U723 ( .A1(G61), .A2(n649), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U725 ( .A1(G86), .A2(n652), .ZN(n655) );
  NAND2_X1 U726 ( .A1(G48), .A2(n653), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT85), .B(n658), .ZN(G305) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(KEYINPUT88), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n659), .B(n667), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(G288), .ZN(n663) );
  XNOR2_X1 U733 ( .A(G166), .B(G299), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n661), .B(G290), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n664), .B(G305), .ZN(n890) );
  XNOR2_X1 U737 ( .A(n665), .B(n890), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n666), .A2(G868), .ZN(n669) );
  OR2_X1 U739 ( .A1(G868), .A2(n667), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U748 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  NAND2_X1 U749 ( .A1(G108), .A2(G120), .ZN(n674) );
  NOR2_X1 U750 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U751 ( .A1(G69), .A2(n675), .ZN(n901) );
  NAND2_X1 U752 ( .A1(n901), .A2(G567), .ZN(n680) );
  NOR2_X1 U753 ( .A1(G219), .A2(G220), .ZN(n676) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U755 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U756 ( .A1(G96), .A2(n678), .ZN(n902) );
  NAND2_X1 U757 ( .A1(n902), .A2(G2106), .ZN(n679) );
  NAND2_X1 U758 ( .A1(n680), .A2(n679), .ZN(n826) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U760 ( .A1(n826), .A2(n681), .ZN(n825) );
  NAND2_X1 U761 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U762 ( .A1(n878), .A2(G138), .ZN(n684) );
  NAND2_X1 U763 ( .A1(G126), .A2(n874), .ZN(n682) );
  XOR2_X1 U764 ( .A(KEYINPUT89), .B(n682), .Z(n683) );
  NAND2_X1 U765 ( .A1(n684), .A2(n683), .ZN(n688) );
  NAND2_X1 U766 ( .A1(G102), .A2(n879), .ZN(n686) );
  NAND2_X1 U767 ( .A1(G114), .A2(n875), .ZN(n685) );
  NAND2_X1 U768 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U769 ( .A1(n688), .A2(n687), .ZN(G164) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n771) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n770) );
  INV_X1 U773 ( .A(n770), .ZN(n689) );
  NAND2_X1 U774 ( .A1(n771), .A2(n689), .ZN(n740) );
  NAND2_X1 U775 ( .A1(G8), .A2(n740), .ZN(n766) );
  NOR2_X1 U776 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NAND2_X1 U777 ( .A1(n751), .A2(KEYINPUT33), .ZN(n690) );
  NOR2_X1 U778 ( .A1(n766), .A2(n690), .ZN(n756) );
  NOR2_X1 U779 ( .A1(n740), .A2(G2084), .ZN(n691) );
  XNOR2_X1 U780 ( .A(n691), .B(KEYINPUT95), .ZN(n723) );
  INV_X1 U781 ( .A(n723), .ZN(n692) );
  NAND2_X1 U782 ( .A1(G8), .A2(n692), .ZN(n738) );
  XNOR2_X1 U783 ( .A(G2078), .B(KEYINPUT25), .ZN(n903) );
  NOR2_X1 U784 ( .A1(n740), .A2(n903), .ZN(n694) );
  INV_X1 U785 ( .A(n740), .ZN(n705) );
  INV_X1 U786 ( .A(G1961), .ZN(n984) );
  NOR2_X1 U787 ( .A1(n705), .A2(n984), .ZN(n693) );
  NOR2_X1 U788 ( .A1(n694), .A2(n693), .ZN(n727) );
  NAND2_X1 U789 ( .A1(G171), .A2(n727), .ZN(n721) );
  NAND2_X1 U790 ( .A1(G1956), .A2(n740), .ZN(n695) );
  XNOR2_X1 U791 ( .A(KEYINPUT97), .B(n695), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n705), .A2(G2072), .ZN(n696) );
  XNOR2_X1 U793 ( .A(KEYINPUT27), .B(n696), .ZN(n697) );
  NOR2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n700) );
  NOR2_X1 U795 ( .A1(n961), .A2(n700), .ZN(n699) );
  XOR2_X1 U796 ( .A(n699), .B(KEYINPUT28), .Z(n716) );
  NAND2_X1 U797 ( .A1(n961), .A2(n700), .ZN(n714) );
  INV_X1 U798 ( .A(G1996), .ZN(n904) );
  NOR2_X1 U799 ( .A1(n740), .A2(n904), .ZN(n701) );
  XOR2_X1 U800 ( .A(n701), .B(KEYINPUT26), .Z(n703) );
  NAND2_X1 U801 ( .A1(n740), .A2(G1341), .ZN(n702) );
  NAND2_X1 U802 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U803 ( .A1(n977), .A2(n704), .ZN(n709) );
  NAND2_X1 U804 ( .A1(G1348), .A2(n740), .ZN(n707) );
  NAND2_X1 U805 ( .A1(G2067), .A2(n705), .ZN(n706) );
  NAND2_X1 U806 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U807 ( .A1(n960), .A2(n710), .ZN(n708) );
  OR2_X1 U808 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n960), .A2(n710), .ZN(n711) );
  NAND2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U811 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n719) );
  XNOR2_X1 U813 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n734) );
  NOR2_X1 U815 ( .A1(n766), .A2(G1966), .ZN(n722) );
  XNOR2_X1 U816 ( .A(n722), .B(KEYINPUT96), .ZN(n735) );
  NAND2_X1 U817 ( .A1(G8), .A2(n723), .ZN(n724) );
  NOR2_X1 U818 ( .A1(n735), .A2(n724), .ZN(n725) );
  XOR2_X1 U819 ( .A(KEYINPUT30), .B(n725), .Z(n726) );
  NOR2_X1 U820 ( .A1(G168), .A2(n726), .ZN(n730) );
  NOR2_X1 U821 ( .A1(G171), .A2(n727), .ZN(n728) );
  XNOR2_X1 U822 ( .A(KEYINPUT100), .B(n728), .ZN(n729) );
  NOR2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n732) );
  XNOR2_X1 U824 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n731) );
  XNOR2_X1 U825 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U826 ( .A1(n734), .A2(n733), .ZN(n739) );
  INV_X1 U827 ( .A(n739), .ZN(n736) );
  NOR2_X1 U828 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n749) );
  NAND2_X1 U830 ( .A1(n739), .A2(G286), .ZN(n745) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n766), .ZN(n742) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U834 ( .A1(n743), .A2(G303), .ZN(n744) );
  NAND2_X1 U835 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U836 ( .A1(G8), .A2(n746), .ZN(n747) );
  XNOR2_X1 U837 ( .A(KEYINPUT32), .B(n747), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n760) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n968) );
  NAND2_X1 U841 ( .A1(n760), .A2(n968), .ZN(n752) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n964) );
  NAND2_X1 U843 ( .A1(n752), .A2(n964), .ZN(n753) );
  NOR2_X1 U844 ( .A1(n753), .A2(n766), .ZN(n754) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n754), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n957) );
  NAND2_X1 U848 ( .A1(n757), .A2(n957), .ZN(n763) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U850 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U852 ( .A1(n761), .A2(n766), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n769) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U855 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  NOR2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U857 ( .A(n767), .B(KEYINPUT94), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n802) );
  NOR2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n816) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(KEYINPUT90), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G140), .A2(n878), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G104), .A2(n879), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U864 ( .A(n775), .B(n774), .ZN(n781) );
  XNOR2_X1 U865 ( .A(KEYINPUT35), .B(KEYINPUT91), .ZN(n779) );
  NAND2_X1 U866 ( .A1(G128), .A2(n874), .ZN(n777) );
  NAND2_X1 U867 ( .A1(G116), .A2(n875), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U869 ( .A(n779), .B(n778), .ZN(n780) );
  NOR2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U871 ( .A(n782), .B(KEYINPUT36), .ZN(n862) );
  XNOR2_X1 U872 ( .A(KEYINPUT37), .B(G2067), .ZN(n814) );
  NOR2_X1 U873 ( .A1(n862), .A2(n814), .ZN(n949) );
  NAND2_X1 U874 ( .A1(n816), .A2(n949), .ZN(n811) );
  NAND2_X1 U875 ( .A1(G119), .A2(n874), .ZN(n784) );
  NAND2_X1 U876 ( .A1(G131), .A2(n878), .ZN(n783) );
  NAND2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G95), .A2(n879), .ZN(n786) );
  NAND2_X1 U879 ( .A1(G107), .A2(n875), .ZN(n785) );
  NAND2_X1 U880 ( .A1(n786), .A2(n785), .ZN(n787) );
  OR2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n854) );
  NAND2_X1 U882 ( .A1(G1991), .A2(n854), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G129), .A2(n874), .ZN(n790) );
  NAND2_X1 U884 ( .A1(G117), .A2(n875), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n879), .A2(G105), .ZN(n791) );
  XOR2_X1 U887 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U889 ( .A(n794), .B(KEYINPUT92), .ZN(n796) );
  NAND2_X1 U890 ( .A1(G141), .A2(n878), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n856) );
  NAND2_X1 U892 ( .A1(G1996), .A2(n856), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n932) );
  NAND2_X1 U894 ( .A1(n932), .A2(n816), .ZN(n799) );
  XNOR2_X1 U895 ( .A(n799), .B(KEYINPUT93), .ZN(n808) );
  INV_X1 U896 ( .A(n808), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n811), .A2(n800), .ZN(n801) );
  NOR2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n804) );
  XNOR2_X1 U899 ( .A(G1986), .B(G290), .ZN(n970) );
  NAND2_X1 U900 ( .A1(n970), .A2(n816), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n819) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n856), .ZN(n945) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n854), .ZN(n937) );
  NOR2_X1 U905 ( .A1(n805), .A2(n937), .ZN(n806) );
  XNOR2_X1 U906 ( .A(n806), .B(KEYINPUT102), .ZN(n807) );
  NOR2_X1 U907 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n945), .A2(n809), .ZN(n810) );
  XNOR2_X1 U909 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U911 ( .A(KEYINPUT103), .B(n813), .Z(n815) );
  NAND2_X1 U912 ( .A1(n862), .A2(n814), .ZN(n931) );
  NAND2_X1 U913 ( .A1(n815), .A2(n931), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U919 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n823) );
  XOR2_X1 U921 ( .A(KEYINPUT105), .B(n823), .Z(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U923 ( .A(n826), .ZN(G319) );
  XOR2_X1 U924 ( .A(G2096), .B(KEYINPUT43), .Z(n828) );
  XNOR2_X1 U925 ( .A(G2072), .B(KEYINPUT106), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U927 ( .A(n829), .B(G2678), .Z(n831) );
  XNOR2_X1 U928 ( .A(G2067), .B(G2090), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U930 ( .A(KEYINPUT42), .B(G2100), .Z(n833) );
  XNOR2_X1 U931 ( .A(G2078), .B(G2084), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(G227) );
  XOR2_X1 U934 ( .A(G1956), .B(G1961), .Z(n837) );
  XNOR2_X1 U935 ( .A(G1976), .B(G1966), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U937 ( .A(n838), .B(G2474), .Z(n840) );
  XNOR2_X1 U938 ( .A(G1986), .B(G1971), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U940 ( .A(KEYINPUT41), .B(G1981), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(G229) );
  NAND2_X1 U944 ( .A1(G124), .A2(n874), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n845), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U946 ( .A1(G100), .A2(n879), .ZN(n846) );
  XOR2_X1 U947 ( .A(KEYINPUT107), .B(n846), .Z(n847) );
  NAND2_X1 U948 ( .A1(n848), .A2(n847), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G136), .A2(n878), .ZN(n850) );
  NAND2_X1 U950 ( .A1(G112), .A2(n875), .ZN(n849) );
  NAND2_X1 U951 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U952 ( .A1(n852), .A2(n851), .ZN(G162) );
  XOR2_X1 U953 ( .A(G164), .B(n936), .Z(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U955 ( .A(G160), .B(G162), .Z(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n864) );
  XOR2_X1 U958 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n860) );
  XNOR2_X1 U959 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n887) );
  NAND2_X1 U963 ( .A1(n879), .A2(G103), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n865), .B(KEYINPUT108), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G139), .A2(n878), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U967 ( .A(KEYINPUT109), .B(n868), .Z(n873) );
  NAND2_X1 U968 ( .A1(G127), .A2(n874), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G115), .A2(n875), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n871), .Z(n872) );
  NOR2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n926) );
  NAND2_X1 U973 ( .A1(G130), .A2(n874), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G118), .A2(n875), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U976 ( .A1(G142), .A2(n878), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G106), .A2(n879), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U979 ( .A(KEYINPUT45), .B(n882), .Z(n883) );
  NOR2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n926), .B(n885), .ZN(n886) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U983 ( .A1(G37), .A2(n888), .ZN(G395) );
  XOR2_X1 U984 ( .A(n977), .B(n960), .Z(n889) );
  XOR2_X1 U985 ( .A(n889), .B(KEYINPUT112), .Z(n892) );
  XNOR2_X1 U986 ( .A(G171), .B(n890), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U988 ( .A(G286), .B(n893), .Z(n894) );
  NOR2_X1 U989 ( .A1(G37), .A2(n894), .ZN(G397) );
  NOR2_X1 U990 ( .A1(G227), .A2(G229), .ZN(n895) );
  XOR2_X1 U991 ( .A(KEYINPUT49), .B(n895), .Z(n896) );
  NAND2_X1 U992 ( .A1(G319), .A2(n896), .ZN(n897) );
  NOR2_X1 U993 ( .A1(G401), .A2(n897), .ZN(n900) );
  NOR2_X1 U994 ( .A1(G395), .A2(G397), .ZN(n898) );
  XOR2_X1 U995 ( .A(KEYINPUT113), .B(n898), .Z(n899) );
  NAND2_X1 U996 ( .A1(n900), .A2(n899), .ZN(G225) );
  XOR2_X1 U997 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U999 ( .A(G120), .ZN(G236) );
  INV_X1 U1000 ( .A(G108), .ZN(G238) );
  INV_X1 U1001 ( .A(G96), .ZN(G221) );
  INV_X1 U1002 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1003 ( .A1(n902), .A2(n901), .ZN(G325) );
  INV_X1 U1004 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1005 ( .A(G27), .B(n903), .ZN(n912) );
  XOR2_X1 U1006 ( .A(G2067), .B(G26), .Z(n906) );
  XNOR2_X1 U1007 ( .A(n904), .B(G32), .ZN(n905) );
  NAND2_X1 U1008 ( .A1(n906), .A2(n905), .ZN(n910) );
  XOR2_X1 U1009 ( .A(G1991), .B(G25), .Z(n907) );
  NAND2_X1 U1010 ( .A1(n907), .A2(G28), .ZN(n908) );
  XNOR2_X1 U1011 ( .A(KEYINPUT120), .B(n908), .ZN(n909) );
  NOR2_X1 U1012 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(G33), .B(G2072), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1016 ( .A(KEYINPUT53), .B(n915), .Z(n919) );
  XNOR2_X1 U1017 ( .A(KEYINPUT54), .B(G34), .ZN(n916) );
  XNOR2_X1 U1018 ( .A(n916), .B(KEYINPUT121), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(G2084), .B(n917), .ZN(n918) );
  NAND2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(G35), .B(G2090), .ZN(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n922), .A2(KEYINPUT55), .ZN(n1016) );
  INV_X1 U1024 ( .A(n922), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(G29), .A2(KEYINPUT55), .ZN(n923) );
  NAND2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(G11), .A2(n925), .ZN(n1014) );
  INV_X1 U1028 ( .A(KEYINPUT55), .ZN(n955) );
  XOR2_X1 U1029 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1032 ( .A(KEYINPUT50), .B(n929), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(n930), .B(KEYINPUT118), .ZN(n935) );
  INV_X1 U1034 ( .A(n931), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n943) );
  XOR2_X1 U1037 ( .A(G160), .B(G2084), .Z(n940) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(KEYINPUT115), .B(n938), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1041 ( .A(KEYINPUT116), .B(n941), .Z(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n951) );
  XOR2_X1 U1043 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1045 ( .A(KEYINPUT117), .B(n946), .Z(n947) );
  XNOR2_X1 U1046 ( .A(n947), .B(KEYINPUT51), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(n952), .B(KEYINPUT52), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(KEYINPUT119), .B(n953), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n956), .A2(G29), .ZN(n1012) );
  XNOR2_X1 U1053 ( .A(G16), .B(KEYINPUT56), .ZN(n983) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(n959), .B(KEYINPUT57), .ZN(n981) );
  XNOR2_X1 U1057 ( .A(G171), .B(G1961), .ZN(n975) );
  XNOR2_X1 U1058 ( .A(n960), .B(G1348), .ZN(n973) );
  XOR2_X1 U1059 ( .A(n961), .B(G1956), .Z(n962) );
  XNOR2_X1 U1060 ( .A(KEYINPUT122), .B(n962), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(G1971), .A2(G303), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(KEYINPUT123), .B(n971), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT124), .B(n976), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G1341), .B(n977), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n1009) );
  INV_X1 U1074 ( .A(G16), .ZN(n1007) );
  XNOR2_X1 U1075 ( .A(G5), .B(n984), .ZN(n1002) );
  XNOR2_X1 U1076 ( .A(G1981), .B(G6), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n985), .B(G4), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n986), .B(G1348), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G1341), .B(G19), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(G1956), .B(G20), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(n993), .B(KEYINPUT60), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G1976), .B(G23), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n997) );
  XOR2_X1 U1089 ( .A(G1986), .B(G24), .Z(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT58), .B(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G21), .B(G1966), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1099 ( .A(KEYINPUT126), .B(n1010), .Z(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(n1017), .B(KEYINPUT127), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1018), .ZN(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

