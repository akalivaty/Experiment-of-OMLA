//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT66), .B(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n209), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n207), .ZN(new_n225));
  NOR2_X1   g0025(.A1(G58), .A2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n219), .B(new_n223), .C1(new_n225), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT68), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n235), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  AND2_X1   g0048(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n224), .B1(new_n248), .B2(KEYINPUT70), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT7), .B1(new_n254), .B2(new_n207), .ZN(new_n257));
  OAI21_X1  g0057(.A(G68), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT16), .ZN(new_n259));
  INV_X1    g0059(.A(G58), .ZN(new_n260));
  INV_X1    g0060(.A(G68), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(G20), .B1(new_n262), .B2(new_n226), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G159), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n258), .A2(new_n259), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT7), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n269), .B1(new_n274), .B2(G20), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n261), .B1(new_n275), .B2(new_n255), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT16), .B1(new_n276), .B2(new_n266), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n251), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n280), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n224), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n206), .A2(G13), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n207), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  OR3_X1    g0086(.A1(new_n207), .A2(KEYINPUT71), .A3(G1), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT71), .B1(new_n207), .B2(G1), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n285), .A2(new_n289), .B1(new_n286), .B2(new_n284), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n278), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n274), .A2(G223), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n274), .A2(G226), .A3(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G87), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  OAI211_X1 g0098(.A(G1), .B(G13), .C1(new_n271), .C2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G274), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n299), .A2(new_n302), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n305), .B1(new_n307), .B2(G232), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(G190), .B2(new_n309), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT17), .B1(new_n292), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n301), .A2(new_n315), .A3(new_n308), .ZN(new_n316));
  AOI21_X1  g0116(.A(G169), .B1(new_n301), .B2(new_n308), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT18), .B1(new_n292), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT18), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n318), .B(new_n321), .C1(new_n291), .C2(new_n278), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n292), .A2(KEYINPUT17), .A3(new_n312), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n314), .A2(new_n320), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n274), .A2(G238), .A3(G1698), .ZN(new_n325));
  INV_X1    g0125(.A(G107), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n274), .A2(new_n293), .ZN(new_n327));
  INV_X1    g0127(.A(G232), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n325), .B1(new_n326), .B2(new_n274), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n300), .ZN(new_n330));
  INV_X1    g0130(.A(new_n210), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n305), .B1(new_n307), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT72), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT72), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n334), .A2(new_n310), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(G190), .B1(new_n334), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n287), .A2(new_n288), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n285), .A2(G77), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT73), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT15), .B(G87), .Z(new_n344));
  NOR2_X1   g0144(.A1(new_n271), .A2(G20), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n344), .A2(new_n345), .B1(G20), .B2(G77), .ZN(new_n346));
  INV_X1    g0146(.A(new_n264), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n286), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n282), .B1(new_n211), .B2(new_n284), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n339), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n350), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n334), .A2(new_n336), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G179), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n334), .A2(G169), .A3(new_n336), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n324), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT69), .B(G226), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n304), .B1(new_n306), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n274), .A2(G223), .A3(G1698), .ZN(new_n362));
  INV_X1    g0162(.A(G222), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n362), .B1(new_n211), .B2(new_n274), .C1(new_n327), .C2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n361), .B1(new_n364), .B2(new_n300), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(G179), .B2(new_n365), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n203), .A2(G20), .ZN(new_n369));
  INV_X1    g0169(.A(new_n345), .ZN(new_n370));
  INV_X1    g0170(.A(G150), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n286), .A2(new_n370), .B1(new_n371), .B2(new_n347), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n251), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n284), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n251), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n340), .A2(G50), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n376), .A2(new_n377), .B1(G50), .B2(new_n375), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n368), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(KEYINPUT75), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n374), .B2(new_n378), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT9), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(KEYINPUT9), .A3(new_n383), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n365), .A2(G190), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n310), .B2(new_n365), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT10), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n384), .B2(new_n385), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT10), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(new_n387), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n380), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT77), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n299), .A2(G238), .A3(new_n302), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n304), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(G226), .B(new_n293), .C1(new_n252), .C2(new_n253), .ZN(new_n402));
  OAI211_X1 g0202(.A(G232), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n300), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n398), .A2(new_n304), .A3(KEYINPUT76), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n401), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT13), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n401), .A2(new_n406), .A3(new_n410), .A4(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G190), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n397), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n409), .A2(KEYINPUT77), .A3(G190), .A4(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n283), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(G20), .A3(new_n261), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(KEYINPUT12), .ZN(new_n419));
  OR2_X1    g0219(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n420));
  NAND2_X1  g0220(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n419), .B1(KEYINPUT79), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(KEYINPUT79), .B2(new_n422), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n264), .A2(G50), .B1(G20), .B2(new_n261), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n370), .B2(new_n211), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n282), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT11), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n285), .A2(G68), .A3(new_n340), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n424), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n412), .B2(G200), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n416), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n409), .A2(G179), .A3(new_n411), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n366), .B1(new_n409), .B2(new_n411), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI211_X1 g0236(.A(KEYINPUT14), .B(new_n366), .C1(new_n409), .C2(new_n411), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT74), .B1(new_n351), .B2(new_n356), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n359), .A2(new_n396), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n206), .A2(G45), .ZN(new_n443));
  OR2_X1    g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  NAND2_X1  g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G274), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n300), .A2(new_n446), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(G270), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n274), .A2(G264), .A3(G1698), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n274), .A2(G257), .A3(new_n293), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n254), .A2(G303), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n300), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G169), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  INV_X1    g0258(.A(G97), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n458), .B(new_n207), .C1(G33), .C2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT83), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G20), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n282), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n461), .B1(new_n282), .B2(new_n463), .ZN(new_n465));
  OAI211_X1 g0265(.A(KEYINPUT20), .B(new_n460), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n463), .B1(new_n249), .B2(new_n250), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT83), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n282), .A2(new_n461), .A3(new_n463), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(KEYINPUT84), .A3(KEYINPUT20), .A4(new_n460), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT20), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n468), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n375), .A2(G116), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n271), .A2(G1), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n376), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n480), .B2(G116), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n457), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n482), .A2(KEYINPUT86), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT21), .B1(new_n482), .B2(KEYINPUT86), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n454), .A2(new_n300), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n449), .A2(G270), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n447), .ZN(new_n488));
  OAI211_X1 g0288(.A(KEYINPUT21), .B(G169), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n450), .A2(G179), .A3(new_n455), .ZN(new_n490));
  AOI221_X4 g0290(.A(KEYINPUT85), .B1(new_n489), .B2(new_n490), .C1(new_n477), .C2(new_n481), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT85), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n477), .A2(new_n481), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n490), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n456), .A2(new_n310), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(G190), .B2(new_n456), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(new_n477), .A3(new_n481), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n485), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n274), .A2(G250), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n293), .B1(new_n501), .B2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(G1698), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(G244), .C1(new_n253), .C2(new_n252), .ZN(new_n505));
  INV_X1    g0305(.A(G244), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n272), .B2(new_n273), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n505), .B(new_n458), .C1(new_n507), .C2(KEYINPUT4), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n300), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n448), .B1(G257), .B2(new_n449), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n366), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n509), .A2(new_n510), .A3(G179), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n375), .A2(G97), .ZN(new_n514));
  XNOR2_X1  g0314(.A(G97), .B(G107), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n516), .A2(new_n459), .A3(G107), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(G20), .B1(G77), .B2(new_n264), .ZN(new_n521));
  OAI21_X1  g0321(.A(G107), .B1(new_n256), .B2(new_n257), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n514), .B1(new_n523), .B2(new_n282), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n480), .A2(G97), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n512), .A2(new_n513), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n518), .B1(new_n516), .B2(new_n515), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n527), .A2(new_n207), .B1(new_n211), .B2(new_n347), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n326), .B1(new_n275), .B2(new_n255), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n282), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n514), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(G200), .B1(new_n509), .B2(new_n510), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n509), .A2(new_n510), .A3(new_n413), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT80), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n513), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n532), .B1(new_n538), .B2(new_n511), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT80), .ZN(new_n540));
  INV_X1    g0340(.A(new_n535), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n533), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n539), .B(new_n540), .C1(new_n542), .C2(new_n532), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n443), .A2(G250), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n300), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n274), .A2(G238), .A3(new_n293), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n274), .A2(G244), .A3(G1698), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n548), .C1(new_n271), .C2(new_n462), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n546), .B1(new_n549), .B2(new_n300), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT82), .B1(new_n551), .B2(new_n413), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT82), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n553), .A3(G190), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G87), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(new_n459), .A3(new_n326), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n557), .B(KEYINPUT81), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT19), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n207), .B1(new_n404), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n254), .A2(G20), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n562), .A2(G68), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n282), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n480), .A2(G87), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n375), .A2(new_n344), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n550), .A2(new_n310), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n344), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n285), .B1(G1), .B2(new_n271), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n566), .B(new_n569), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n550), .A2(G179), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n366), .B2(new_n550), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n555), .A2(new_n572), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n537), .A2(new_n543), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n574), .A2(new_n326), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n417), .A2(G20), .A3(new_n326), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n581), .B(KEYINPUT25), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n556), .A2(KEYINPUT87), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n274), .A2(new_n207), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT22), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT88), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n207), .B2(G107), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT23), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n588), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n274), .A2(KEYINPUT22), .A3(new_n207), .A4(new_n584), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n587), .A2(new_n594), .A3(KEYINPUT24), .A4(new_n595), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n596), .A2(new_n282), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n587), .A2(new_n594), .A3(new_n595), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT89), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  AND4_X1   g0401(.A1(KEYINPUT89), .A2(new_n600), .A3(new_n282), .A4(new_n596), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n583), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n274), .A2(G250), .A3(new_n293), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n274), .A2(G257), .A3(G1698), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G294), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n300), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n449), .A2(G264), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n447), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT90), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n607), .A2(new_n300), .B1(new_n449), .B2(G264), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT90), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n447), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(G169), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n315), .B2(new_n610), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n603), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n600), .A2(new_n282), .A3(new_n596), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT89), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n597), .A2(KEYINPUT89), .A3(new_n600), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(G190), .B1(new_n611), .B2(new_n614), .ZN(new_n623));
  AOI21_X1  g0423(.A(G200), .B1(new_n612), .B2(new_n447), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n622), .B(new_n583), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n579), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n442), .A2(new_n500), .A3(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n323), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n313), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n356), .A2(new_n432), .ZN(new_n631));
  INV_X1    g0431(.A(new_n438), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n320), .A2(new_n322), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT92), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n320), .A2(KEYINPUT92), .A3(new_n322), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n392), .A2(new_n395), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n380), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n577), .A2(new_n575), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n578), .A2(new_n526), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(KEYINPUT26), .B2(new_n642), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n493), .A2(new_n494), .ZN(new_n645));
  INV_X1    g0445(.A(new_n457), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n493), .A2(KEYINPUT86), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n482), .A2(KEYINPUT86), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n645), .B(new_n617), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n526), .A2(new_n536), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n625), .A2(new_n652), .A3(new_n578), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n651), .A2(KEYINPUT91), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT91), .B1(new_n651), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n644), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n640), .B1(new_n657), .B2(new_n442), .ZN(G369));
  OR3_X1    g0458(.A1(new_n283), .A2(KEYINPUT27), .A3(G20), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT27), .B1(new_n283), .B2(G20), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n493), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n500), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n485), .A2(new_n493), .A3(new_n645), .A4(new_n663), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n603), .A2(new_n663), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n617), .A2(new_n671), .A3(new_n625), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT93), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  INV_X1    g0475(.A(new_n617), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n674), .A2(new_n675), .B1(new_n676), .B2(new_n663), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n663), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n485), .A2(new_n496), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n674), .A2(new_n682), .A3(new_n680), .A4(new_n675), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n220), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n558), .A2(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n228), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n627), .A2(new_n500), .A3(new_n663), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n509), .A2(new_n510), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n490), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT94), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n550), .A2(new_n612), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n695), .A2(KEYINPUT94), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(G179), .B1(new_n450), .B2(new_n455), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n610), .A3(new_n551), .A4(new_n693), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n698), .B1(new_n694), .B2(new_n697), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n663), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT31), .B(new_n663), .C1(new_n702), .C2(new_n703), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT95), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n706), .A2(KEYINPUT95), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n692), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n668), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n656), .A2(new_n680), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n653), .B1(new_n682), .B2(new_n676), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n663), .B1(new_n644), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n714), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n691), .B1(new_n721), .B2(G1), .ZN(G364));
  AND2_X1   g0522(.A1(new_n207), .A2(G13), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G45), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n687), .A2(G1), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(G330), .B1(new_n665), .B2(new_n666), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n669), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n725), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n665), .B2(new_n666), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n685), .A2(new_n254), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n734), .A2(G355), .B1(new_n462), .B2(new_n685), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n229), .A2(G45), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n246), .B2(G45), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n685), .A2(new_n274), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n735), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n224), .B1(G20), .B2(new_n366), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n731), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT96), .Z(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n207), .A2(new_n413), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n315), .A2(new_n310), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G326), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n254), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n746), .A2(new_n315), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n315), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n746), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n752), .A2(G303), .B1(new_n755), .B2(G322), .ZN(new_n756));
  INV_X1    g0556(.A(G311), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n207), .A2(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n753), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n747), .A2(new_n758), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  OAI221_X1 g0561(.A(new_n756), .B1(new_n757), .B2(new_n759), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n413), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n207), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n750), .B(new_n762), .C1(G294), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n758), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n767), .A2(G179), .A3(G200), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT97), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT97), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n767), .A2(G179), .A3(new_n310), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT99), .Z(new_n774));
  AOI22_X1  g0574(.A1(new_n772), .A2(G329), .B1(new_n774), .B2(G283), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n274), .B1(new_n751), .B2(new_n556), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT98), .ZN(new_n780));
  INV_X1    g0580(.A(new_n748), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G50), .A2(new_n781), .B1(new_n755), .B2(G58), .ZN(new_n782));
  INV_X1    g0582(.A(new_n760), .ZN(new_n783));
  INV_X1    g0583(.A(new_n759), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G68), .A2(new_n783), .B1(new_n784), .B2(G77), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n782), .B(new_n785), .C1(new_n459), .C2(new_n764), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n780), .B(new_n786), .C1(G107), .C2(new_n774), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n766), .A2(new_n775), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n741), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n745), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n728), .B1(new_n733), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n727), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  AOI211_X1 g0593(.A(new_n352), .B(new_n663), .C1(new_n354), .C2(new_n355), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n350), .A2(new_n663), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n339), .B2(new_n350), .ZN(new_n796));
  INV_X1    g0596(.A(new_n356), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n715), .B(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n728), .B1(new_n799), .B2(new_n714), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n714), .B2(new_n799), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n774), .A2(G87), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n757), .B2(new_n771), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT100), .Z(new_n804));
  AOI22_X1  g0604(.A1(G283), .A2(new_n783), .B1(new_n784), .B2(G116), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  INV_X1    g0606(.A(G303), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(new_n806), .B2(new_n754), .C1(new_n807), .C2(new_n748), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n254), .B1(new_n751), .B2(new_n326), .C1(new_n459), .C2(new_n764), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n781), .A2(G137), .B1(new_n784), .B2(G159), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT101), .B(G143), .Z(new_n812));
  OAI221_X1 g0612(.A(new_n811), .B1(new_n371), .B2(new_n760), .C1(new_n754), .C2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT34), .Z(new_n814));
  INV_X1    g0614(.A(new_n774), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n261), .ZN(new_n816));
  INV_X1    g0616(.A(G132), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n771), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G50), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n274), .B1(new_n751), .B2(new_n819), .C1(new_n260), .C2(new_n764), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n814), .A2(new_n816), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n741), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n741), .A2(new_n729), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n725), .B1(new_n211), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(new_n798), .C2(new_n730), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n801), .A2(new_n825), .ZN(G384));
  OAI211_X1 g0626(.A(G116), .B(new_n225), .C1(new_n520), .C2(KEYINPUT35), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(KEYINPUT35), .B2(new_n520), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT36), .ZN(new_n829));
  OR3_X1    g0629(.A1(new_n228), .A2(new_n211), .A3(new_n262), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n819), .A2(G68), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n206), .B(G13), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n434), .A2(new_n435), .ZN(new_n834));
  INV_X1    g0634(.A(new_n437), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(new_n835), .A3(new_n433), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n836), .A2(KEYINPUT102), .A3(new_n430), .A4(new_n663), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n430), .A2(new_n663), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n432), .A2(new_n438), .A3(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n430), .B(new_n663), .C1(new_n436), .C2(new_n437), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT102), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n837), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n656), .A2(new_n680), .A3(new_n798), .ZN(new_n845));
  INV_X1    g0645(.A(new_n794), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n259), .A2(KEYINPUT103), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n258), .A2(new_n267), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(KEYINPUT103), .B(new_n259), .C1(new_n276), .C2(new_n266), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n850), .A3(new_n282), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n851), .A2(KEYINPUT104), .A3(new_n290), .ZN(new_n852));
  INV_X1    g0652(.A(new_n661), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n318), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT104), .B1(new_n851), .B2(new_n290), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n292), .A2(new_n312), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT37), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n292), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n318), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n853), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n857), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n852), .A2(new_n855), .A3(new_n661), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n324), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n847), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n853), .B1(new_n636), .B2(new_n637), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT39), .B1(new_n870), .B2(new_n868), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n636), .A2(new_n630), .A3(new_n637), .ZN(new_n875));
  INV_X1    g0675(.A(new_n862), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n861), .A2(new_n862), .A3(new_n857), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n875), .A2(new_n876), .B1(new_n878), .B2(new_n864), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n869), .B(new_n874), .C1(new_n879), .C2(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n873), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n632), .A2(new_n680), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n872), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n871), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n442), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n717), .A2(new_n886), .A3(new_n720), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n640), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n885), .B(new_n888), .Z(new_n889));
  OAI21_X1  g0689(.A(new_n869), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n843), .A2(new_n798), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n495), .B(new_n491), .C1(new_n483), .C2(new_n484), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n579), .A2(new_n626), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(new_n499), .A4(new_n680), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n707), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n703), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n699), .A3(new_n701), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n898), .A2(KEYINPUT105), .A3(KEYINPUT31), .A4(new_n663), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n896), .A2(new_n899), .A3(new_n706), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n891), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n890), .B1(new_n901), .B2(KEYINPUT107), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n894), .A2(new_n900), .ZN(new_n903));
  INV_X1    g0703(.A(new_n891), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT40), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n870), .A2(new_n868), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n907), .A2(KEYINPUT40), .ZN(new_n908));
  AOI211_X1 g0708(.A(KEYINPUT106), .B(new_n891), .C1(new_n894), .C2(new_n900), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT106), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n903), .B2(new_n904), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n908), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n442), .B1(new_n894), .B2(new_n900), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n913), .B(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n915), .A2(new_n668), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n889), .A2(new_n916), .B1(new_n206), .B2(new_n723), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n889), .A2(new_n916), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n833), .B1(new_n917), .B2(new_n918), .ZN(G367));
  NAND2_X1  g0719(.A1(new_n532), .A2(new_n663), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n652), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n526), .A2(new_n663), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT110), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n683), .B2(new_n681), .ZN(new_n926));
  OR3_X1    g0726(.A1(new_n926), .A2(KEYINPUT42), .A3(new_n683), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT42), .B1(new_n926), .B2(new_n683), .ZN(new_n928));
  INV_X1    g0728(.A(new_n925), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n539), .B1(new_n929), .B2(new_n617), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n680), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n570), .A2(new_n663), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n641), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n578), .B2(new_n933), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT108), .ZN(new_n936));
  XNOR2_X1  g0736(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(KEYINPUT43), .B2(new_n936), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n679), .A2(new_n929), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n927), .A2(new_n928), .A3(new_n931), .A4(new_n938), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n941), .B1(new_n940), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n686), .B(KEYINPUT41), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n926), .A2(KEYINPUT44), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT44), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n948), .B(new_n925), .C1(new_n683), .C2(new_n681), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n683), .A2(new_n925), .A3(new_n681), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT45), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n947), .A2(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n678), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n950), .B(new_n951), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n679), .B(new_n956), .C1(new_n947), .C2(new_n949), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n677), .B1(new_n892), .B2(new_n663), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n683), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(new_n669), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n955), .A2(new_n957), .A3(new_n721), .A4(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n946), .B1(new_n961), .B2(new_n721), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n724), .A2(G1), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n945), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n744), .B1(new_n220), .B2(new_n573), .C1(new_n239), .C2(new_n739), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT111), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n967), .A2(new_n728), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n772), .A2(G137), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n764), .A2(new_n261), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n754), .A2(new_n371), .B1(new_n759), .B2(new_n819), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n254), .B(new_n973), .C1(G77), .C2(new_n773), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n751), .A2(new_n260), .B1(new_n760), .B2(new_n776), .ZN(new_n975));
  INV_X1    g0775(.A(new_n812), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n975), .B1(new_n781), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n970), .A2(new_n972), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n751), .A2(new_n462), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n979), .A2(KEYINPUT46), .B1(new_n326), .B2(new_n764), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(KEYINPUT46), .B2(new_n979), .ZN(new_n981));
  INV_X1    g0781(.A(G283), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n760), .A2(new_n806), .B1(new_n759), .B2(new_n982), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n274), .B(new_n983), .C1(G97), .C2(new_n773), .ZN(new_n984));
  INV_X1    g0784(.A(G317), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n981), .B(new_n984), .C1(new_n985), .C2(new_n771), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n748), .A2(new_n757), .B1(new_n754), .B2(new_n807), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT112), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n978), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT47), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n741), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n969), .B1(new_n991), .B2(new_n992), .C1(new_n936), .C2(new_n732), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n964), .A2(new_n993), .ZN(G387));
  OAI22_X1  g0794(.A1(new_n748), .A2(new_n776), .B1(new_n754), .B2(new_n819), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n573), .A2(new_n764), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n760), .A2(new_n286), .B1(new_n759), .B2(new_n261), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n274), .B1(new_n751), .B2(new_n211), .ZN(new_n998));
  NOR4_X1   g0798(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n371), .B2(new_n771), .C1(new_n815), .C2(new_n459), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n765), .A2(G283), .B1(new_n752), .B2(G294), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n781), .A2(G322), .B1(new_n784), .B2(G303), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n757), .B2(new_n760), .C1(new_n985), .C2(new_n754), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n274), .B1(new_n773), .B2(G116), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1007), .B(new_n1008), .C1(new_n749), .C2(new_n771), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n741), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n688), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1013), .A2(new_n734), .B1(new_n326), .B2(new_n685), .ZN(new_n1014));
  INV_X1    g0814(.A(G45), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n234), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n286), .A2(G50), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT50), .ZN(new_n1018));
  AOI21_X1  g0818(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n1013), .C2(KEYINPUT113), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1013), .A2(KEYINPUT113), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n738), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1014), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n725), .B1(new_n1023), .B2(new_n744), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1012), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT114), .Z(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n677), .B2(new_n731), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n960), .B2(new_n963), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n960), .A2(new_n721), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n686), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n960), .A2(new_n721), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(G393));
  AOI21_X1  g0832(.A(new_n743), .B1(G97), .B2(new_n685), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n738), .A2(new_n243), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n725), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n772), .A2(G322), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n774), .A2(G107), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n752), .A2(G283), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n274), .B1(new_n784), .B2(G294), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n764), .A2(new_n462), .B1(new_n760), .B2(new_n807), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT116), .Z(new_n1042));
  OAI22_X1  g0842(.A1(new_n748), .A2(new_n985), .B1(new_n754), .B2(new_n757), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n748), .A2(new_n371), .B1(new_n754), .B2(new_n776), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT51), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n802), .B(new_n1047), .C1(new_n771), .C2(new_n812), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n751), .A2(new_n261), .B1(new_n760), .B2(new_n819), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n764), .A2(new_n211), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n274), .B1(new_n759), .B2(new_n286), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1040), .A2(new_n1045), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1035), .B1(new_n789), .B2(new_n1054), .C1(new_n925), .C2(new_n732), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT115), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n947), .A2(new_n949), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n679), .B1(new_n1058), .B2(new_n956), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n954), .A2(new_n678), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n955), .A2(new_n957), .A3(KEYINPUT115), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1056), .B1(new_n1063), .B2(new_n963), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1029), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(new_n686), .A3(new_n961), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(KEYINPUT117), .A3(new_n1066), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n955), .A2(new_n957), .A3(KEYINPUT115), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT115), .B1(new_n955), .B2(new_n957), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n963), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n1066), .A3(new_n1055), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT117), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1067), .A2(new_n1073), .ZN(G390));
  AOI21_X1  g0874(.A(new_n816), .B1(G294), .B2(new_n772), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n781), .A2(G283), .B1(new_n784), .B2(G97), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G107), .A2(new_n783), .B1(new_n755), .B2(G116), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n274), .B(new_n1050), .C1(G87), .C2(new_n752), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n254), .B1(new_n773), .B2(G50), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n776), .B2(new_n764), .ZN(new_n1081));
  INV_X1    g0881(.A(G128), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n748), .A2(new_n1082), .B1(new_n754), .B2(new_n817), .ZN(new_n1083));
  INV_X1    g0883(.A(G137), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT54), .B(G143), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n760), .A2(new_n1084), .B1(new_n759), .B2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1081), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n751), .A2(new_n371), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT53), .ZN(new_n1089));
  INV_X1    g0889(.A(G125), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1087), .B(new_n1089), .C1(new_n1090), .C2(new_n771), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n789), .B1(new_n1079), .B2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n725), .B(new_n1092), .C1(new_n286), .C2(new_n823), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n881), .B2(new_n730), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n873), .B(new_n880), .C1(new_n847), .C2(new_n883), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n796), .A2(new_n797), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n794), .B1(new_n719), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n882), .B(new_n890), .C1(new_n1097), .C2(new_n844), .ZN(new_n1098));
  OAI211_X1 g0898(.A(G330), .B(new_n904), .C1(new_n692), .C2(new_n712), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1095), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n845), .A2(new_n846), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n883), .B1(new_n1101), .B2(new_n843), .ZN(new_n1102));
  OAI211_X1 g0902(.A(KEYINPUT118), .B(new_n1098), .C1(new_n1102), .C2(new_n881), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n798), .A2(G330), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n903), .A2(new_n843), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT118), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1100), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n963), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1094), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(G330), .B(new_n798), .C1(new_n692), .C2(new_n712), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n844), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1106), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n903), .A2(new_n1105), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n844), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1115), .A2(new_n1101), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n914), .A2(G330), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n887), .A2(new_n640), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1100), .B(new_n1122), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1122), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n687), .B1(new_n1110), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1112), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(G378));
  INV_X1    g0927(.A(new_n885), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n661), .B1(new_n381), .B2(new_n383), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n396), .A2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1129), .B(new_n380), .C1(new_n392), .C2(new_n395), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1133));
  NOR3_X1   g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1133), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n380), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n395), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n394), .B1(new_n393), .B2(new_n387), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n1129), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n396), .A2(new_n1130), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1135), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1134), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n913), .B2(G330), .ZN(new_n1144));
  OAI21_X1  g0944(.A(KEYINPUT120), .B1(new_n1134), .B2(new_n1142), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1133), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1140), .A2(new_n1141), .A3(new_n1135), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT120), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n668), .B(new_n1150), .C1(new_n906), .C2(new_n912), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1128), .B1(new_n1144), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1150), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n913), .A2(G330), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n668), .B1(new_n906), .B2(new_n912), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n885), .C1(new_n1155), .C2(new_n1143), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1121), .ZN(new_n1157));
  AOI221_X4 g0957(.A(KEYINPUT57), .B1(new_n1152), .B2(new_n1156), .C1(new_n1123), .C2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1123), .A2(new_n1157), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n686), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n823), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n728), .B1(G50), .B2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT119), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1150), .A2(new_n730), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n748), .A2(new_n1090), .B1(new_n760), .B2(new_n817), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1085), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n752), .A2(new_n1169), .B1(new_n755), .B2(G128), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1084), .B2(new_n759), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1168), .B(new_n1171), .C1(G150), .C2(new_n765), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n772), .A2(G124), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G33), .B(G41), .C1(new_n773), .C2(G159), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n274), .A2(G41), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G97), .A2(new_n783), .B1(new_n755), .B2(G107), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n771), .C2(new_n982), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n773), .A2(G58), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n211), .B2(new_n751), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n573), .A2(new_n759), .B1(new_n462), .B2(new_n748), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1181), .A2(new_n971), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1179), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n819), .C1(G33), .C2(G41), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1178), .A2(new_n1186), .A3(new_n1187), .A4(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1166), .B(new_n1167), .C1(new_n741), .C2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1161), .B2(new_n963), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1163), .A2(new_n1192), .ZN(G375));
  OAI21_X1  g0993(.A(new_n728), .B1(G68), .B2(new_n1164), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n752), .A2(G159), .B1(new_n783), .B2(new_n1169), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1084), .B2(new_n754), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n772), .B2(G128), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n764), .A2(new_n819), .B1(new_n759), .B2(new_n371), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT123), .Z(new_n1199));
  NAND3_X1  g0999(.A1(new_n781), .A2(KEYINPUT122), .A3(G132), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT122), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n748), .B2(new_n817), .ZN(new_n1202));
  AND4_X1   g1002(.A1(new_n274), .A2(new_n1182), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1197), .A2(new_n1199), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n274), .B1(new_n774), .B2(G77), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT121), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n772), .A2(G303), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n996), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n751), .A2(new_n459), .B1(new_n760), .B2(new_n462), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G294), .B2(new_n781), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G283), .A2(new_n755), .B1(new_n784), .B2(G107), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1204), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1194), .B1(new_n1213), .B2(new_n741), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n843), .B2(new_n730), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1119), .B2(new_n1111), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1122), .A2(new_n946), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1115), .A2(new_n1101), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(new_n1157), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1217), .B1(new_n1218), .B2(new_n1222), .ZN(G381));
  NAND4_X1  g1023(.A1(new_n1067), .A2(new_n1073), .A3(new_n964), .A4(new_n993), .ZN(new_n1224));
  OR2_X1    g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1224), .A2(G384), .A3(G381), .A4(new_n1225), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT124), .Z(new_n1227));
  NAND3_X1  g1027(.A1(new_n1163), .A2(new_n1126), .A3(new_n1192), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1227), .A2(new_n1228), .ZN(G407));
  NAND2_X1  g1029(.A1(new_n662), .A2(G213), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(G213), .B(new_n1231), .C1(new_n1227), .C2(new_n1228), .ZN(G409));
  XNOR2_X1  g1032(.A(G393), .B(new_n792), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT117), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1234));
  AND4_X1   g1034(.A1(KEYINPUT117), .A2(new_n1070), .A3(new_n1066), .A4(new_n1055), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1234), .A2(G387), .A3(new_n1235), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1067), .A2(new_n1073), .B1(new_n964), .B2(new_n993), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1233), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G390), .A2(G387), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1233), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1224), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1238), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1230), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n686), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT60), .B1(new_n1221), .B2(new_n1157), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1119), .A2(new_n1121), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1245), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(new_n1216), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(G384), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n801), .B(new_n825), .C1(new_n1249), .C2(new_n1216), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1163), .A2(G378), .A3(new_n1192), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1192), .B1(new_n1255), .B2(new_n946), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1126), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1244), .B(new_n1253), .C1(new_n1254), .C2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1243), .B1(new_n1258), .B2(KEYINPUT63), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1244), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT126), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1244), .A2(KEYINPUT125), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1251), .A2(new_n1252), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1244), .A2(G2897), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1264), .B(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1261), .A2(new_n1262), .A3(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT126), .B1(new_n1260), .B2(new_n1267), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1253), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1230), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1259), .A2(new_n1269), .A3(new_n1270), .A4(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1273), .A2(KEYINPUT62), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1242), .B1(new_n1260), .B2(new_n1267), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1260), .B2(new_n1272), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1276), .B1(new_n1281), .B2(new_n1282), .ZN(G405));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1254), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1238), .A2(new_n1241), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(new_n1284), .A3(new_n1254), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G378), .B1(new_n1163), .B2(new_n1192), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1272), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1289), .B(new_n1291), .ZN(G402));
endmodule


