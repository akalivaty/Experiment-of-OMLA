//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(new_n203), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n210), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n213), .B1(new_n217), .B2(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  AND2_X1   g0045(.A1(new_n245), .A2(new_n214), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n204), .A2(G20), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n249), .A2(new_n251), .B1(G150), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n246), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n245), .A2(new_n214), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G20), .ZN(new_n261));
  OAI21_X1  g0061(.A(G50), .B1(new_n261), .B2(G1), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n260), .A2(new_n262), .B1(G50), .B2(new_n256), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT9), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n271), .A3(G274), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n250), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G223), .A3(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G77), .ZN(new_n283));
  INV_X1    g0083(.A(G222), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G1698), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n286), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n282), .B1(new_n283), .B2(new_n281), .C1(new_n284), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n271), .ZN(new_n293));
  AOI211_X1 g0093(.A(new_n273), .B(new_n277), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G190), .ZN(new_n295));
  INV_X1    g0095(.A(G200), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n266), .B(new_n295), .C1(new_n296), .C2(new_n294), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT10), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT68), .B(G179), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n300), .B(KEYINPUT69), .Z(new_n301));
  INV_X1    g0101(.A(new_n264), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n301), .B(new_n302), .C1(G169), .C2(new_n294), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n249), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT15), .B(G87), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(KEYINPUT70), .A3(new_n251), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT70), .B1(new_n306), .B2(new_n251), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n258), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n283), .B1(new_n255), .B2(G20), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n259), .A2(new_n311), .B1(new_n283), .B2(new_n257), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G238), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n286), .A2(new_n288), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n281), .B1(new_n315), .B2(new_n285), .C1(new_n316), .C2(new_n230), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n293), .C1(G107), .C2(new_n281), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n273), .B1(G244), .B2(new_n276), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G200), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n314), .B(new_n321), .C1(new_n322), .C2(new_n320), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n318), .A2(new_n299), .A3(new_n319), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n325), .A2(new_n313), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n298), .A2(new_n303), .A3(new_n323), .A4(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT12), .B1(new_n256), .B2(G68), .ZN(new_n330));
  OR3_X1    g0130(.A1(new_n256), .A2(KEYINPUT12), .A3(G68), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n203), .B1(new_n255), .B2(G20), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n330), .A2(new_n331), .B1(new_n259), .B2(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n334));
  INV_X1    g0134(.A(new_n251), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(new_n283), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n336), .A2(new_n258), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(KEYINPUT11), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n271), .A2(G238), .A3(new_n274), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n272), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n272), .A2(new_n341), .A3(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n289), .A2(new_n290), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n286), .A2(new_n288), .A3(G226), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G232), .A2(G1698), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT71), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n293), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n346), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT13), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n346), .A2(new_n359), .A3(new_n356), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n340), .B1(new_n361), .B2(G200), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT73), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n359), .B1(new_n346), .B2(new_n356), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT73), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n364), .A2(new_n366), .A3(G190), .A4(new_n360), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n340), .B(KEYINPUT74), .ZN(new_n369));
  INV_X1    g0169(.A(new_n360), .ZN(new_n370));
  OAI21_X1  g0170(.A(G169), .B1(new_n370), .B2(new_n365), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n364), .A2(new_n366), .A3(G179), .A4(new_n360), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n361), .A2(new_n374), .A3(G169), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n368), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n377), .A2(KEYINPUT75), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(KEYINPUT75), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n329), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n272), .B1(new_n230), .B2(new_n275), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT79), .B(G190), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  AND2_X1   g0184(.A1(KEYINPUT76), .A2(G33), .ZN(new_n385));
  NOR2_X1   g0185(.A1(KEYINPUT76), .A2(G33), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT3), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n279), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n286), .A2(new_n288), .A3(G223), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G226), .A2(G1698), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n388), .A2(new_n391), .B1(G33), .B2(G87), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n382), .B(new_n384), .C1(new_n392), .C2(new_n271), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT67), .B(G1698), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT76), .B(G33), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n290), .B1(new_n396), .B2(KEYINPUT3), .ZN(new_n397));
  INV_X1    g0197(.A(G87), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n395), .A2(new_n397), .B1(new_n250), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n381), .B1(new_n399), .B2(new_n293), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n393), .B1(new_n400), .B2(G200), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G58), .A2(G68), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT77), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(KEYINPUT77), .A2(G58), .A3(G68), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n218), .A3(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(G20), .B1(G159), .B2(new_n252), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n397), .B2(new_n261), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n387), .A2(new_n408), .A3(new_n261), .A4(new_n279), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G68), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT16), .B(new_n407), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n289), .A2(new_n408), .A3(G20), .ZN(new_n414));
  OR2_X1    g0214(.A1(KEYINPUT76), .A2(G33), .ZN(new_n415));
  NAND2_X1  g0215(.A1(KEYINPUT76), .A2(G33), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n278), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n279), .A2(new_n261), .A3(new_n280), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n408), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n203), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n407), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n413), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n412), .A2(new_n423), .A3(new_n258), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n248), .B1(new_n255), .B2(G20), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n259), .B1(new_n257), .B2(new_n248), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n401), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n401), .A2(new_n424), .A3(KEYINPUT17), .A4(new_n426), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT80), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(KEYINPUT80), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n424), .A2(new_n426), .ZN(new_n435));
  INV_X1    g0235(.A(new_n299), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n382), .B(new_n436), .C1(new_n392), .C2(new_n271), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n400), .B2(new_n324), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n435), .A2(KEYINPUT18), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT18), .B1(new_n435), .B2(new_n438), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT78), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n435), .A2(new_n438), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT78), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n433), .A2(new_n434), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n380), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT86), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n286), .A2(new_n288), .A3(G250), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G257), .A2(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n388), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G294), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n415), .B2(new_n416), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n449), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  AOI211_X1 g0257(.A(KEYINPUT86), .B(new_n455), .C1(new_n388), .C2(new_n452), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n293), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n255), .A2(G45), .ZN(new_n460));
  OR2_X1    g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G274), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n215), .B2(new_n270), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g0266(.A(KEYINPUT5), .B(G41), .ZN(new_n467));
  INV_X1    g0267(.A(new_n460), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n467), .A2(new_n468), .B1(new_n215), .B2(new_n270), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G264), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n459), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G200), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n459), .A2(G190), .A3(new_n466), .A4(new_n470), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT25), .B1(new_n257), .B2(new_n207), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n255), .A2(G33), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n246), .A2(new_n256), .A3(new_n476), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n474), .A2(new_n475), .B1(new_n477), .B2(new_n207), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n415), .B2(new_n416), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n261), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n261), .A2(G87), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n347), .B2(new_n485), .ZN(new_n486));
  OR3_X1    g0286(.A1(new_n261), .A2(KEYINPUT23), .A3(G107), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT23), .B1(new_n261), .B2(G107), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n483), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT22), .A2(G87), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n397), .A2(G20), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n480), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(new_n488), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n261), .B2(new_n482), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n388), .A2(KEYINPUT22), .A3(new_n261), .A4(G87), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(new_n495), .A3(new_n479), .A4(new_n486), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n478), .B1(new_n497), .B2(new_n258), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n472), .A2(new_n473), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n459), .A2(G179), .A3(new_n466), .A4(new_n470), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n279), .A2(new_n387), .B1(new_n450), .B2(new_n451), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT86), .B1(new_n501), .B2(new_n455), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n453), .A2(new_n449), .A3(new_n456), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n271), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n466), .ZN(new_n505));
  INV_X1    g0305(.A(new_n470), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n500), .B1(new_n507), .B2(new_n324), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n498), .B1(new_n508), .B2(KEYINPUT87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n471), .A2(G169), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT87), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n500), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n499), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  OAI211_X1 g0315(.A(G250), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n516));
  NAND2_X1  g0316(.A1(KEYINPUT4), .A2(G244), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n515), .B(new_n516), .C1(new_n291), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n394), .A2(G244), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n397), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT82), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n286), .A2(new_n288), .A3(G244), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT4), .B1(new_n388), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n525), .A2(new_n518), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n293), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n469), .A2(G257), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n466), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(G190), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n519), .A2(new_n522), .A3(KEYINPUT82), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n526), .B1(new_n525), .B2(new_n518), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n271), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(G200), .B1(new_n535), .B2(new_n530), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n257), .A2(new_n206), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n477), .B2(new_n206), .ZN(new_n538));
  XOR2_X1   g0338(.A(KEYINPUT81), .B(KEYINPUT6), .Z(new_n539));
  NAND2_X1  g0339(.A1(new_n207), .A2(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n208), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(G20), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n252), .A2(G77), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n417), .A2(new_n414), .B1(new_n419), .B2(new_n408), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n545), .B(new_n546), .C1(new_n207), .C2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n538), .B1(new_n548), .B2(new_n258), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n532), .A2(new_n536), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n530), .A2(new_n436), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n549), .B1(new_n528), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n324), .B1(new_n535), .B2(new_n530), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n353), .B2(new_n354), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n557), .A2(G20), .B1(G87), .B2(new_n208), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n278), .B1(new_n415), .B2(new_n416), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n261), .B(G68), .C1(new_n559), .C2(new_n290), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n556), .B1(new_n335), .B2(new_n206), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n258), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n305), .A2(new_n257), .ZN(new_n564));
  AND4_X1   g0364(.A1(new_n214), .A2(new_n256), .A3(new_n245), .A4(new_n476), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n306), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n460), .A2(G250), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n465), .A2(new_n468), .B1(new_n568), .B2(new_n271), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G244), .A2(G1698), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n316), .B2(new_n315), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n482), .B1(new_n571), .B2(new_n388), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n569), .B1(new_n572), .B2(new_n271), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n324), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n299), .B(new_n569), .C1(new_n572), .C2(new_n271), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n567), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(G200), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n562), .A2(new_n258), .B1(new_n257), .B2(new_n305), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n565), .A2(G87), .ZN(new_n579));
  OAI211_X1 g0379(.A(G190), .B(new_n569), .C1(new_n572), .C2(new_n271), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n469), .A2(G270), .B1(new_n465), .B2(new_n463), .ZN(new_n583));
  INV_X1    g0383(.A(G303), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n281), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n286), .A2(new_n288), .A3(G257), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G264), .A2(G1698), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n388), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n583), .B(new_n383), .C1(new_n589), .C2(new_n271), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n256), .A2(G116), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n477), .B2(new_n481), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n515), .B(new_n261), .C1(G33), .C2(new_n206), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n481), .A2(G20), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n258), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n594), .A2(KEYINPUT20), .A3(new_n258), .A4(new_n595), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n593), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n279), .A2(new_n387), .B1(new_n586), .B2(new_n587), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n293), .B1(new_n602), .B2(new_n585), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n296), .B1(new_n603), .B2(new_n583), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT83), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n583), .B1(new_n589), .B2(new_n271), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT83), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n600), .A4(new_n590), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n598), .A2(new_n599), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n591), .B1(new_n565), .B2(G116), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n324), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n606), .A3(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n612), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n615), .A2(G179), .A3(new_n603), .A4(new_n583), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT21), .B1(new_n613), .B2(new_n606), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT84), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n610), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n620), .B1(new_n610), .B2(new_n619), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n555), .B(new_n582), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n448), .A2(new_n514), .A3(new_n624), .ZN(G372));
  INV_X1    g0425(.A(new_n303), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n439), .A2(new_n440), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n433), .A2(new_n434), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n362), .A2(new_n367), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n376), .A2(new_n369), .B1(new_n631), .B2(new_n327), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n628), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n626), .B1(new_n633), .B2(new_n298), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n498), .B1(new_n510), .B2(new_n500), .ZN(new_n635));
  INV_X1    g0435(.A(new_n619), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT88), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n497), .A2(new_n258), .ZN(new_n639));
  INV_X1    g0439(.A(new_n478), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n502), .A2(new_n503), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n506), .B1(new_n642), .B2(new_n293), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n324), .B1(new_n643), .B2(new_n466), .ZN(new_n644));
  INV_X1    g0444(.A(G179), .ZN(new_n645));
  NOR4_X1   g0445(.A1(new_n504), .A2(new_n645), .A3(new_n505), .A4(new_n506), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n641), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT88), .B1(new_n647), .B2(new_n619), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n472), .A2(new_n473), .A3(new_n498), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n550), .A3(new_n582), .A4(new_n554), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n638), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n552), .A2(new_n553), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT26), .B1(new_n652), .B2(new_n582), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n576), .A2(new_n581), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n554), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n576), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n634), .B1(new_n448), .B2(new_n658), .ZN(G369));
  INV_X1    g0459(.A(G330), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n610), .A2(new_n619), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT84), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n621), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n255), .A2(new_n261), .A3(G13), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT27), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G213), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n615), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n619), .A2(new_n670), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n660), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT87), .B1(new_n644), .B2(new_n646), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n512), .A3(new_n641), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n641), .A2(KEYINPUT89), .A3(new_n669), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  INV_X1    g0477(.A(new_n669), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n498), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n675), .A2(new_n680), .A3(new_n649), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n509), .A2(new_n512), .A3(new_n669), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n635), .A2(new_n678), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n619), .A2(new_n669), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n513), .A2(new_n680), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(G399));
  NAND2_X1  g0488(.A1(new_n211), .A2(new_n267), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n255), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n692));
  INV_X1    g0492(.A(new_n219), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n691), .A2(new_n692), .B1(new_n693), .B2(new_n690), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  OAI21_X1  g0495(.A(new_n678), .B1(new_n651), .B2(new_n657), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n650), .B1(new_n675), .B2(new_n619), .ZN(new_n699));
  OAI211_X1 g0499(.A(KEYINPUT29), .B(new_n678), .C1(new_n699), .C2(new_n657), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n583), .B(G179), .C1(new_n589), .C2(new_n271), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n573), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n643), .A2(new_n528), .A3(new_n702), .A4(new_n531), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n535), .A2(new_n530), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n643), .A4(new_n702), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n528), .A2(new_n531), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n606), .A2(new_n573), .A3(new_n299), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n471), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n678), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT90), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT90), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(new_n717), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n550), .A2(new_n554), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n654), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n513), .A2(new_n663), .A3(new_n721), .A4(new_n678), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n712), .A2(new_n669), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT91), .A3(new_n713), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT91), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n709), .B1(new_n643), .B2(new_n466), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n704), .A2(new_n703), .B1(new_n726), .B2(new_n708), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n678), .B1(new_n727), .B2(new_n707), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n725), .B1(new_n728), .B2(KEYINPUT31), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n719), .A2(new_n722), .A3(new_n724), .A4(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n698), .A2(new_n700), .B1(G330), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n695), .B1(new_n731), .B2(G1), .ZN(G364));
  INV_X1    g0532(.A(new_n673), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n671), .A2(new_n660), .A3(new_n672), .ZN(new_n734));
  INV_X1    g0534(.A(G13), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G45), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(KEYINPUT92), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n691), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n733), .A2(new_n734), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n742), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n281), .A2(new_n211), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n746), .B1(G116), .B2(new_n211), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n240), .A2(G45), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n397), .A2(new_n211), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n268), .B2(new_n693), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n214), .B1(G20), .B2(new_n324), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n744), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n261), .A2(G179), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(new_n322), .A3(new_n296), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G159), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n322), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n261), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n762), .A2(KEYINPUT32), .B1(G97), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n759), .A2(new_n322), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n207), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n347), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n766), .B(new_n769), .C1(KEYINPUT32), .C2(new_n762), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT96), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT96), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n398), .ZN(new_n776));
  OR3_X1    g0576(.A1(new_n299), .A2(KEYINPUT93), .A3(new_n261), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT93), .B1(new_n299), .B2(new_n261), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n296), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n384), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n770), .B(new_n776), .C1(G58), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n296), .B1(new_n777), .B2(new_n778), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT94), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(KEYINPUT94), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n784), .A2(new_n322), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n780), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n782), .B1(new_n203), .B2(new_n786), .C1(new_n283), .C2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n784), .A2(new_n383), .A3(new_n785), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT95), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n784), .A2(KEYINPUT95), .A3(new_n383), .A4(new_n785), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G50), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n281), .B1(new_n761), .B2(G329), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n797), .B1(new_n798), .B2(new_n767), .C1(new_n454), .C2(new_n764), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n775), .A2(new_n584), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(G311), .C2(new_n787), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  INV_X1    g0602(.A(new_n781), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n804));
  INV_X1    g0604(.A(G317), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n801), .B1(new_n802), .B2(new_n803), .C1(new_n786), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n792), .A2(new_n793), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n808), .A2(G326), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n789), .A2(new_n796), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n758), .B1(new_n810), .B2(new_n755), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n671), .A2(new_n672), .A3(new_n754), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n743), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NOR2_X1   g0615(.A1(new_n755), .A2(new_n752), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n742), .B1(new_n283), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n327), .A2(new_n678), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n313), .A2(new_n669), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n323), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n818), .B1(new_n820), .B2(new_n327), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n786), .A2(new_n798), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n767), .A2(new_n398), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n347), .B1(new_n760), .B2(new_n825), .C1(new_n764), .C2(new_n206), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n824), .B(new_n826), .C1(new_n774), .C2(G107), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n827), .B1(new_n803), .B2(new_n454), .C1(new_n481), .C2(new_n788), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n823), .B(new_n828), .C1(G303), .C2(new_n808), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n787), .A2(G159), .B1(new_n781), .B2(G143), .ZN(new_n830));
  INV_X1    g0630(.A(G150), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n786), .C1(new_n794), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT34), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n388), .B1(new_n835), .B2(new_n760), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n764), .A2(new_n202), .B1(new_n767), .B2(new_n203), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(new_n774), .C2(G50), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n829), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n755), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n817), .B1(new_n822), .B2(new_n753), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n696), .A2(new_n821), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(KEYINPUT98), .ZN(new_n844));
  INV_X1    g0644(.A(new_n650), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n647), .A2(KEYINPUT88), .A3(new_n619), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n637), .B1(new_n635), .B2(new_n636), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n576), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n652), .A2(KEYINPUT26), .A3(new_n582), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n655), .B1(new_n554), .B2(new_n654), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n669), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(new_n822), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n844), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n730), .A2(G330), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n744), .B1(new_n855), .B2(new_n856), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n842), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  NOR2_X1   g0660(.A1(new_n736), .A2(new_n255), .ZN(new_n861));
  INV_X1    g0661(.A(new_n667), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n628), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n818), .B1(new_n696), .B2(new_n821), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n376), .A2(new_n369), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n369), .A2(new_n669), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n631), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n369), .B(new_n669), .C1(new_n368), .C2(new_n376), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n409), .A2(new_n411), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT16), .B1(new_n874), .B2(new_n407), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n412), .A2(new_n258), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n426), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n862), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n441), .A2(new_n446), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n878), .B1(new_n629), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n438), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n878), .A3(new_n427), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n435), .A2(new_n862), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n442), .A2(new_n884), .A3(new_n885), .A4(new_n427), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n873), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n886), .ZN(new_n889));
  OAI211_X1 g0689(.A(KEYINPUT38), .B(new_n889), .C1(new_n447), .C2(new_n878), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n863), .B1(new_n872), .B2(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n435), .B(new_n862), .C1(new_n627), .C2(new_n431), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n442), .A2(new_n884), .A3(new_n427), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n886), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n894), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n890), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n888), .B2(new_n890), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT101), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n435), .A2(KEYINPUT18), .A3(new_n438), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n445), .B1(new_n444), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n440), .A2(KEYINPUT78), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n429), .A2(KEYINPUT80), .A3(new_n430), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT80), .B1(new_n429), .B2(new_n430), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n906), .A2(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n878), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n912), .B2(new_n889), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n880), .A2(new_n887), .A3(new_n873), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT39), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT101), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n890), .A2(new_n900), .A3(new_n901), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n866), .A2(new_n669), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n904), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n892), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n700), .B1(new_n853), .B2(KEYINPUT29), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n634), .B1(new_n448), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n723), .A2(new_n713), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n675), .A2(new_n649), .A3(new_n678), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n925), .B(new_n715), .C1(new_n624), .C2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n821), .B1(new_n868), .B2(new_n869), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n890), .A2(new_n900), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT102), .A4(KEYINPUT40), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT102), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n910), .A2(new_n911), .B1(new_n886), .B2(new_n883), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n899), .B1(new_n933), .B2(KEYINPUT38), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n927), .A2(KEYINPUT40), .A3(new_n928), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n891), .A2(new_n929), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n931), .A2(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n723), .A2(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n448), .B1(new_n722), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n660), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n939), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n861), .B1(new_n924), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n924), .B2(new_n943), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n693), .A2(G77), .A3(new_n404), .A4(new_n405), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n201), .A2(G68), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(G1), .A3(new_n735), .ZN(new_n949));
  INV_X1    g0749(.A(new_n217), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT35), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n541), .A2(new_n544), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n950), .B(G116), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n945), .A2(new_n949), .A3(new_n956), .ZN(G367));
  OAI221_X1 g0757(.A(new_n756), .B1(new_n211), .B2(new_n305), .C1(new_n236), .C2(new_n749), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n744), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n754), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n578), .A2(new_n579), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n669), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n582), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(KEYINPUT103), .C1(new_n576), .C2(new_n962), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n962), .A2(new_n576), .A3(KEYINPUT103), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n774), .A2(G116), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n454), .B2(new_n786), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT108), .Z(new_n970));
  NOR2_X1   g0770(.A1(new_n767), .A2(new_n206), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n397), .B1(new_n805), .B2(new_n760), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(G107), .C2(new_n765), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n803), .B2(new_n584), .C1(new_n798), .C2(new_n788), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G311), .B2(new_n808), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n764), .A2(new_n203), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n281), .B1(new_n760), .B2(new_n832), .C1(new_n283), .C2(new_n767), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(new_n774), .C2(G58), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n803), .B2(new_n831), .C1(new_n201), .C2(new_n788), .ZN(new_n979));
  INV_X1    g0779(.A(new_n786), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(G159), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n808), .A2(G143), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n970), .A2(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n983), .A2(KEYINPUT47), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n755), .B1(new_n983), .B2(KEYINPUT47), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n959), .B1(new_n960), .B2(new_n966), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n740), .A2(new_n255), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n686), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n681), .A2(new_n682), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n673), .A2(new_n687), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n856), .A2(new_n922), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT106), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n990), .A2(new_n993), .A3(new_n687), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n993), .B1(new_n990), .B2(new_n687), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n995), .A2(new_n996), .A3(new_n673), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT107), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT107), .ZN(new_n999));
  INV_X1    g0799(.A(new_n996), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(new_n994), .A3(new_n733), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n731), .A2(new_n999), .A3(new_n1001), .A4(new_n991), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n684), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n687), .A2(new_n685), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT104), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n652), .A2(new_n1006), .A3(new_n669), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT104), .B1(new_n554), .B2(new_n678), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n549), .A2(new_n678), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1007), .A2(new_n1008), .B1(new_n555), .B2(new_n1010), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1005), .A2(KEYINPUT44), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT44), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n555), .A2(new_n1010), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n687), .A2(new_n1017), .A3(new_n685), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n687), .A2(new_n1017), .A3(KEYINPUT45), .A4(new_n685), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1004), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n684), .C1(new_n1013), .C2(new_n1012), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n731), .B1(new_n1003), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n689), .B(KEYINPUT41), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n988), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n684), .A2(new_n1011), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n554), .B1(new_n1011), .B2(new_n675), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n678), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT42), .B1(new_n687), .B2(new_n1011), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(KEYINPUT105), .A3(new_n1038), .ZN(new_n1039));
  OR3_X1    g0839(.A1(new_n687), .A2(new_n1011), .A3(KEYINPUT42), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT105), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1034), .B(new_n1035), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NOR4_X1   g0844(.A1(new_n1041), .A2(new_n1042), .A3(KEYINPUT43), .A4(new_n966), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1032), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1035), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n1033), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n1031), .A3(new_n1043), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n986), .B1(new_n1030), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT109), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(KEYINPUT109), .B(new_n986), .C1(new_n1030), .C2(new_n1050), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(G387));
  INV_X1    g0855(.A(new_n971), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n774), .A2(G77), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n397), .B1(G150), .B2(new_n761), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n765), .A2(new_n306), .ZN(new_n1059));
  AND4_X1   g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n803), .B2(new_n795), .C1(new_n203), .C2(new_n788), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n249), .B2(new_n980), .ZN(new_n1062));
  INV_X1    g0862(.A(G159), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1062), .B1(new_n794), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n787), .A2(G303), .B1(new_n781), .B2(G317), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n825), .B2(new_n786), .C1(new_n794), .C2(new_n802), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n774), .A2(G294), .B1(G283), .B2(new_n765), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT49), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1068), .A2(KEYINPUT49), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(KEYINPUT110), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n767), .A2(new_n481), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n388), .B(new_n1076), .C1(G326), .C2(new_n761), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT110), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1064), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n755), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n745), .A2(new_n692), .B1(G107), .B2(new_n211), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n233), .A2(new_n268), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n692), .ZN(new_n1084));
  AOI211_X1 g0884(.A(G45), .B(new_n1084), .C1(G68), .C2(G77), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n248), .A2(G50), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT50), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n749), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1082), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n744), .B1(new_n1089), .B2(new_n757), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n683), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n754), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1001), .A2(new_n991), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1081), .A2(new_n1092), .B1(new_n988), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1003), .B(new_n690), .C1(new_n731), .C2(new_n1093), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(G393));
  AND2_X1   g0896(.A1(new_n1003), .A2(new_n1026), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n690), .B1(new_n1003), .B2(new_n1026), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1023), .A2(new_n1025), .A3(new_n988), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n794), .A2(new_n831), .B1(new_n1063), .B2(new_n803), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT51), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n397), .B1(G143), .B2(new_n761), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n824), .B1(G77), .B2(new_n765), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n775), .C2(new_n203), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n249), .B2(new_n787), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1102), .B(new_n1106), .C1(new_n201), .C2(new_n786), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n808), .A2(G317), .B1(G311), .B2(new_n781), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT111), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT52), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n281), .B(new_n768), .C1(G322), .C2(new_n761), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n481), .B2(new_n764), .C1(new_n775), .C2(new_n798), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G294), .B2(new_n787), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1110), .B(new_n1113), .C1(new_n584), .C2(new_n786), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1109), .A2(KEYINPUT52), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n755), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1011), .A2(new_n754), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n756), .B1(new_n206), .B2(new_n211), .C1(new_n243), .C2(new_n749), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1117), .A2(new_n744), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1100), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1099), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G390));
  AOI21_X1  g0923(.A(new_n919), .B1(new_n864), .B2(new_n870), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT101), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n699), .A2(new_n657), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(new_n669), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n820), .A2(new_n327), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1130), .A2(new_n1131), .B1(new_n327), .B2(new_n678), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(new_n871), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n930), .B1(new_n866), .B2(new_n669), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n730), .A2(G330), .A3(new_n822), .A4(new_n870), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1128), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n927), .A2(G330), .A3(new_n928), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT112), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n660), .B1(new_n722), .B2(new_n940), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT112), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n928), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1124), .B1(new_n904), .B2(new_n918), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1137), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n380), .A2(new_n447), .A3(new_n1140), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(new_n634), .C1(new_n448), .C2(new_n922), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1140), .A2(new_n822), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n871), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1132), .A2(new_n1151), .A3(new_n1136), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n730), .A2(G330), .A3(new_n822), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1154), .A2(new_n871), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n864), .B1(new_n1155), .B2(new_n1143), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT113), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n871), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n1142), .A3(new_n1139), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT113), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n864), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1153), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1147), .B1(new_n1149), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1138), .A2(KEYINPUT112), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1141), .B1(new_n1140), .B2(new_n928), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(KEYINPUT113), .B(new_n865), .C1(new_n1166), .C2(new_n1158), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1160), .B1(new_n1159), .B2(new_n864), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1152), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1149), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1169), .A2(new_n1137), .A3(new_n1146), .A4(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1163), .A2(new_n690), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n753), .B1(new_n904), .B2(new_n918), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n347), .B1(new_n761), .B2(G125), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n201), .B2(new_n767), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT114), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n774), .A2(G150), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1176), .B(new_n1179), .C1(G159), .C2(new_n765), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT54), .B(G143), .Z(new_n1181));
  AOI22_X1  g0981(.A1(new_n787), .A2(new_n1181), .B1(new_n781), .B2(G132), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(new_n832), .C2(new_n786), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G128), .B2(new_n808), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n803), .A2(new_n481), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n764), .A2(new_n283), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n347), .B1(new_n760), .B2(new_n454), .C1(new_n203), .C2(new_n767), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n1185), .A2(new_n776), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n206), .B2(new_n788), .C1(new_n207), .C2(new_n786), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G283), .B2(new_n808), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n755), .B1(new_n1184), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n816), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1191), .B(new_n744), .C1(new_n249), .C2(new_n1192), .ZN(new_n1193));
  OR3_X1    g0993(.A1(new_n1173), .A2(KEYINPUT116), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT116), .B1(new_n1173), .B2(new_n1193), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1137), .A2(new_n1146), .A3(new_n988), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1172), .A2(new_n1199), .ZN(G378));
  AOI21_X1  g1000(.A(new_n742), .B1(new_n201), .B2(new_n816), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT121), .Z(new_n1202));
  NAND2_X1  g1002(.A1(new_n298), .A2(new_n303), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n264), .A2(new_n667), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1202), .B1(new_n1212), .B2(new_n753), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1063), .B2(new_n767), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n808), .A2(G125), .B1(G150), .B2(new_n765), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT119), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n781), .A2(G128), .B1(new_n774), .B2(new_n1181), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT118), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n980), .A2(G132), .B1(G137), .B2(new_n787), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT120), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1215), .B1(new_n1222), .B2(KEYINPUT59), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(KEYINPUT59), .B2(new_n1222), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n980), .A2(G97), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n388), .A2(G41), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n767), .A2(new_n202), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n976), .B1(G283), .B2(new_n761), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1057), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n306), .B2(new_n787), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n781), .A2(KEYINPUT117), .A3(G107), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT117), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n803), .B2(new_n207), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1225), .A2(new_n1230), .A3(new_n1231), .A4(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G116), .B2(new_n808), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT58), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1226), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1237), .B(new_n795), .C1(G33), .C2(G41), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1235), .A2(KEYINPUT58), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1224), .A2(new_n1236), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1213), .B1(new_n1240), .B2(new_n755), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n931), .A2(new_n936), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n937), .A2(new_n938), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1242), .A2(new_n1212), .A3(G330), .A4(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1212), .B1(new_n939), .B2(G330), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n921), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1242), .A2(G330), .A3(new_n1243), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1212), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1250), .A2(new_n920), .A3(new_n892), .A4(new_n1244), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1241), .B1(new_n1252), .B2(new_n988), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1170), .B1(new_n1147), .B2(new_n1162), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT57), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n690), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT57), .B1(new_n1254), .B2(new_n1252), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1253), .B1(new_n1258), .B2(new_n1259), .ZN(G375));
  NAND2_X1  g1060(.A1(new_n1162), .A2(new_n1149), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1029), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n744), .B1(G68), .B2(new_n1192), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1059), .B1(new_n803), .B2(new_n798), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT123), .Z(new_n1266));
  OAI21_X1  g1066(.A(new_n347), .B1(new_n767), .B2(new_n283), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT122), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n775), .A2(new_n206), .B1(new_n584), .B2(new_n760), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(G107), .C2(new_n787), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1266), .B(new_n1270), .C1(new_n481), .C2(new_n786), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n794), .A2(new_n454), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n794), .A2(new_n835), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n980), .A2(new_n1181), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n787), .A2(G150), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n781), .A2(G137), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n397), .B1(G128), .B2(new_n761), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1277), .B(new_n1227), .C1(new_n795), .C2(new_n764), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G159), .B2(new_n774), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .A4(new_n1279), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n1271), .A2(new_n1272), .B1(new_n1273), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1264), .B1(new_n1281), .B2(new_n755), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n871), .A2(new_n752), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1162), .B2(new_n987), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1263), .A2(new_n1286), .ZN(G381));
  NOR2_X1   g1087(.A1(G393), .A2(G396), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n859), .A3(new_n1122), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(G387), .A2(G381), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n689), .B1(new_n1262), .B2(new_n1147), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1198), .B1(new_n1291), .B2(new_n1171), .ZN(new_n1292));
  INV_X1    g1092(.A(G375), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1292), .A3(new_n1293), .ZN(G407));
  NAND2_X1  g1094(.A1(new_n668), .A2(G213), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1293), .A2(new_n1292), .A3(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(G407), .A2(G213), .A3(new_n1297), .ZN(G409));
  AOI21_X1  g1098(.A(new_n814), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1288), .A2(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1051), .A2(new_n1122), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1051), .A2(new_n1122), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1053), .A2(new_n1054), .A3(new_n1122), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1053), .A2(KEYINPUT124), .A3(new_n1054), .A4(new_n1122), .ZN(new_n1307));
  OAI22_X1  g1107(.A1(new_n1288), .A2(new_n1299), .B1(new_n1051), .B2(new_n1122), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AND4_X1   g1109(.A1(KEYINPUT125), .A2(new_n1306), .A3(new_n1307), .A4(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1308), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT125), .B1(new_n1311), .B2(new_n1307), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1303), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1296), .A2(G2897), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1317), .A2(KEYINPUT60), .A3(new_n1149), .A4(new_n1152), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n690), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT60), .B1(new_n1162), .B2(new_n1149), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1261), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(G384), .B1(new_n1323), .B2(new_n1286), .ZN(new_n1324));
  AOI211_X1 g1124(.A(new_n859), .B(new_n1285), .C1(new_n1320), .C2(new_n1322), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1316), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1170), .B(new_n1153), .C1(new_n1157), .C2(new_n1161), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(KEYINPUT60), .B2(new_n1262), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1286), .B1(new_n1328), .B2(new_n1319), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n859), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1323), .A2(G384), .A3(new_n1286), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1331), .A3(new_n1315), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1326), .A2(new_n1332), .ZN(new_n1333));
  OAI211_X1 g1133(.A(G378), .B(new_n1253), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1254), .A2(new_n1029), .A3(new_n1252), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1253), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1292), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1296), .B1(new_n1334), .B2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1314), .B1(new_n1333), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT62), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1334), .A2(new_n1337), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1342));
  AND4_X1   g1142(.A1(new_n1340), .A2(new_n1341), .A3(new_n1295), .A4(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1340), .B1(new_n1338), .B2(new_n1342), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1339), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1330), .A2(new_n1331), .A3(new_n1315), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1315), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1341), .A2(new_n1295), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT61), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT63), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1351), .B1(new_n1349), .B2(new_n1352), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1350), .A2(new_n1313), .A3(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1338), .A2(KEYINPUT63), .A3(new_n1342), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(KEYINPUT126), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT126), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1338), .A2(new_n1357), .A3(KEYINPUT63), .A4(new_n1342), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1356), .A2(new_n1358), .ZN(new_n1359));
  OAI22_X1  g1159(.A1(new_n1313), .A2(new_n1345), .B1(new_n1354), .B2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(new_n1313), .A2(KEYINPUT127), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(G375), .A2(new_n1292), .ZN(new_n1362));
  AND3_X1   g1162(.A1(new_n1362), .A2(new_n1334), .A3(new_n1352), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1352), .B1(new_n1362), .B2(new_n1334), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT127), .ZN(new_n1367));
  OAI211_X1 g1167(.A(new_n1367), .B(new_n1303), .C1(new_n1310), .C2(new_n1312), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1361), .A2(new_n1366), .A3(new_n1368), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1365), .A2(new_n1313), .A3(KEYINPUT127), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(G402));
endmodule


