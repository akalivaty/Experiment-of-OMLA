

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809;

  XNOR2_X1 U374 ( .A(G143), .B(G131), .ZN(n500) );
  XNOR2_X2 U375 ( .A(n435), .B(n482), .ZN(n683) );
  NAND2_X1 U376 ( .A1(n453), .A2(n450), .ZN(n455) );
  XNOR2_X1 U377 ( .A(n435), .B(n534), .ZN(n689) );
  XNOR2_X2 U378 ( .A(n404), .B(n682), .ZN(n684) );
  XNOR2_X2 U379 ( .A(n605), .B(KEYINPUT32), .ZN(n694) );
  NOR2_X1 U380 ( .A1(n806), .A2(n807), .ZN(n398) );
  XNOR2_X2 U381 ( .A(n632), .B(KEYINPUT30), .ZN(n409) );
  NAND2_X1 U382 ( .A1(n353), .A2(n393), .ZN(n391) );
  AND2_X1 U383 ( .A1(n694), .A2(n608), .ZN(n353) );
  XNOR2_X2 U384 ( .A(n365), .B(n688), .ZN(n690) );
  XNOR2_X2 U385 ( .A(n488), .B(KEYINPUT19), .ZN(n489) );
  XNOR2_X2 U386 ( .A(G902), .B(KEYINPUT15), .ZN(n667) );
  XOR2_X1 U387 ( .A(KEYINPUT99), .B(KEYINPUT80), .Z(n540) );
  INV_X1 U388 ( .A(G237), .ZN(n491) );
  NOR2_X1 U389 ( .A1(n618), .A2(n738), .ZN(n638) );
  INV_X1 U390 ( .A(KEYINPUT64), .ZN(n473) );
  AND2_X2 U391 ( .A1(n646), .A2(n753), .ZN(n636) );
  AND2_X2 U392 ( .A1(n371), .A2(n372), .ZN(n453) );
  NAND2_X2 U393 ( .A1(n615), .A2(n614), .ZN(n617) );
  AND2_X2 U394 ( .A1(n599), .A2(n598), .ZN(n615) );
  XNOR2_X1 U395 ( .A(n644), .B(KEYINPUT36), .ZN(n363) );
  INV_X1 U396 ( .A(n722), .ZN(n725) );
  AND2_X1 U397 ( .A1(n658), .A2(KEYINPUT78), .ZN(n357) );
  NOR2_X2 U398 ( .A1(n363), .A2(n602), .ZN(n731) );
  AND2_X1 U399 ( .A1(n649), .A2(n648), .ZN(n721) );
  XNOR2_X1 U400 ( .A(n375), .B(n368), .ZN(n753) );
  AND2_X1 U401 ( .A1(n618), .A2(n575), .ZN(n734) );
  OR2_X1 U402 ( .A1(G902), .A2(n776), .ZN(n526) );
  XNOR2_X1 U403 ( .A(n514), .B(n515), .ZN(n557) );
  INV_X1 U404 ( .A(KEYINPUT33), .ZN(n388) );
  INV_X1 U405 ( .A(KEYINPUT90), .ZN(n370) );
  INV_X1 U406 ( .A(KEYINPUT2), .ZN(n426) );
  INV_X1 U407 ( .A(KEYINPUT41), .ZN(n366) );
  NAND2_X1 U408 ( .A1(n433), .A2(n469), .ZN(n432) );
  NOR2_X1 U409 ( .A1(n429), .A2(n426), .ZN(n672) );
  AND2_X1 U410 ( .A1(n354), .A2(n449), .ZN(n372) );
  XNOR2_X1 U411 ( .A(n396), .B(n386), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n731), .B(n370), .ZN(n362) );
  XNOR2_X1 U413 ( .A(n647), .B(KEYINPUT107), .ZN(n649) );
  XNOR2_X1 U414 ( .A(n367), .B(n366), .ZN(n767) );
  NAND2_X1 U415 ( .A1(n629), .A2(n628), .ZN(n460) );
  NAND2_X1 U416 ( .A1(n753), .A2(n383), .ZN(n367) );
  XNOR2_X1 U417 ( .A(n389), .B(n388), .ZN(n766) );
  BUF_X1 U418 ( .A(n590), .Z(n735) );
  AND2_X1 U419 ( .A1(n734), .A2(n640), .ZN(n390) );
  XNOR2_X1 U420 ( .A(G478), .B(n526), .ZN(n594) );
  XNOR2_X1 U421 ( .A(n579), .B(n536), .ZN(n590) );
  NOR2_X1 U422 ( .A1(n624), .A2(n623), .ZN(n642) );
  BUF_X1 U423 ( .A(n689), .Z(n365) );
  XOR2_X1 U424 ( .A(G140), .B(G113), .Z(n501) );
  XNOR2_X1 U425 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n502) );
  INV_X1 U426 ( .A(KEYINPUT38), .ZN(n368) );
  XOR2_X1 U427 ( .A(KEYINPUT16), .B(KEYINPUT77), .Z(n471) );
  XOR2_X1 U428 ( .A(G137), .B(G140), .Z(n552) );
  NAND2_X1 U429 ( .A1(n354), .A2(n376), .ZN(n429) );
  NAND2_X1 U430 ( .A1(n356), .A2(n355), .ZN(n361) );
  INV_X1 U431 ( .A(n721), .ZN(n355) );
  NAND2_X1 U432 ( .A1(n659), .A2(n357), .ZN(n356) );
  NAND2_X1 U433 ( .A1(n359), .A2(n358), .ZN(n364) );
  NAND2_X1 U434 ( .A1(n439), .A2(n430), .ZN(n358) );
  NAND2_X1 U435 ( .A1(n361), .A2(n360), .ZN(n359) );
  NAND2_X1 U436 ( .A1(n721), .A2(KEYINPUT78), .ZN(n360) );
  NAND2_X1 U437 ( .A1(n364), .A2(n362), .ZN(n400) );
  NAND2_X1 U438 ( .A1(n409), .A2(n634), .ZN(n635) );
  INV_X2 U439 ( .A(KEYINPUT74), .ZN(n437) );
  INV_X1 U440 ( .A(n375), .ZN(n630) );
  INV_X1 U441 ( .A(n780), .ZN(n369) );
  NAND2_X1 U442 ( .A1(n671), .A2(KEYINPUT88), .ZN(n371) );
  INV_X1 U443 ( .A(n576), .ZN(n373) );
  BUF_X1 U444 ( .A(n728), .Z(n374) );
  XNOR2_X1 U445 ( .A(n578), .B(KEYINPUT31), .ZN(n728) );
  NAND2_X2 U446 ( .A1(n487), .A2(n752), .ZN(n490) );
  BUF_X1 U447 ( .A(n487), .Z(n375) );
  XNOR2_X2 U448 ( .A(n490), .B(n489), .ZN(n650) );
  XNOR2_X2 U449 ( .A(n617), .B(n616), .ZN(n671) );
  XNOR2_X1 U450 ( .A(KEYINPUT69), .B(G101), .ZN(n479) );
  XNOR2_X1 U451 ( .A(n419), .B(n394), .ZN(n393) );
  XNOR2_X1 U452 ( .A(KEYINPUT35), .B(n600), .ZN(n394) );
  INV_X1 U453 ( .A(KEYINPUT70), .ZN(n600) );
  NOR2_X1 U454 ( .A1(n454), .A2(n387), .ZN(n449) );
  XNOR2_X1 U455 ( .A(n551), .B(n438), .ZN(n793) );
  INV_X1 U456 ( .A(n552), .ZN(n438) );
  XOR2_X1 U457 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n475) );
  AND2_X1 U458 ( .A1(n766), .A2(n385), .ZN(n417) );
  NOR2_X1 U459 ( .A1(G902), .A2(n549), .ZN(n413) );
  XNOR2_X1 U460 ( .A(n401), .B(n550), .ZN(n619) );
  INV_X1 U461 ( .A(KEYINPUT78), .ZN(n430) );
  XNOR2_X1 U462 ( .A(n400), .B(n431), .ZN(n399) );
  INV_X1 U463 ( .A(KEYINPUT72), .ZN(n431) );
  XNOR2_X1 U464 ( .A(n398), .B(KEYINPUT46), .ZN(n397) );
  INV_X1 U465 ( .A(KEYINPUT65), .ZN(n467) );
  XNOR2_X1 U466 ( .A(G116), .B(KEYINPUT5), .ZN(n542) );
  XOR2_X1 U467 ( .A(KEYINPUT86), .B(KEYINPUT8), .Z(n515) );
  OR2_X1 U468 ( .A1(n670), .A2(KEYINPUT65), .ZN(n466) );
  XNOR2_X1 U469 ( .A(G104), .B(G122), .ZN(n503) );
  NAND2_X1 U470 ( .A1(n486), .A2(G214), .ZN(n752) );
  XNOR2_X1 U471 ( .A(n513), .B(n512), .ZN(n595) );
  NAND2_X1 U472 ( .A1(n445), .A2(n448), .ZN(n444) );
  NAND2_X1 U473 ( .A1(n447), .A2(n564), .ZN(n446) );
  XNOR2_X1 U474 ( .A(G110), .B(G107), .ZN(n480) );
  XNOR2_X1 U475 ( .A(G128), .B(G119), .ZN(n558) );
  XNOR2_X1 U476 ( .A(n793), .B(n555), .ZN(n556) );
  XNOR2_X1 U477 ( .A(G134), .B(G107), .ZN(n516) );
  XOR2_X1 U478 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n517) );
  INV_X1 U479 ( .A(n429), .ZN(n427) );
  NAND2_X1 U480 ( .A1(n416), .A2(n420), .ZN(n419) );
  NOR2_X1 U481 ( .A1(n418), .A2(n417), .ZN(n416) );
  NAND2_X1 U482 ( .A1(G902), .A2(n549), .ZN(n414) );
  INV_X1 U483 ( .A(KEYINPUT22), .ZN(n464) );
  INV_X1 U484 ( .A(n800), .ZN(n428) );
  OR2_X1 U485 ( .A1(n799), .A2(G952), .ZN(n704) );
  XNOR2_X1 U486 ( .A(n442), .B(n441), .ZN(n807) );
  INV_X1 U487 ( .A(KEYINPUT42), .ZN(n441) );
  OR2_X1 U488 ( .A1(n767), .A2(n460), .ZN(n442) );
  NAND2_X1 U489 ( .A1(n459), .A2(n458), .ZN(n723) );
  INV_X1 U490 ( .A(n655), .ZN(n458) );
  AND2_X1 U491 ( .A1(n666), .A2(n808), .ZN(n376) );
  AND2_X1 U492 ( .A1(n753), .A2(n752), .ZN(n377) );
  AND2_X1 U493 ( .A1(n377), .A2(n656), .ZN(n378) );
  XOR2_X1 U494 ( .A(n485), .B(n484), .Z(n379) );
  NOR2_X1 U495 ( .A1(n735), .A2(n640), .ZN(n380) );
  AND2_X1 U496 ( .A1(n673), .A2(n467), .ZN(n381) );
  AND2_X1 U497 ( .A1(n440), .A2(n575), .ZN(n382) );
  INV_X1 U498 ( .A(G902), .ZN(n564) );
  INV_X1 U499 ( .A(n755), .ZN(n440) );
  AND2_X1 U500 ( .A1(n440), .A2(n752), .ZN(n383) );
  NOR2_X1 U501 ( .A1(n735), .A2(n570), .ZN(n384) );
  INV_X1 U502 ( .A(n376), .ZN(n454) );
  AND2_X1 U503 ( .A1(n717), .A2(n722), .ZN(n756) );
  XOR2_X1 U504 ( .A(n593), .B(KEYINPUT34), .Z(n385) );
  XNOR2_X1 U505 ( .A(n660), .B(KEYINPUT89), .ZN(n386) );
  AND2_X1 U506 ( .A1(n667), .A2(KEYINPUT88), .ZN(n387) );
  NAND2_X1 U507 ( .A1(n590), .A2(n390), .ZN(n389) );
  OR2_X2 U508 ( .A1(n443), .A2(n444), .ZN(n579) );
  NAND2_X1 U509 ( .A1(n391), .A2(n606), .ZN(n613) );
  XNOR2_X2 U510 ( .A(n395), .B(n379), .ZN(n487) );
  NAND2_X1 U511 ( .A1(n683), .A2(n667), .ZN(n395) );
  NAND2_X1 U512 ( .A1(n399), .A2(n397), .ZN(n396) );
  INV_X1 U513 ( .A(n401), .ZN(n576) );
  XNOR2_X1 U514 ( .A(n401), .B(n572), .ZN(n640) );
  NAND2_X1 U515 ( .A1(n734), .A2(n373), .ZN(n580) );
  NAND2_X1 U516 ( .A1(n743), .A2(n373), .ZN(n744) );
  NAND2_X2 U517 ( .A1(n411), .A2(n415), .ZN(n401) );
  AND2_X1 U518 ( .A1(n412), .A2(n414), .ZN(n411) );
  NAND2_X1 U519 ( .A1(n689), .A2(n535), .ZN(n445) );
  NAND2_X1 U520 ( .A1(n422), .A2(n432), .ZN(n402) );
  NAND2_X1 U521 ( .A1(n422), .A2(n432), .ZN(n403) );
  NAND2_X2 U522 ( .A1(n422), .A2(n432), .ZN(n775) );
  BUF_X1 U523 ( .A(n683), .Z(n404) );
  NAND2_X1 U524 ( .A1(n453), .A2(n450), .ZN(n405) );
  NOR2_X1 U525 ( .A1(n592), .A2(n385), .ZN(n421) );
  XNOR2_X1 U526 ( .A(n410), .B(n472), .ZN(n788) );
  XNOR2_X1 U527 ( .A(n410), .B(n537), .ZN(n546) );
  NAND2_X1 U528 ( .A1(n452), .A2(n451), .ZN(n450) );
  XNOR2_X1 U529 ( .A(n419), .B(KEYINPUT35), .ZN(n406) );
  XNOR2_X1 U530 ( .A(n405), .B(KEYINPUT87), .ZN(n407) );
  BUF_X1 U531 ( .A(n797), .Z(n408) );
  XNOR2_X1 U532 ( .A(n455), .B(KEYINPUT87), .ZN(n434) );
  OR2_X2 U533 ( .A1(n728), .A2(n710), .ZN(n586) );
  INV_X1 U534 ( .A(n735), .ZN(n602) );
  NAND2_X1 U535 ( .A1(n457), .A2(n421), .ZN(n420) );
  NAND2_X1 U536 ( .A1(n456), .A2(n648), .ZN(n418) );
  XNOR2_X2 U537 ( .A(n462), .B(n461), .ZN(n410) );
  NAND2_X1 U538 ( .A1(n674), .A2(n413), .ZN(n412) );
  OR2_X1 U539 ( .A1(n674), .A2(G472), .ZN(n415) );
  AND2_X2 U540 ( .A1(n423), .A2(n425), .ZN(n422) );
  NAND2_X1 U541 ( .A1(n434), .A2(n381), .ZN(n423) );
  NAND2_X1 U542 ( .A1(n424), .A2(n465), .ZN(n425) );
  NAND2_X1 U543 ( .A1(n468), .A2(n467), .ZN(n424) );
  NAND2_X1 U544 ( .A1(n369), .A2(n427), .ZN(n765) );
  XNOR2_X1 U545 ( .A(n429), .B(n428), .ZN(n798) );
  XNOR2_X2 U546 ( .A(n547), .B(n481), .ZN(n435) );
  XNOR2_X2 U547 ( .A(n797), .B(n479), .ZN(n547) );
  XNOR2_X2 U548 ( .A(n521), .B(KEYINPUT4), .ZN(n797) );
  INV_X1 U549 ( .A(n407), .ZN(n433) );
  NAND2_X1 U550 ( .A1(n436), .A2(n380), .ZN(n573) );
  NAND2_X1 U551 ( .A1(n436), .A2(n604), .ZN(n605) );
  NAND2_X1 U552 ( .A1(n436), .A2(n384), .ZN(n608) );
  XNOR2_X2 U553 ( .A(n530), .B(n464), .ZN(n436) );
  XNOR2_X2 U554 ( .A(n437), .B(G119), .ZN(n462) );
  NOR2_X2 U555 ( .A1(n635), .A2(n579), .ZN(n646) );
  NAND2_X1 U556 ( .A1(n659), .A2(n658), .ZN(n439) );
  NOR2_X1 U557 ( .A1(n689), .A2(n446), .ZN(n443) );
  INV_X1 U558 ( .A(n535), .ZN(n447) );
  NAND2_X1 U559 ( .A1(n535), .A2(G902), .ZN(n448) );
  NOR2_X1 U560 ( .A1(n667), .A2(KEYINPUT88), .ZN(n451) );
  INV_X1 U561 ( .A(n671), .ZN(n452) );
  NAND2_X1 U562 ( .A1(n592), .A2(n385), .ZN(n456) );
  INV_X1 U563 ( .A(n766), .ZN(n457) );
  INV_X1 U564 ( .A(n460), .ZN(n459) );
  NOR2_X1 U565 ( .A1(n651), .A2(n460), .ZN(n652) );
  XNOR2_X1 U566 ( .A(n547), .B(n548), .ZN(n674) );
  XNOR2_X2 U567 ( .A(G113), .B(KEYINPUT3), .ZN(n461) );
  XNOR2_X2 U568 ( .A(n795), .B(G146), .ZN(n537) );
  XNOR2_X2 U569 ( .A(G131), .B(G134), .ZN(n795) );
  XNOR2_X2 U570 ( .A(n463), .B(G143), .ZN(n521) );
  XNOR2_X2 U571 ( .A(G128), .B(KEYINPUT84), .ZN(n463) );
  NAND2_X1 U572 ( .A1(n673), .A2(n466), .ZN(n465) );
  INV_X1 U573 ( .A(n673), .ZN(n468) );
  AND2_X1 U574 ( .A1(n670), .A2(KEYINPUT65), .ZN(n469) );
  XNOR2_X2 U575 ( .A(n563), .B(n562), .ZN(n695) );
  BUF_X1 U576 ( .A(n591), .Z(n582) );
  BUF_X1 U577 ( .A(n521), .Z(n523) );
  OR2_X1 U578 ( .A1(n642), .A2(n641), .ZN(n470) );
  INV_X1 U579 ( .A(KEYINPUT47), .ZN(n653) );
  INV_X1 U580 ( .A(G137), .ZN(n541) );
  XNOR2_X1 U581 ( .A(n542), .B(n541), .ZN(n543) );
  INV_X1 U582 ( .A(n752), .ZN(n641) );
  XNOR2_X1 U583 ( .A(n544), .B(n543), .ZN(n545) );
  NOR2_X2 U584 ( .A1(n643), .A2(n470), .ZN(n662) );
  INV_X1 U585 ( .A(KEYINPUT1), .ZN(n536) );
  XNOR2_X1 U586 ( .A(n522), .B(n471), .ZN(n472) );
  XNOR2_X1 U587 ( .A(n511), .B(G475), .ZN(n512) );
  BUF_X1 U588 ( .A(n680), .Z(n681) );
  XOR2_X1 U589 ( .A(G116), .B(G122), .Z(n522) );
  XNOR2_X2 U590 ( .A(n473), .B(G953), .ZN(n799) );
  NAND2_X1 U591 ( .A1(G224), .A2(n799), .ZN(n474) );
  XNOR2_X1 U592 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X2 U593 ( .A(G146), .B(G125), .ZN(n507) );
  XNOR2_X1 U594 ( .A(KEYINPUT18), .B(n507), .ZN(n476) );
  XNOR2_X1 U595 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U596 ( .A(n788), .B(n478), .ZN(n482) );
  XNOR2_X1 U597 ( .A(n480), .B(G104), .ZN(n786) );
  XNOR2_X1 U598 ( .A(n786), .B(KEYINPUT75), .ZN(n481) );
  NAND2_X1 U599 ( .A1(n564), .A2(n491), .ZN(n486) );
  NAND2_X1 U600 ( .A1(n486), .A2(G210), .ZN(n485) );
  INV_X1 U601 ( .A(KEYINPUT93), .ZN(n483) );
  XNOR2_X1 U602 ( .A(n483), .B(KEYINPUT94), .ZN(n484) );
  INV_X1 U603 ( .A(KEYINPUT67), .ZN(n488) );
  XOR2_X1 U604 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n494) );
  INV_X1 U605 ( .A(n491), .ZN(n492) );
  NAND2_X1 U606 ( .A1(G234), .A2(n492), .ZN(n493) );
  XNOR2_X1 U607 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U608 ( .A1(G952), .A2(n495), .ZN(n764) );
  OR2_X1 U609 ( .A1(n764), .A2(G953), .ZN(n620) );
  NAND2_X1 U610 ( .A1(G902), .A2(n495), .ZN(n621) );
  INV_X1 U611 ( .A(G898), .ZN(n783) );
  NAND2_X1 U612 ( .A1(G953), .A2(n783), .ZN(n790) );
  OR2_X1 U613 ( .A1(n621), .A2(n790), .ZN(n496) );
  NAND2_X1 U614 ( .A1(n620), .A2(n496), .ZN(n497) );
  NAND2_X1 U615 ( .A1(n650), .A2(n497), .ZN(n499) );
  INV_X1 U616 ( .A(KEYINPUT0), .ZN(n498) );
  XNOR2_X2 U617 ( .A(n499), .B(n498), .ZN(n591) );
  XNOR2_X1 U618 ( .A(n501), .B(n500), .ZN(n506) );
  INV_X1 U619 ( .A(n502), .ZN(n504) );
  XNOR2_X1 U620 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U621 ( .A(n506), .B(n505), .Z(n510) );
  NOR2_X2 U622 ( .A1(G953), .A2(G237), .ZN(n538) );
  NAND2_X1 U623 ( .A1(G214), .A2(n538), .ZN(n508) );
  XNOR2_X1 U624 ( .A(KEYINPUT10), .B(n507), .ZN(n551) );
  XNOR2_X1 U625 ( .A(n508), .B(n551), .ZN(n509) );
  XNOR2_X1 U626 ( .A(n510), .B(n509), .ZN(n701) );
  NOR2_X1 U627 ( .A1(G902), .A2(n701), .ZN(n513) );
  XNOR2_X1 U628 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n511) );
  NAND2_X1 U629 ( .A1(G234), .A2(n799), .ZN(n514) );
  NAND2_X1 U630 ( .A1(G217), .A2(n557), .ZN(n520) );
  XNOR2_X1 U631 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U632 ( .A(n518), .B(KEYINPUT7), .Z(n519) );
  XNOR2_X1 U633 ( .A(n520), .B(n519), .ZN(n525) );
  XOR2_X1 U634 ( .A(n523), .B(n522), .Z(n524) );
  XNOR2_X1 U635 ( .A(n525), .B(n524), .ZN(n776) );
  OR2_X1 U636 ( .A1(n595), .A2(n594), .ZN(n755) );
  NAND2_X1 U637 ( .A1(n667), .A2(G234), .ZN(n527) );
  XNOR2_X1 U638 ( .A(n527), .B(KEYINPUT20), .ZN(n565) );
  AND2_X1 U639 ( .A1(n565), .A2(G221), .ZN(n529) );
  INV_X1 U640 ( .A(KEYINPUT21), .ZN(n528) );
  XNOR2_X1 U641 ( .A(n529), .B(n528), .ZN(n738) );
  INV_X1 U642 ( .A(n738), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n591), .A2(n382), .ZN(n530) );
  XOR2_X1 U644 ( .A(n552), .B(KEYINPUT81), .Z(n532) );
  NAND2_X1 U645 ( .A1(n799), .A2(G227), .ZN(n531) );
  XNOR2_X1 U646 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U647 ( .A(n537), .B(n533), .ZN(n534) );
  XNOR2_X1 U648 ( .A(KEYINPUT73), .B(G469), .ZN(n535) );
  NAND2_X1 U649 ( .A1(n538), .A2(G210), .ZN(n539) );
  XNOR2_X1 U650 ( .A(n540), .B(n539), .ZN(n544) );
  XNOR2_X1 U651 ( .A(n546), .B(n545), .ZN(n548) );
  INV_X1 U652 ( .A(G472), .ZN(n549) );
  INV_X1 U653 ( .A(KEYINPUT105), .ZN(n550) );
  XOR2_X1 U654 ( .A(KEYINPUT23), .B(KEYINPUT97), .Z(n554) );
  XNOR2_X1 U655 ( .A(G110), .B(KEYINPUT95), .ZN(n553) );
  XNOR2_X1 U656 ( .A(n554), .B(n553), .ZN(n555) );
  INV_X1 U657 ( .A(n556), .ZN(n563) );
  NAND2_X1 U658 ( .A1(G221), .A2(n557), .ZN(n561) );
  XOR2_X1 U659 ( .A(KEYINPUT24), .B(KEYINPUT96), .Z(n559) );
  XNOR2_X1 U660 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U661 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U662 ( .A1(n695), .A2(n564), .ZN(n569) );
  XOR2_X1 U663 ( .A(KEYINPUT25), .B(KEYINPUT98), .Z(n567) );
  NAND2_X1 U664 ( .A1(G217), .A2(n565), .ZN(n566) );
  XNOR2_X1 U665 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X2 U666 ( .A(n569), .B(n568), .ZN(n618) );
  INV_X1 U667 ( .A(n618), .ZN(n739) );
  NAND2_X1 U668 ( .A1(n619), .A2(n739), .ZN(n570) );
  XNOR2_X1 U669 ( .A(n608), .B(G110), .ZN(G12) );
  INV_X1 U670 ( .A(KEYINPUT103), .ZN(n571) );
  XNOR2_X1 U671 ( .A(n571), .B(KEYINPUT6), .ZN(n572) );
  XNOR2_X1 U672 ( .A(n573), .B(KEYINPUT91), .ZN(n574) );
  NAND2_X1 U673 ( .A1(n574), .A2(n618), .ZN(n680) );
  AND2_X1 U674 ( .A1(n576), .A2(n734), .ZN(n577) );
  AND2_X1 U675 ( .A1(n735), .A2(n577), .ZN(n746) );
  NAND2_X1 U676 ( .A1(n582), .A2(n746), .ZN(n578) );
  NOR2_X1 U677 ( .A1(n580), .A2(n579), .ZN(n581) );
  AND2_X1 U678 ( .A1(n582), .A2(n581), .ZN(n710) );
  XOR2_X1 U679 ( .A(n595), .B(KEYINPUT101), .Z(n585) );
  INV_X1 U680 ( .A(n585), .ZN(n583) );
  NAND2_X1 U681 ( .A1(n583), .A2(n594), .ZN(n717) );
  INV_X1 U682 ( .A(n594), .ZN(n584) );
  NAND2_X1 U683 ( .A1(n585), .A2(n584), .ZN(n722) );
  INV_X1 U684 ( .A(n756), .ZN(n656) );
  NAND2_X1 U685 ( .A1(n586), .A2(n656), .ZN(n587) );
  NAND2_X1 U686 ( .A1(n680), .A2(n587), .ZN(n589) );
  INV_X1 U687 ( .A(KEYINPUT104), .ZN(n588) );
  XNOR2_X1 U688 ( .A(n589), .B(n588), .ZN(n599) );
  INV_X1 U689 ( .A(n591), .ZN(n592) );
  INV_X1 U690 ( .A(KEYINPUT76), .ZN(n593) );
  AND2_X1 U691 ( .A1(n595), .A2(n594), .ZN(n648) );
  NAND2_X1 U692 ( .A1(n406), .A2(KEYINPUT44), .ZN(n597) );
  INV_X1 U693 ( .A(KEYINPUT92), .ZN(n596) );
  NAND2_X1 U694 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U695 ( .A(n640), .B(KEYINPUT83), .ZN(n601) );
  NAND2_X1 U696 ( .A1(n601), .A2(n739), .ZN(n603) );
  NOR2_X1 U697 ( .A1(n603), .A2(n602), .ZN(n604) );
  INV_X1 U698 ( .A(KEYINPUT44), .ZN(n606) );
  AND2_X1 U699 ( .A1(KEYINPUT70), .A2(KEYINPUT44), .ZN(n607) );
  AND2_X1 U700 ( .A1(n608), .A2(n607), .ZN(n609) );
  AND2_X1 U701 ( .A1(n694), .A2(n609), .ZN(n611) );
  NAND2_X1 U702 ( .A1(n406), .A2(KEYINPUT92), .ZN(n610) );
  NAND2_X1 U703 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U704 ( .A1(n613), .A2(n612), .ZN(n614) );
  INV_X1 U705 ( .A(KEYINPUT45), .ZN(n616) );
  INV_X1 U706 ( .A(n619), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n638), .A2(n631), .ZN(n625) );
  INV_X1 U708 ( .A(n620), .ZN(n624) );
  OR2_X1 U709 ( .A1(n799), .A2(n621), .ZN(n622) );
  NOR2_X1 U710 ( .A1(G900), .A2(n622), .ZN(n623) );
  NOR2_X1 U711 ( .A1(n625), .A2(n642), .ZN(n626) );
  XNOR2_X1 U712 ( .A(n626), .B(KEYINPUT28), .ZN(n629) );
  INV_X1 U713 ( .A(KEYINPUT108), .ZN(n627) );
  XNOR2_X1 U714 ( .A(n579), .B(n627), .ZN(n628) );
  AND2_X1 U715 ( .A1(n631), .A2(n752), .ZN(n632) );
  INV_X1 U716 ( .A(n734), .ZN(n633) );
  NOR2_X1 U717 ( .A1(n633), .A2(n642), .ZN(n634) );
  XNOR2_X1 U718 ( .A(n636), .B(KEYINPUT39), .ZN(n661) );
  NOR2_X1 U719 ( .A1(n661), .A2(n722), .ZN(n637) );
  XNOR2_X1 U720 ( .A(n637), .B(KEYINPUT40), .ZN(n806) );
  AND2_X1 U721 ( .A1(n725), .A2(n638), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n643) );
  INV_X1 U723 ( .A(n630), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n662), .A2(n645), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  INV_X1 U726 ( .A(n650), .ZN(n655) );
  OR2_X1 U727 ( .A1(n655), .A2(n756), .ZN(n651) );
  NOR2_X1 U728 ( .A1(KEYINPUT85), .A2(n652), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(n653), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n723), .A2(n656), .ZN(n657) );
  NAND2_X1 U731 ( .A1(KEYINPUT85), .A2(n657), .ZN(n658) );
  XOR2_X1 U732 ( .A(KEYINPUT48), .B(KEYINPUT71), .Z(n660) );
  NOR2_X1 U733 ( .A1(n717), .A2(n661), .ZN(n733) );
  INV_X1 U734 ( .A(n733), .ZN(n666) );
  NAND2_X1 U735 ( .A1(n662), .A2(n602), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n663), .B(KEYINPUT43), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n664), .A2(n630), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(KEYINPUT106), .ZN(n808) );
  INV_X1 U739 ( .A(n667), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n668), .A2(KEYINPUT2), .ZN(n669) );
  XNOR2_X1 U741 ( .A(n669), .B(KEYINPUT66), .ZN(n670) );
  BUF_X1 U742 ( .A(n671), .Z(n780) );
  NAND2_X1 U743 ( .A1(n672), .A2(n452), .ZN(n673) );
  NAND2_X1 U744 ( .A1(n403), .A2(G472), .ZN(n677) );
  BUF_X1 U745 ( .A(n674), .Z(n675) );
  XNOR2_X1 U746 ( .A(n675), .B(KEYINPUT62), .ZN(n676) );
  XNOR2_X1 U747 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U748 ( .A1(n678), .A2(n704), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n679), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U750 ( .A(n681), .B(G101), .ZN(G3) );
  NAND2_X1 U751 ( .A1(n775), .A2(G210), .ZN(n685) );
  XNOR2_X1 U752 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n682) );
  XNOR2_X1 U753 ( .A(n685), .B(n684), .ZN(n686) );
  INV_X1 U754 ( .A(n704), .ZN(n779) );
  NOR2_X2 U755 ( .A1(n686), .A2(n779), .ZN(n687) );
  XNOR2_X1 U756 ( .A(n687), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U757 ( .A1(n775), .A2(G469), .ZN(n691) );
  XOR2_X1 U758 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n688) );
  XNOR2_X1 U759 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X2 U760 ( .A1(n692), .A2(n779), .ZN(n693) );
  XNOR2_X1 U761 ( .A(n693), .B(KEYINPUT122), .ZN(G54) );
  XNOR2_X1 U762 ( .A(n694), .B(G119), .ZN(G21) );
  XOR2_X1 U763 ( .A(n406), .B(G122), .Z(G24) );
  NAND2_X1 U764 ( .A1(n402), .A2(G217), .ZN(n697) );
  XNOR2_X1 U765 ( .A(n695), .B(KEYINPUT124), .ZN(n696) );
  XNOR2_X1 U766 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U767 ( .A1(n698), .A2(n704), .ZN(n699) );
  XNOR2_X1 U768 ( .A(n699), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U769 ( .A1(n403), .A2(G475), .ZN(n703) );
  XOR2_X1 U770 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n700) );
  XNOR2_X1 U771 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U772 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n707) );
  XOR2_X1 U774 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n706) );
  XNOR2_X1 U775 ( .A(n707), .B(n706), .ZN(G60) );
  XOR2_X1 U776 ( .A(G104), .B(KEYINPUT109), .Z(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n725), .ZN(n708) );
  XNOR2_X1 U778 ( .A(n709), .B(n708), .ZN(G6) );
  INV_X1 U779 ( .A(n717), .ZN(n727) );
  NAND2_X1 U780 ( .A1(n710), .A2(n727), .ZN(n716) );
  XOR2_X1 U781 ( .A(KEYINPUT112), .B(KEYINPUT27), .Z(n712) );
  XNOR2_X1 U782 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n711) );
  XNOR2_X1 U783 ( .A(n712), .B(n711), .ZN(n714) );
  XOR2_X1 U784 ( .A(G107), .B(KEYINPUT26), .Z(n713) );
  XNOR2_X1 U785 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U786 ( .A(n716), .B(n715), .ZN(G9) );
  NOR2_X1 U787 ( .A1(n723), .A2(n717), .ZN(n719) );
  XNOR2_X1 U788 ( .A(KEYINPUT29), .B(KEYINPUT113), .ZN(n718) );
  XNOR2_X1 U789 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U790 ( .A(G128), .B(n720), .Z(G30) );
  XOR2_X1 U791 ( .A(G143), .B(n721), .Z(G45) );
  NOR2_X1 U792 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U793 ( .A(G146), .B(n724), .Z(G48) );
  NAND2_X1 U794 ( .A1(n374), .A2(n725), .ZN(n726) );
  XNOR2_X1 U795 ( .A(n726), .B(G113), .ZN(G15) );
  NAND2_X1 U796 ( .A1(n374), .A2(n727), .ZN(n729) );
  XNOR2_X1 U797 ( .A(n729), .B(KEYINPUT114), .ZN(n730) );
  XNOR2_X1 U798 ( .A(G116), .B(n730), .ZN(G18) );
  XNOR2_X1 U799 ( .A(n731), .B(G125), .ZN(n732) );
  XNOR2_X1 U800 ( .A(n732), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U801 ( .A(G134), .B(n733), .Z(G36) );
  OR2_X1 U802 ( .A1(n735), .A2(n734), .ZN(n737) );
  XOR2_X1 U803 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n736) );
  XNOR2_X1 U804 ( .A(n737), .B(n736), .ZN(n745) );
  NAND2_X1 U805 ( .A1(n739), .A2(n738), .ZN(n742) );
  XNOR2_X1 U806 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n740) );
  XNOR2_X1 U807 ( .A(n740), .B(KEYINPUT116), .ZN(n741) );
  XNOR2_X1 U808 ( .A(n742), .B(n741), .ZN(n743) );
  OR2_X1 U809 ( .A1(n745), .A2(n744), .ZN(n748) );
  INV_X1 U810 ( .A(n746), .ZN(n747) );
  AND2_X1 U811 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U812 ( .A(n749), .B(KEYINPUT119), .ZN(n750) );
  XNOR2_X1 U813 ( .A(KEYINPUT51), .B(n750), .ZN(n751) );
  NOR2_X1 U814 ( .A1(n767), .A2(n751), .ZN(n761) );
  NOR2_X1 U815 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U816 ( .A1(n755), .A2(n754), .ZN(n757) );
  NOR2_X1 U817 ( .A1(n757), .A2(n378), .ZN(n758) );
  NOR2_X1 U818 ( .A1(n758), .A2(n766), .ZN(n759) );
  XNOR2_X1 U819 ( .A(n759), .B(KEYINPUT120), .ZN(n760) );
  NOR2_X1 U820 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U821 ( .A(n762), .B(KEYINPUT52), .ZN(n763) );
  NOR2_X1 U822 ( .A1(n764), .A2(n763), .ZN(n771) );
  XNOR2_X1 U823 ( .A(n765), .B(KEYINPUT2), .ZN(n769) );
  NOR2_X1 U824 ( .A1(n767), .A2(n766), .ZN(n768) );
  OR2_X1 U825 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U826 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U827 ( .A(n772), .B(KEYINPUT121), .ZN(n773) );
  NOR2_X1 U828 ( .A1(G953), .A2(n773), .ZN(n774) );
  XNOR2_X1 U829 ( .A(KEYINPUT53), .B(n774), .ZN(G75) );
  NAND2_X1 U830 ( .A1(n402), .A2(G478), .ZN(n777) );
  XNOR2_X1 U831 ( .A(n776), .B(n777), .ZN(n778) );
  NOR2_X1 U832 ( .A1(n779), .A2(n778), .ZN(G63) );
  OR2_X1 U833 ( .A1(n780), .A2(G953), .ZN(n785) );
  NAND2_X1 U834 ( .A1(G953), .A2(G224), .ZN(n781) );
  XOR2_X1 U835 ( .A(KEYINPUT61), .B(n781), .Z(n782) );
  OR2_X1 U836 ( .A1(n783), .A2(n782), .ZN(n784) );
  AND2_X1 U837 ( .A1(n785), .A2(n784), .ZN(n792) );
  XOR2_X1 U838 ( .A(G101), .B(n786), .Z(n787) );
  XNOR2_X1 U839 ( .A(n788), .B(n787), .ZN(n789) );
  NAND2_X1 U840 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U841 ( .A(n792), .B(n791), .ZN(G69) );
  XOR2_X1 U842 ( .A(n793), .B(KEYINPUT126), .Z(n794) );
  XNOR2_X1 U843 ( .A(n795), .B(n794), .ZN(n796) );
  XOR2_X1 U844 ( .A(n408), .B(n796), .Z(n800) );
  NAND2_X1 U845 ( .A1(n799), .A2(n798), .ZN(n805) );
  XNOR2_X1 U846 ( .A(n800), .B(G227), .ZN(n801) );
  XNOR2_X1 U847 ( .A(n801), .B(KEYINPUT127), .ZN(n802) );
  NAND2_X1 U848 ( .A1(n802), .A2(G900), .ZN(n803) );
  NAND2_X1 U849 ( .A1(G953), .A2(n803), .ZN(n804) );
  NAND2_X1 U850 ( .A1(n805), .A2(n804), .ZN(G72) );
  XOR2_X1 U851 ( .A(n806), .B(G131), .Z(G33) );
  XOR2_X1 U852 ( .A(G137), .B(n807), .Z(G39) );
  XOR2_X1 U853 ( .A(G140), .B(n808), .Z(n809) );
  XNOR2_X1 U854 ( .A(KEYINPUT115), .B(n809), .ZN(G42) );
endmodule

