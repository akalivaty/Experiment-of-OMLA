//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n607, new_n608, new_n609, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n645, new_n646, new_n649, new_n650, new_n652, new_n653, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT65), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(new_n463), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT66), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n474), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT68), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n480), .A3(new_n477), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n473), .A2(new_n479), .A3(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n464), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n469), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  AND4_X1   g066(.A1(KEYINPUT69), .A2(new_n461), .A3(new_n463), .A4(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(new_n477), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n477), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI211_X1 g074(.A(KEYINPUT4), .B(new_n498), .C1(new_n469), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n496), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT71), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n509), .B1(new_n506), .B2(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n503), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT5), .B1(new_n514), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT72), .B1(new_n516), .B2(KEYINPUT73), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n508), .A2(new_n512), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(new_n519), .ZN(new_n525));
  INV_X1    g100(.A(new_n515), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n527), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n522), .B(new_n524), .C1(new_n503), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n528), .A2(new_n503), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n531), .A2(new_n532), .A3(new_n522), .A4(new_n524), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(G166));
  AOI22_X1  g109(.A1(new_n504), .A2(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(new_n527), .A3(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(G51), .A3(G543), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n523), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n514), .A2(G543), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n549), .A2(KEYINPUT72), .B1(G543), .B2(new_n518), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n508), .B(new_n512), .C1(new_n550), .C2(new_n515), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n547), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n503), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(G171));
  NAND3_X1  g130(.A1(new_n535), .A2(new_n527), .A3(G81), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n535), .A2(G43), .A3(G543), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n558), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n520), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n563), .A2(new_n564), .A3(G651), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n564), .B1(new_n563), .B2(G651), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n559), .A2(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT78), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n556), .A2(new_n557), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT77), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n563), .A2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT76), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n563), .A2(new_n564), .A3(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n568), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G860), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT79), .Z(G153));
  AND3_X1   g156(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G36), .ZN(G176));
  NAND2_X1  g158(.A1(G1), .A2(G3), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT8), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(G188));
  NAND4_X1  g161(.A1(new_n508), .A2(new_n512), .A3(G53), .A4(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT9), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(KEYINPUT80), .A3(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT9), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n523), .A2(new_n593), .A3(new_n594), .A4(G53), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT81), .B1(new_n587), .B2(KEYINPUT9), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n527), .A2(G65), .ZN(new_n599));
  NAND2_X1  g174(.A1(G78), .A2(G543), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT82), .Z(new_n601));
  AOI21_X1  g176(.A(new_n503), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n521), .A2(G91), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n598), .A2(new_n603), .A3(new_n604), .ZN(G299));
  OAI221_X1 g180(.A(new_n547), .B1(new_n548), .B2(new_n551), .C1(new_n553), .C2(new_n503), .ZN(G301));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n607));
  NOR2_X1   g182(.A1(G166), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(KEYINPUT83), .B1(new_n530), .B2(new_n533), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(G303));
  INV_X1    g185(.A(G74), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n503), .B1(new_n520), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n521), .B2(G87), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n535), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G49), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n523), .A2(KEYINPUT84), .A3(G49), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n613), .A2(new_n617), .A3(new_n618), .ZN(G288));
  NAND2_X1  g194(.A1(new_n521), .A2(G86), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n527), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G48), .ZN(new_n622));
  OAI221_X1 g197(.A(new_n620), .B1(new_n621), .B2(new_n503), .C1(new_n622), .C2(new_n615), .ZN(G305));
  AOI22_X1  g198(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(new_n503), .ZN(new_n625));
  INV_X1    g200(.A(G47), .ZN(new_n626));
  INV_X1    g201(.A(G85), .ZN(new_n627));
  OAI22_X1  g202(.A1(new_n615), .A2(new_n626), .B1(new_n551), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(G290));
  INV_X1    g205(.A(G92), .ZN(new_n631));
  OAI21_X1  g206(.A(KEYINPUT10), .B1(new_n551), .B2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G66), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(new_n525), .B2(new_n526), .ZN(new_n634));
  AND2_X1   g209(.A1(G79), .A2(G543), .ZN(new_n635));
  OAI21_X1  g210(.A(G651), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n523), .A2(G54), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT10), .ZN(new_n638));
  NAND4_X1  g213(.A1(new_n535), .A2(new_n527), .A3(new_n638), .A4(G92), .ZN(new_n639));
  NAND4_X1  g214(.A1(new_n632), .A2(new_n636), .A3(new_n637), .A4(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G868), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(G171), .B2(new_n641), .ZN(G284));
  OAI21_X1  g218(.A(new_n642), .B1(G171), .B2(new_n641), .ZN(G321));
  NAND2_X1  g219(.A1(G286), .A2(G868), .ZN(new_n645));
  INV_X1    g220(.A(G299), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(G868), .ZN(G297));
  OAI21_X1  g222(.A(new_n645), .B1(new_n646), .B2(G868), .ZN(G280));
  INV_X1    g223(.A(new_n640), .ZN(new_n649));
  INV_X1    g224(.A(G559), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n649), .B1(new_n650), .B2(G860), .ZN(G148));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G868), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n579), .B2(G868), .ZN(G323));
  XNOR2_X1  g229(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g230(.A1(new_n486), .A2(G135), .ZN(new_n656));
  INV_X1    g231(.A(G123), .ZN(new_n657));
  NOR2_X1   g232(.A1(G99), .A2(G2105), .ZN(new_n658));
  OAI21_X1  g233(.A(G2104), .B1(new_n477), .B2(G111), .ZN(new_n659));
  OAI221_X1 g234(.A(new_n656), .B1(new_n483), .B2(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(G2096), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT13), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT85), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(new_n666), .ZN(G156));
  XNOR2_X1  g242(.A(KEYINPUT15), .B(G2430), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2435), .ZN(new_n669));
  XOR2_X1   g244(.A(G2427), .B(G2438), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT14), .ZN(new_n672));
  XOR2_X1   g247(.A(G2451), .B(G2454), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT16), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1341), .B(G1348), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2443), .B(G2446), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G14), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT86), .Z(G401));
  XOR2_X1   g256(.A(G2072), .B(G2078), .Z(new_n682));
  XOR2_X1   g257(.A(G2067), .B(G2678), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n682), .B1(new_n686), .B2(KEYINPUT18), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G2096), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2100), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n686), .A2(KEYINPUT17), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n684), .A2(new_n685), .ZN(new_n691));
  AOI21_X1  g266(.A(KEYINPUT18), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n689), .B(new_n692), .Z(G227));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT87), .Z(new_n697));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT19), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT88), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT20), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n694), .A2(new_n695), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(new_n699), .A3(new_n696), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n702), .B(new_n705), .C1(new_n699), .C2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT22), .B(G1981), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G24), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n629), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT89), .B(G29), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n484), .A2(G119), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n486), .A2(G131), .ZN(new_n722));
  OR2_X1    g297(.A1(G95), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G107), .C2(new_n477), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n720), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT35), .B(G1991), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n727), .B(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n731));
  INV_X1    g306(.A(G22), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G16), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n714), .A2(KEYINPUT90), .A3(G22), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n733), .B(new_n734), .C1(G166), .C2(new_n714), .ZN(new_n735));
  INV_X1    g310(.A(G1971), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G23), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n613), .A2(new_n617), .A3(new_n618), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT33), .B(G1976), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n714), .A2(G6), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n620), .B1(new_n622), .B2(new_n615), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n621), .A2(new_n503), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n743), .B1(new_n746), .B2(new_n714), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT32), .B(G1981), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n737), .A2(new_n742), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT34), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n718), .B(new_n730), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n754), .B(new_n755), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n714), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n649), .B2(new_n714), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT92), .B(G1348), .Z(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n714), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n714), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(G1966), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT97), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n714), .A2(G5), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G171), .B2(new_n714), .ZN(new_n767));
  INV_X1    g342(.A(G1961), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n473), .A2(new_n479), .A3(new_n481), .ZN(new_n770));
  INV_X1    g345(.A(G29), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT94), .B(G34), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT24), .ZN(new_n773));
  OAI22_X1  g348(.A1(new_n770), .A2(new_n771), .B1(new_n719), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2084), .ZN(new_n775));
  OR2_X1    g350(.A1(G29), .A2(G33), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT25), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n486), .A2(G139), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n477), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n776), .B1(new_n781), .B2(new_n771), .ZN(new_n782));
  INV_X1    g357(.A(G2072), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n769), .A2(new_n775), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n763), .A2(G1966), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n477), .A2(G105), .A3(G2104), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT95), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G141), .B2(new_n486), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n484), .A2(G129), .ZN(new_n791));
  NAND3_X1  g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT26), .Z(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G32), .B(new_n794), .S(G29), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT27), .B(G1996), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n719), .ZN(new_n798));
  INV_X1    g373(.A(G28), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(KEYINPUT30), .ZN(new_n800));
  AOI21_X1  g375(.A(G29), .B1(new_n799), .B2(KEYINPUT30), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n797), .B1(new_n660), .B2(new_n798), .C1(new_n800), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n795), .A2(new_n796), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n786), .A2(new_n787), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n798), .A2(G27), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G164), .B2(new_n798), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G2078), .Z(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT31), .B(G11), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n765), .A2(new_n805), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT98), .ZN(new_n811));
  NOR2_X1   g386(.A1(G16), .A2(G19), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n579), .B2(G16), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G1341), .Z(new_n814));
  NAND3_X1  g389(.A1(new_n714), .A2(KEYINPUT23), .A3(G20), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT23), .ZN(new_n816));
  INV_X1    g391(.A(G20), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G16), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n815), .B(new_n818), .C1(new_n646), .C2(new_n714), .ZN(new_n819));
  INV_X1    g394(.A(G1956), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n798), .A2(G26), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT93), .Z(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(KEYINPUT28), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n486), .A2(G140), .ZN(new_n825));
  OR2_X1    g400(.A1(G104), .A2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n827));
  INV_X1    g402(.A(G128), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n825), .B(new_n827), .C1(new_n828), .C2(new_n483), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G29), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n823), .A2(KEYINPUT28), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n824), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G2067), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n814), .A2(new_n821), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n810), .B2(KEYINPUT98), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n756), .A2(new_n761), .A3(new_n811), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n798), .A2(G35), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G162), .B2(new_n798), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT29), .Z(new_n840));
  INV_X1    g415(.A(G2090), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT99), .Z(new_n843));
  NOR2_X1   g418(.A1(new_n840), .A2(new_n841), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n837), .A2(new_n843), .A3(new_n844), .ZN(G311));
  INV_X1    g420(.A(G311), .ZN(G150));
  AOI22_X1  g421(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n503), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  INV_X1    g424(.A(G93), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n615), .A2(new_n849), .B1(new_n551), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NOR2_X1   g430(.A1(new_n567), .A2(KEYINPUT78), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n577), .B1(new_n572), .B2(new_n576), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n567), .A2(new_n852), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT39), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n649), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n861), .B(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n855), .B1(new_n864), .B2(G860), .ZN(G145));
  XNOR2_X1  g440(.A(new_n794), .B(new_n726), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n496), .A2(new_n501), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n781), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n866), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n770), .B(new_n490), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n486), .A2(G142), .ZN(new_n871));
  INV_X1    g446(.A(G130), .ZN(new_n872));
  NOR2_X1   g447(.A1(G106), .A2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(new_n477), .B2(G118), .ZN(new_n874));
  OAI221_X1 g449(.A(new_n871), .B1(new_n483), .B2(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n660), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n870), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n869), .B(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n829), .B(new_n663), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(KEYINPUT100), .B(G37), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g458(.A1(new_n853), .A2(new_n641), .ZN(new_n884));
  NAND2_X1  g459(.A1(G299), .A2(new_n640), .ZN(new_n885));
  INV_X1    g460(.A(new_n604), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n592), .B2(new_n597), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(new_n603), .A3(new_n649), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n649), .B1(new_n887), .B2(new_n603), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n590), .A2(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n892));
  NOR4_X1   g467(.A1(new_n892), .A2(new_n640), .A3(new_n602), .A4(new_n886), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n888), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n652), .B(KEYINPUT101), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n860), .B(new_n897), .ZN(new_n898));
  MUX2_X1   g473(.A(new_n889), .B(new_n896), .S(new_n898), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n746), .A2(G288), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n739), .A2(G305), .ZN(new_n901));
  NAND3_X1  g476(.A1(G166), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(G166), .B1(new_n900), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g479(.A(G290), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n901), .ZN(new_n906));
  INV_X1    g481(.A(G166), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n629), .A3(new_n902), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT42), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n899), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n884), .B1(new_n912), .B2(new_n641), .ZN(G295));
  OAI21_X1  g488(.A(new_n884), .B1(new_n912), .B2(new_n641), .ZN(G331));
  AND2_X1   g489(.A1(new_n905), .A2(new_n909), .ZN(new_n915));
  OAI21_X1  g490(.A(G171), .B1(new_n543), .B2(new_n544), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n541), .A2(new_n542), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n541), .A2(new_n542), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(G301), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n858), .A2(new_n920), .A3(new_n859), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n919), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n852), .B1(new_n568), .B2(new_n578), .ZN(new_n923));
  INV_X1    g498(.A(new_n859), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n896), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n921), .A2(new_n925), .B1(new_n885), .B2(new_n888), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n915), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n921), .A2(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n889), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n896), .A2(new_n921), .A3(new_n925), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n910), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n881), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT104), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n928), .A2(new_n932), .A3(new_n935), .A4(new_n881), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(KEYINPUT43), .A3(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n928), .A2(new_n932), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(KEYINPUT44), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n937), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n939), .B1(new_n938), .B2(new_n940), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT103), .B1(new_n933), .B2(KEYINPUT43), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n946), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n946), .A2(KEYINPUT106), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(G397));
  XNOR2_X1  g533(.A(new_n829), .B(new_n833), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT108), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n867), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G160), .A2(G40), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n969));
  INV_X1    g544(.A(new_n966), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n794), .B(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n968), .B(new_n969), .C1(new_n970), .C2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT110), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n725), .B(new_n729), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n975), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n966), .B1(KEYINPUT111), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n974), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n629), .A2(new_n717), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n970), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT48), .Z(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n974), .A2(new_n729), .A3(new_n726), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(G2067), .B2(new_n829), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n966), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n970), .B2(G1996), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n966), .B1(new_n960), .B2(new_n794), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n966), .A2(KEYINPUT46), .A3(new_n971), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n995));
  XNOR2_X1  g570(.A(new_n994), .B(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n986), .A2(new_n989), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n983), .A2(KEYINPUT107), .ZN(new_n998));
  NAND2_X1  g573(.A1(G290), .A2(G1986), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n980), .B1(new_n966), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G40), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n770), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n867), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n964), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n736), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n867), .A2(new_n961), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(new_n1003), .A3(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(G2090), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1005), .A2(KEYINPUT112), .A3(new_n736), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1008), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1016), .A2(G8), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n1018));
  NAND4_X1  g593(.A1(G303), .A2(new_n1018), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT55), .B(G8), .C1(new_n608), .C2(new_n609), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT114), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n608), .A2(new_n609), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1017), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT115), .B(G1981), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n746), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(G305), .A2(KEYINPUT116), .A3(G1981), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT116), .B1(G305), .B2(G1981), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n965), .A2(new_n962), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(new_n1024), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT49), .B(new_n1029), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1037), .B1(new_n1040), .B2(G288), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1037), .B(new_n1043), .C1(new_n1040), .C2(G288), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1027), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1039), .A2(new_n1040), .A3(new_n739), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1029), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1046), .B1(new_n1037), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n962), .A2(new_n1010), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n1003), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1011), .B1(new_n867), .B2(new_n961), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n965), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1051), .B(new_n1054), .C1(KEYINPUT50), .C2(new_n962), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1006), .B1(new_n1055), .B2(G2090), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G8), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1057), .A2(new_n1025), .A3(new_n1021), .A4(new_n1019), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1045), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1027), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1966), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1005), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2084), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1009), .A2(new_n1063), .A3(new_n1003), .A4(new_n1012), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(G168), .A3(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G286), .A2(KEYINPUT123), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT123), .B1(new_n1065), .B2(G8), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT51), .B1(new_n1071), .B2(KEYINPUT122), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT62), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  OR3_X1    g650(.A1(new_n1005), .A2(new_n1075), .A3(G2078), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1013), .A2(new_n768), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1075), .B1(new_n1005), .B2(G2078), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1079), .A2(G171), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1070), .A2(new_n1072), .A3(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1060), .A2(new_n1074), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1055), .A2(new_n820), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT56), .B(G2072), .Z(new_n1085));
  OR2_X1    g660(.A1(new_n1005), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n598), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(G299), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1087), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1013), .A2(new_n760), .B1(new_n1036), .B2(new_n833), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n649), .A2(KEYINPUT60), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n649), .A2(KEYINPUT60), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n964), .A2(new_n971), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1099), .A2(KEYINPUT121), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n965), .B2(new_n962), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(KEYINPUT121), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n579), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1104), .B2(new_n579), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1093), .B(new_n1098), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1098), .B(new_n1088), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1094), .A2(new_n640), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1109), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1045), .B1(new_n1017), .B2(new_n1026), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1117), .A2(new_n1073), .A3(new_n1058), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1079), .A2(G301), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1076), .A2(G171), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(KEYINPUT124), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1119), .A2(KEYINPUT124), .A3(KEYINPUT54), .A4(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1118), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1049), .B(new_n1083), .C1(new_n1116), .C2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(G8), .A3(G168), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT118), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1128), .A2(new_n1131), .A3(G8), .A4(G168), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1027), .A2(new_n1058), .A3(new_n1059), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1135), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1026), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1016), .A2(G8), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1142), .A2(new_n1117), .A3(new_n1133), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1138), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(KEYINPUT125), .B(new_n1001), .C1(new_n1127), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT119), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1142), .A2(new_n1117), .A3(new_n1133), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(new_n1137), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1114), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1118), .B(new_n1125), .C1(new_n1151), .C2(new_n1109), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1150), .A2(new_n1049), .A3(new_n1152), .A4(new_n1083), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT125), .B1(new_n1153), .B2(new_n1001), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n997), .B1(new_n1146), .B2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g730(.A(G227), .ZN(new_n1157));
  AND4_X1   g731(.A1(G319), .A2(new_n882), .A3(new_n680), .A4(new_n1157), .ZN(new_n1158));
  AND4_X1   g732(.A1(new_n712), .A2(new_n949), .A3(new_n951), .A4(new_n1158), .ZN(G308));
  NAND4_X1  g733(.A1(new_n712), .A2(new_n949), .A3(new_n951), .A4(new_n1158), .ZN(G225));
endmodule


