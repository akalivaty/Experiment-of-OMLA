//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1296, new_n1297, new_n1298, new_n1299;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT65), .Z(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n459), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n462), .A2(new_n470), .ZN(G160));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT66), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n459), .A2(new_n476), .A3(G2105), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT67), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT68), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n465), .A2(G136), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g060(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(G162));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n461), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n474), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n461), .C1(new_n472), .C2(new_n473), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n465), .A2(new_n493), .A3(G138), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT69), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .A3(G543), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n498), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT70), .B(G88), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(G50), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n507), .B1(new_n498), .B2(new_n500), .ZN(new_n508));
  AND2_X1   g083(.A1(G75), .A2(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(G651), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n506), .A2(KEYINPUT71), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT71), .B1(new_n506), .B2(new_n510), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n516), .A2(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(KEYINPUT7), .ZN(new_n518));
  AOI22_X1  g093(.A1(G51), .A2(new_n505), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n503), .A2(G89), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n499), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT5), .B1(new_n499), .B2(G543), .ZN(new_n522));
  OAI211_X1 g097(.A(G63), .B(G651), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n519), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(G168));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n498), .A2(new_n500), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G64), .ZN(new_n528));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT6), .B(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n527), .A2(G90), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n505), .A2(G52), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(new_n527), .A2(G56), .ZN(new_n536));
  NAND2_X1  g111(.A1(G68), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n526), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n527), .A2(G81), .A3(new_n531), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n505), .A2(G43), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT73), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n550));
  INV_X1    g125(.A(G65), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n498), .B2(new_n500), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(KEYINPUT6), .A2(G651), .ZN(new_n556));
  NOR2_X1   g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n503), .A2(G91), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n555), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n559), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n531), .A2(KEYINPUT74), .A3(G53), .A4(G543), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT9), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n550), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n555), .A2(new_n561), .A3(new_n562), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT9), .ZN(new_n569));
  NOR3_X1   g144(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT75), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n517), .A2(new_n518), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n531), .A2(G51), .A3(G543), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n523), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n527), .A2(G89), .A3(new_n531), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT76), .A4(new_n523), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G286));
  NAND2_X1  g156(.A1(new_n503), .A2(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n505), .A2(G49), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  AOI22_X1  g160(.A1(new_n503), .A2(G86), .B1(new_n505), .B2(G48), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n498), .B2(new_n500), .ZN(new_n588));
  AND2_X1   g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n503), .A2(G85), .B1(new_n505), .B2(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n526), .B2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n505), .A2(G54), .ZN(new_n596));
  AND2_X1   g171(.A1(G79), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n527), .B2(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n596), .B1(new_n598), .B2(new_n526), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n503), .A2(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n503), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n595), .B1(G868), .B2(new_n604), .ZN(G284));
  OAI21_X1  g180(.A(new_n595), .B1(G868), .B2(new_n604), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(G286), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n607), .ZN(G297));
  AOI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n607), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n604), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n604), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n478), .A2(G123), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n465), .A2(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n461), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2096), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XOR2_X1   g200(.A(KEYINPUT77), .B(KEYINPUT13), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(G2096), .ZN(new_n631));
  NAND4_X1  g206(.A1(new_n623), .A2(new_n629), .A3(new_n630), .A4(new_n631), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(G14), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT78), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT17), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n653), .B1(new_n650), .B2(new_n652), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n651), .B2(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(new_n652), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n657), .A2(new_n653), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  OR3_X1    g235(.A1(new_n654), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n661), .A2(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT79), .B(G2096), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(G2100), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n663), .B1(new_n662), .B2(new_n664), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT80), .ZN(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n678), .C1(new_n669), .C2(new_n677), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT81), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n684), .A2(new_n687), .A3(new_n685), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(G305), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G16), .ZN(new_n694));
  OR2_X1    g269(.A1(G6), .A2(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(KEYINPUT32), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT32), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n694), .A2(new_n698), .A3(new_n695), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G1981), .ZN(new_n701));
  INV_X1    g276(.A(G1981), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n697), .A2(new_n702), .A3(new_n699), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(G303), .A2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G22), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT83), .Z(new_n710));
  NAND3_X1  g285(.A1(new_n706), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n707), .B1(new_n706), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n708), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT33), .B(G1976), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n704), .A2(new_n705), .A3(new_n711), .A4(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G25), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n477), .A3(G119), .ZN(new_n722));
  INV_X1    g297(.A(G95), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n723), .A2(new_n461), .A3(KEYINPUT82), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT82), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G95), .B2(G2105), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G107), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n467), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  AOI22_X1  g304(.A1(G131), .A2(new_n465), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n721), .B1(new_n732), .B2(new_n720), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  XOR2_X1   g309(.A(new_n733), .B(new_n734), .Z(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G24), .ZN(new_n736));
  INV_X1    g311(.A(G290), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G16), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1986), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n719), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n718), .A2(new_n711), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n705), .B1(new_n743), .B2(new_n704), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT36), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n704), .ZN(new_n746));
  OAI21_X1  g321(.A(KEYINPUT34), .B1(new_n746), .B2(new_n742), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n747), .A2(new_n748), .A3(new_n719), .A4(new_n740), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(new_n461), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT86), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n465), .A2(G139), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(KEYINPUT85), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT85), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n465), .A2(new_n757), .A3(G139), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n752), .B2(new_n753), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n720), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n720), .B2(G33), .ZN(new_n766));
  INV_X1    g341(.A(G2072), .ZN(new_n767));
  INV_X1    g342(.A(G1348), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n604), .A2(G16), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G4), .B2(G16), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n768), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n771), .B(new_n772), .C1(new_n767), .C2(new_n766), .ZN(new_n773));
  NOR2_X1   g348(.A1(G27), .A2(G29), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G164), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT90), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2078), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n475), .A2(new_n477), .A3(G129), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT26), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g359(.A(G141), .B(new_n461), .C1(new_n472), .C2(new_n473), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n468), .A2(G105), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n779), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(KEYINPUT87), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n779), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n793), .A2(KEYINPUT88), .A3(G29), .ZN(new_n794));
  INV_X1    g369(.A(G32), .ZN(new_n795));
  AOI21_X1  g370(.A(KEYINPUT88), .B1(new_n720), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n792), .B2(new_n720), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT27), .B(G1996), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n708), .A2(G20), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT23), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n609), .B2(new_n708), .ZN(new_n803));
  INV_X1    g378(.A(G1956), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n778), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n720), .A2(G35), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G162), .B2(new_n720), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT29), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT29), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(new_n807), .C1(G162), .C2(new_n720), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G2090), .ZN(new_n813));
  NOR2_X1   g388(.A1(G168), .A2(new_n708), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n708), .B2(G21), .ZN(new_n815));
  INV_X1    g390(.A(G1966), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT89), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n720), .A2(G26), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT28), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT84), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n465), .A2(new_n821), .A3(G140), .ZN(new_n822));
  OAI211_X1 g397(.A(G140), .B(new_n461), .C1(new_n472), .C2(new_n473), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT84), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n475), .A2(new_n477), .A3(G128), .ZN(new_n826));
  OR2_X1    g401(.A1(G104), .A2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n827), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n820), .B1(new_n829), .B2(new_n720), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G2067), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n818), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G2090), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n809), .A2(new_n833), .A3(new_n811), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n542), .A2(G16), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G16), .B2(G19), .ZN(new_n836));
  INV_X1    g411(.A(G1341), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(G171), .A2(G16), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G5), .B2(G16), .ZN(new_n840));
  INV_X1    g415(.A(G1961), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n837), .B2(new_n836), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT24), .ZN(new_n844));
  INV_X1    g419(.A(G34), .ZN(new_n845));
  AOI21_X1  g420(.A(G29), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G160), .B2(new_n720), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(G2084), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT31), .B(G11), .Z(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT30), .B(G28), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n720), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n622), .B2(new_n720), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n848), .A2(G2084), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n849), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n815), .A2(new_n816), .B1(new_n840), .B2(new_n841), .ZN(new_n856));
  AND4_X1   g431(.A1(new_n838), .A2(new_n843), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n813), .A2(new_n832), .A3(new_n834), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n806), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n750), .A2(new_n859), .ZN(G311));
  AND3_X1   g435(.A1(new_n750), .A2(new_n859), .A3(KEYINPUT91), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT91), .B1(new_n750), .B2(new_n859), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(G150));
  NAND2_X1  g438(.A1(new_n505), .A2(G55), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n527), .A2(G93), .A3(new_n531), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n526), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n604), .A2(G559), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n527), .A2(G67), .ZN(new_n872));
  NAND2_X1  g447(.A1(G80), .A2(G543), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n526), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n865), .A2(new_n864), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n540), .B(new_n539), .C1(new_n877), .C2(new_n526), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT92), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT92), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n542), .A2(new_n880), .A3(new_n867), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT93), .B1(new_n542), .B2(new_n867), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT93), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n876), .A2(new_n884), .A3(new_n878), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n871), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n888), .A2(KEYINPUT39), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT94), .Z(new_n890));
  INV_X1    g465(.A(KEYINPUT95), .ZN(new_n891));
  AOI21_X1  g466(.A(G860), .B1(new_n888), .B2(KEYINPUT39), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n869), .B1(new_n893), .B2(new_n894), .ZN(G145));
  XNOR2_X1  g470(.A(KEYINPUT101), .B(G37), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n475), .A2(new_n477), .A3(G130), .ZN(new_n900));
  OAI21_X1  g475(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n901));
  INV_X1    g476(.A(G118), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(G2105), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(G142), .B2(new_n465), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n904), .A3(new_n625), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n625), .B1(new_n900), .B2(new_n904), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n906), .A2(new_n732), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n900), .A2(new_n904), .ZN(new_n909));
  INV_X1    g484(.A(new_n625), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n731), .B1(new_n911), .B2(new_n905), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n899), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n732), .B1(new_n906), .B2(new_n907), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n731), .A3(new_n905), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n898), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n913), .A2(KEYINPUT100), .A3(new_n916), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n789), .A2(new_n829), .A3(new_n791), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n779), .A2(new_n787), .A3(new_n790), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n790), .B1(new_n779), .B2(new_n787), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n494), .A2(new_n492), .ZN(new_n926));
  INV_X1    g501(.A(new_n490), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT96), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G164), .A2(KEYINPUT96), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n921), .A2(new_n925), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n921), .B2(new_n925), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT97), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n760), .A2(new_n764), .A3(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n754), .A2(new_n759), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT97), .B1(new_n938), .B2(new_n763), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n921), .A2(new_n925), .ZN(new_n941));
  INV_X1    g516(.A(new_n932), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n921), .A2(new_n925), .A3(new_n932), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n919), .B(new_n920), .C1(new_n937), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n936), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n947), .A3(new_n944), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n936), .A2(new_n939), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n933), .B2(new_n934), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n913), .A2(KEYINPUT100), .A3(new_n916), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT100), .B1(new_n913), .B2(new_n916), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n948), .B(new_n950), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n946), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n622), .B(G160), .ZN(new_n955));
  XNOR2_X1  g530(.A(G162), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n897), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n950), .A2(new_n948), .A3(new_n917), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT102), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n950), .A2(new_n948), .A3(new_n960), .A4(new_n917), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n951), .A2(new_n952), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n950), .A2(new_n948), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n956), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n957), .A2(KEYINPUT103), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT103), .B1(new_n957), .B2(new_n966), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT40), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n957), .A2(new_n966), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT40), .B1(new_n974), .B2(new_n967), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n971), .A2(new_n975), .ZN(G395));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n614), .B(new_n977), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n879), .A2(new_n881), .B1(new_n883), .B2(new_n885), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n614), .B(KEYINPUT104), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n887), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT41), .ZN(new_n984));
  OAI21_X1  g559(.A(G65), .B1(new_n521), .B2(new_n522), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n553), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n986), .A2(G651), .B1(G91), .B2(new_n503), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(new_n550), .A3(new_n566), .A4(new_n561), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT75), .B1(new_n568), .B2(new_n569), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n988), .A2(new_n989), .A3(new_n604), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n604), .B1(new_n988), .B2(new_n989), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n984), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n602), .A2(new_n603), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n993), .B(new_n596), .C1(new_n526), .C2(new_n598), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n567), .B2(new_n570), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n989), .A3(new_n604), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(KEYINPUT41), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT105), .B1(new_n983), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n996), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n983), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n980), .A2(new_n982), .A3(new_n998), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT42), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1000), .A2(new_n1007), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n512), .A2(new_n513), .A3(new_n714), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n506), .A2(new_n510), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT71), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(G288), .B1(new_n1013), .B2(new_n511), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n693), .A2(G290), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n737), .A2(G305), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1010), .A2(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1016), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1019), .A2(new_n1009), .A3(new_n1014), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1006), .A2(new_n1008), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1023));
  OAI21_X1  g598(.A(G868), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n867), .A2(new_n607), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(G295));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1025), .ZN(G331));
  INV_X1    g602(.A(KEYINPUT106), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n578), .A2(G171), .A3(new_n1028), .A4(new_n579), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n578), .A2(G171), .A3(new_n579), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT106), .B1(G171), .B2(new_n524), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n979), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n979), .A2(new_n1032), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n990), .A2(new_n991), .A3(new_n984), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT41), .B1(new_n995), .B2(new_n996), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n1033), .A2(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G301), .A2(G168), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(KEYINPUT106), .C1(G301), .C2(new_n580), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n887), .A2(new_n1039), .A3(new_n1029), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n979), .A2(new_n1032), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1001), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1021), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1021), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1040), .A2(new_n1001), .A3(new_n1041), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1040), .A2(new_n1041), .B1(new_n992), .B2(new_n997), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G37), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1044), .B1(new_n1050), .B2(KEYINPUT107), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT43), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT107), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1048), .A2(new_n1053), .A3(new_n1049), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1051), .A2(KEYINPUT108), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1021), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT107), .B1(new_n1056), .B2(G37), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1057), .A2(new_n1054), .A3(new_n1052), .A4(new_n1043), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1048), .A2(new_n896), .A3(new_n1043), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT109), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1048), .A2(new_n1043), .A3(new_n1063), .A4(new_n896), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(KEYINPUT43), .A3(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1055), .A2(new_n1060), .A3(KEYINPUT44), .A4(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1057), .A2(new_n1054), .A3(KEYINPUT43), .A4(new_n1043), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT44), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1061), .A2(new_n1052), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1070), .ZN(G397));
  OR2_X1    g646(.A1(new_n792), .A2(G1996), .ZN(new_n1072));
  INV_X1    g647(.A(G2067), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n922), .B(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n792), .A2(G1996), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  XOR2_X1   g651(.A(new_n731), .B(new_n734), .Z(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1384), .B1(new_n926), .B2(new_n927), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT110), .B1(G164), .B2(G1384), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT45), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n472), .A2(new_n473), .ZN(new_n1085));
  INV_X1    g660(.A(G125), .ZN(new_n1086));
  INV_X1    g661(.A(G113), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1085), .A2(new_n1086), .B1(new_n1087), .B2(new_n467), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G2105), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(G40), .A3(new_n469), .A4(new_n466), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1078), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1986), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1094), .A3(new_n737), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(KEYINPUT48), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(KEYINPUT48), .B2(new_n1096), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n732), .A2(new_n734), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1076), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1073), .B2(new_n829), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(new_n1092), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1092), .A2(G1996), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(KEYINPUT46), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1074), .A2(new_n793), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1091), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(KEYINPUT46), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(KEYINPUT127), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1107), .A2(KEYINPUT127), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(KEYINPUT47), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(KEYINPUT47), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1102), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G8), .ZN(new_n1114));
  INV_X1    g689(.A(G40), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n462), .A2(new_n470), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1116), .B2(new_n1079), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n586), .A2(new_n702), .A3(new_n590), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT113), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n586), .A2(new_n1120), .A3(new_n590), .A4(new_n702), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1119), .A2(new_n1121), .B1(G305), .B2(G1981), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1117), .B1(new_n1122), .B2(KEYINPUT49), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G305), .A2(G1981), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(KEYINPUT49), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1122), .A2(KEYINPUT114), .A3(KEYINPUT49), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1123), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n714), .A2(G1976), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1117), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT52), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT112), .B(G1976), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT52), .B1(G288), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1117), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT115), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1117), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT49), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT114), .B1(new_n1122), .B2(KEYINPUT49), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1137), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1138), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT50), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1079), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1152));
  AND4_X1   g727(.A1(new_n833), .A2(new_n1151), .A3(new_n1152), .A4(new_n1116), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT111), .B(G1971), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1090), .B1(new_n1079), .B2(KEYINPUT45), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1083), .B1(G164), .B2(G1384), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(G8), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1013), .A2(G8), .A3(new_n511), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT55), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1013), .A2(KEYINPUT55), .A3(G8), .A4(new_n511), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1163), .B(G8), .C1(new_n1153), .C2(new_n1157), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(G1384), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n928), .A2(KEYINPUT45), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1156), .A2(new_n1169), .A3(new_n1116), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n816), .ZN(new_n1171));
  INV_X1    g746(.A(G2084), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1151), .A2(new_n1152), .A3(new_n1172), .A4(new_n1116), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1174), .A2(KEYINPUT63), .A3(G8), .A4(new_n580), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1167), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1149), .A2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1178));
  NAND4_X1  g753(.A1(new_n1165), .A2(new_n1145), .A3(new_n1146), .A4(new_n1166), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1174), .A2(G8), .A3(new_n580), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1173), .ZN(new_n1183));
  AOI21_X1  g758(.A(G1966), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1184));
  OAI21_X1  g759(.A(G8), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n524), .A2(G8), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1185), .A2(KEYINPUT51), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT51), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1188), .B(G8), .C1(new_n1174), .C2(new_n524), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT120), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1186), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1174), .B2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g767(.A(KEYINPUT120), .B(new_n1186), .C1(new_n1171), .C2(new_n1173), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1187), .B(new_n1189), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(KEYINPUT62), .ZN(new_n1195));
  INV_X1    g770(.A(G2078), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1156), .A2(new_n1169), .A3(new_n1196), .A4(new_n1116), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT121), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1155), .A2(KEYINPUT121), .A3(new_n1196), .A4(new_n1156), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1199), .A2(KEYINPUT53), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT53), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1151), .A2(new_n1152), .A3(new_n1116), .ZN(new_n1203));
  AOI22_X1  g778(.A1(new_n1202), .A2(new_n1197), .B1(new_n1203), .B2(new_n841), .ZN(new_n1204));
  AOI21_X1  g779(.A(G301), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1179), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1191), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(KEYINPUT120), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1174), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1211), .A2(new_n1212), .A3(new_n1187), .A4(new_n1189), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1195), .A2(new_n1207), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1166), .ZN(new_n1215));
  OR2_X1    g790(.A1(G288), .A2(G1976), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1124), .B1(new_n1130), .B2(new_n1216), .ZN(new_n1217));
  AOI22_X1  g792(.A1(new_n1149), .A2(new_n1215), .B1(new_n1117), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1182), .A2(new_n1214), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1179), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT54), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1197), .A2(new_n1202), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1203), .A2(new_n841), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1222), .A2(new_n1223), .A3(G301), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT123), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1088), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n460), .A2(KEYINPUT123), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1226), .A2(new_n1227), .A3(G2105), .ZN(new_n1228));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n470), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n466), .A2(KEYINPUT122), .A3(new_n469), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n1232));
  OAI211_X1 g807(.A(KEYINPUT53), .B(G40), .C1(new_n1232), .C2(G2078), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1233), .B1(new_n1232), .B2(G2078), .ZN(new_n1234));
  NAND4_X1  g809(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .A4(new_n1234), .ZN(new_n1235));
  NOR3_X1   g810(.A1(G164), .A2(new_n1083), .A3(G1384), .ZN(new_n1236));
  NOR2_X1   g811(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1237), .A2(new_n1084), .ZN(new_n1238));
  INV_X1    g813(.A(KEYINPUT125), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1237), .A2(new_n1084), .A3(KEYINPUT125), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1224), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1221), .B1(new_n1242), .B2(new_n1205), .ZN(new_n1243));
  NAND3_X1  g818(.A1(new_n1201), .A2(G301), .A3(new_n1204), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1245));
  AOI21_X1  g820(.A(new_n1245), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1246));
  OAI211_X1 g821(.A(KEYINPUT54), .B(new_n1244), .C1(new_n1246), .C2(G301), .ZN(new_n1247));
  NAND4_X1  g822(.A1(new_n1220), .A2(new_n1243), .A3(new_n1247), .A4(new_n1194), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1116), .A2(new_n1079), .ZN(new_n1249));
  NOR2_X1   g824(.A1(new_n1249), .A2(G2067), .ZN(new_n1250));
  AOI21_X1  g825(.A(new_n1250), .B1(new_n768), .B2(new_n1203), .ZN(new_n1251));
  INV_X1    g826(.A(KEYINPUT60), .ZN(new_n1252));
  NAND3_X1  g827(.A1(new_n1251), .A2(new_n1252), .A3(new_n604), .ZN(new_n1253));
  XOR2_X1   g828(.A(KEYINPUT58), .B(G1341), .Z(new_n1254));
  NAND2_X1  g829(.A1(new_n1249), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g830(.A(new_n1255), .B1(new_n1170), .B2(G1996), .ZN(new_n1256));
  AND2_X1   g831(.A1(new_n1256), .A2(new_n542), .ZN(new_n1257));
  OAI21_X1  g832(.A(new_n1253), .B1(new_n1257), .B2(KEYINPUT59), .ZN(new_n1258));
  AND3_X1   g833(.A1(new_n1256), .A2(KEYINPUT59), .A3(new_n542), .ZN(new_n1259));
  NOR2_X1   g834(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AND2_X1   g835(.A1(new_n1251), .A2(new_n994), .ZN(new_n1261));
  NOR2_X1   g836(.A1(new_n1251), .A2(new_n994), .ZN(new_n1262));
  OAI21_X1  g837(.A(KEYINPUT60), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g838(.A1(new_n563), .A2(new_n566), .ZN(new_n1264));
  NOR2_X1   g839(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1265));
  NAND2_X1  g840(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1266));
  XOR2_X1   g841(.A(new_n1266), .B(KEYINPUT118), .Z(new_n1267));
  INV_X1    g842(.A(new_n1267), .ZN(new_n1268));
  OR3_X1    g843(.A1(new_n1264), .A2(new_n1265), .A3(new_n1268), .ZN(new_n1269));
  OAI21_X1  g844(.A(new_n1268), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1270));
  NAND2_X1  g845(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g846(.A1(new_n1271), .A2(KEYINPUT119), .ZN(new_n1272));
  INV_X1    g847(.A(KEYINPUT119), .ZN(new_n1273));
  NAND3_X1  g848(.A1(new_n1269), .A2(new_n1270), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g849(.A1(new_n1203), .A2(new_n804), .ZN(new_n1275));
  XNOR2_X1  g850(.A(KEYINPUT56), .B(G2072), .ZN(new_n1276));
  NAND3_X1  g851(.A1(new_n1155), .A2(new_n1156), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g852(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g853(.A1(new_n1272), .A2(new_n1274), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g854(.A1(new_n1271), .A2(new_n1275), .A3(new_n1277), .ZN(new_n1280));
  NAND3_X1  g855(.A1(new_n1279), .A2(KEYINPUT61), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g856(.A(KEYINPUT61), .ZN(new_n1282));
  INV_X1    g857(.A(new_n1280), .ZN(new_n1283));
  AOI21_X1  g858(.A(new_n1271), .B1(new_n1277), .B2(new_n1275), .ZN(new_n1284));
  OAI21_X1  g859(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND4_X1  g860(.A1(new_n1260), .A2(new_n1263), .A3(new_n1281), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g861(.A1(new_n1262), .A2(new_n1280), .ZN(new_n1287));
  AND2_X1   g862(.A1(new_n1287), .A2(new_n1279), .ZN(new_n1288));
  AOI22_X1  g863(.A1(new_n1248), .A2(KEYINPUT126), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  OR2_X1    g864(.A1(new_n1248), .A2(KEYINPUT126), .ZN(new_n1290));
  AOI21_X1  g865(.A(new_n1219), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  XOR2_X1   g866(.A(G290), .B(G1986), .Z(new_n1292));
  AOI21_X1  g867(.A(new_n1092), .B1(new_n1078), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g868(.A(new_n1113), .B1(new_n1291), .B2(new_n1293), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g869(.A1(new_n974), .A2(new_n967), .ZN(new_n1296));
  AND2_X1   g870(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1297));
  OAI211_X1 g871(.A(G319), .B(new_n647), .C1(new_n665), .C2(new_n666), .ZN(new_n1298));
  AOI21_X1  g872(.A(new_n1298), .B1(new_n689), .B2(new_n690), .ZN(new_n1299));
  AND3_X1   g873(.A1(new_n1296), .A2(new_n1297), .A3(new_n1299), .ZN(G308));
  NAND3_X1  g874(.A1(new_n1296), .A2(new_n1297), .A3(new_n1299), .ZN(G225));
endmodule


