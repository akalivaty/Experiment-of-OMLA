//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  OR4_X1    g026(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n452));
  OR2_X1    g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  XNOR2_X1  g031(.A(KEYINPUT3), .B(G2104), .ZN(new_n457));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n457), .A2(G137), .A3(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT68), .B1(new_n460), .B2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(new_n458), .A3(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT67), .A4(G125), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n474), .B2(G2105), .ZN(G160));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n466), .A2(new_n468), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n458), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n466), .A2(new_n468), .A3(new_n458), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n478), .A2(KEYINPUT69), .A3(G124), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n481), .A2(new_n483), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n466), .A2(new_n468), .A3(G126), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n460), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G102), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n458), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n457), .A2(KEYINPUT4), .A3(G138), .A4(new_n458), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n492), .A2(new_n494), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT71), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(G62), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT70), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .A3(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n505), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n501), .B1(new_n516), .B2(new_n518), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n519), .A2(G88), .B1(new_n520), .B2(G50), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n513), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT72), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT72), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n524), .A2(KEYINPUT7), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT7), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(new_n520), .A2(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n516), .A2(new_n518), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(G90), .A3(new_n509), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n537), .B1(new_n534), .B2(new_n536), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n505), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n542), .A2(new_n543), .A3(G651), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n543), .B1(new_n542), .B2(G651), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n538), .A2(new_n539), .B1(new_n544), .B2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  AOI22_X1  g122(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n515), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(G43), .B2(new_n520), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n519), .A2(G81), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(new_n554));
  XOR2_X1   g129(.A(new_n554), .B(KEYINPUT75), .Z(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n520), .A2(new_n561), .A3(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n520), .A2(new_n561), .A3(new_n564), .A4(G53), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(KEYINPUT77), .B(G65), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n509), .A2(new_n567), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n515), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n519), .A2(G91), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(G299));
  NAND2_X1  g146(.A1(new_n513), .A2(new_n521), .ZN(G303));
  NAND2_X1  g147(.A1(new_n519), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n520), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n505), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(G48), .B2(new_n520), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n519), .A2(G86), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n505), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G47), .B2(new_n520), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n519), .A2(G85), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(KEYINPUT79), .B(G66), .Z(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n505), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n520), .B2(G54), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n594));
  NAND3_X1  g169(.A1(new_n519), .A2(G92), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n535), .A2(new_n509), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n593), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT80), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n589), .B1(new_n601), .B2(G868), .ZN(G284));
  XOR2_X1   g177(.A(G284), .B(KEYINPUT81), .Z(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G91), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n568), .A2(new_n515), .B1(new_n597), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n565), .B2(new_n563), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n604), .B1(G868), .B2(new_n607), .ZN(G297));
  OAI21_X1  g183(.A(new_n604), .B1(G868), .B2(new_n607), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n601), .B1(new_n610), .B2(G860), .ZN(G148));
  OR2_X1    g186(.A1(new_n553), .A2(G868), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n601), .A2(new_n610), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n478), .A2(G123), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n482), .A2(G135), .ZN(new_n618));
  NOR2_X1   g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(new_n458), .B2(G111), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT83), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n457), .A2(new_n461), .A3(new_n463), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n624), .B(new_n625), .Z(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT13), .B(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2451), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n634), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G14), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT85), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT87), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT17), .ZN(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n646), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n649), .ZN(new_n655));
  INV_X1    g230(.A(new_n651), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n656), .A2(new_n652), .A3(new_n646), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n649), .A2(new_n653), .A3(new_n646), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(G2096), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT88), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  AOI22_X1  g248(.A1(new_n671), .A2(new_n672), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(new_n672), .C2(new_n671), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT22), .B(G1981), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n678), .B(new_n679), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(new_n681), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(G229));
  NOR2_X1   g261(.A1(G4), .A2(G16), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n601), .B2(G16), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1348), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G26), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT91), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n478), .A2(G128), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n482), .A2(G140), .ZN(new_n695));
  OR2_X1    g270(.A1(G104), .A2(G2105), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n696), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n693), .B1(new_n699), .B2(new_n690), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G2067), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n702), .A2(KEYINPUT23), .A3(G20), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT23), .ZN(new_n704));
  INV_X1    g279(.A(G20), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(G16), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n706), .C1(new_n607), .C2(new_n702), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1956), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n689), .A2(new_n701), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n702), .A2(G5), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G171), .B2(new_n702), .ZN(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n622), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n709), .B(new_n713), .C1(new_n690), .C2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G29), .B2(G33), .ZN(new_n717));
  OR3_X1    g292(.A1(new_n716), .A2(G29), .A3(G33), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT94), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT93), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n722), .A2(new_n458), .A3(G103), .A4(G2104), .ZN(new_n723));
  AOI21_X1  g298(.A(KEYINPUT25), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n721), .A2(KEYINPUT25), .A3(new_n723), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n457), .A2(G139), .A3(new_n458), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n457), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n458), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n719), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n726), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(new_n724), .ZN(new_n733));
  NAND2_X1  g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  INV_X1    g309(.A(G127), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n477), .B2(new_n735), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n736), .A2(G2105), .B1(G139), .B2(new_n482), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n733), .A2(new_n737), .A3(KEYINPUT94), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n717), .B(new_n718), .C1(new_n739), .C2(new_n690), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G2072), .Z(new_n741));
  NOR2_X1   g316(.A1(G164), .A2(new_n690), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G27), .B2(new_n690), .ZN(new_n743));
  INV_X1    g318(.A(G2078), .ZN(new_n744));
  NOR2_X1   g319(.A1(G29), .A2(G32), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n478), .A2(G129), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n461), .A2(new_n463), .A3(G105), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n482), .A2(G141), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  NAND4_X1  g325(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n745), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  OAI22_X1  g329(.A1(new_n743), .A2(new_n744), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n741), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n690), .A2(G35), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G162), .B2(new_n690), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT29), .B(G2090), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n743), .A2(new_n744), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n702), .A2(G19), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n553), .B2(new_n702), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1341), .Z(new_n764));
  NAND4_X1  g339(.A1(new_n756), .A2(new_n760), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n753), .A2(new_n754), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT95), .B(G28), .Z(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT30), .Z(new_n768));
  OAI21_X1  g343(.A(new_n766), .B1(G29), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n715), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n702), .A2(G22), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G166), .B2(new_n702), .ZN(new_n774));
  INV_X1    g349(.A(G1971), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G16), .A2(G23), .ZN(new_n777));
  INV_X1    g352(.A(G288), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT33), .B(G1976), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n702), .A2(G6), .ZN(new_n782));
  INV_X1    g357(.A(G305), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n702), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT32), .B(G1981), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n776), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT34), .Z(new_n788));
  AND2_X1   g363(.A1(new_n702), .A2(G24), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G290), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(G1986), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n478), .A2(G119), .B1(new_n482), .B2(G131), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(new_n458), .B2(G107), .ZN(new_n794));
  NOR2_X1   g369(.A1(G95), .A2(G2105), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT89), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n793), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G25), .B(new_n797), .S(G29), .Z(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT35), .B(G1991), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n790), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(G1986), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n788), .A2(new_n792), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT90), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n803), .A2(KEYINPUT90), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n772), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n803), .A2(KEYINPUT90), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n808), .A2(KEYINPUT36), .A3(new_n804), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n771), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n702), .A2(G21), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G168), .B2(new_n702), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1966), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(KEYINPUT24), .A2(G34), .ZN(new_n815));
  NAND2_X1  g390(.A1(KEYINPUT24), .A2(G34), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n815), .A2(new_n690), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G160), .B2(new_n690), .ZN(new_n818));
  INV_X1    g393(.A(G2084), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT31), .B(G11), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n810), .A2(new_n814), .A3(new_n820), .A4(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  AOI22_X1  g398(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(new_n515), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n520), .A2(G55), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n535), .A2(G93), .A3(new_n509), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT96), .ZN(new_n828));
  AOI21_X1  g403(.A(KEYINPUT96), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT97), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(new_n825), .C1(new_n828), .C2(new_n829), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n553), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n553), .A2(new_n830), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT39), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n601), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n838), .B(new_n840), .Z(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT98), .Z(new_n843));
  AND2_X1   g418(.A1(new_n831), .A2(new_n833), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT99), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(new_n487), .B(G160), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n622), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n626), .B(new_n797), .Z(new_n851));
  AND2_X1   g426(.A1(new_n482), .A2(G142), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n478), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(KEYINPUT102), .ZN(new_n855));
  OR2_X1    g430(.A1(G106), .A2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(G2104), .C1(G118), .C2(new_n458), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n851), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n698), .B1(new_n739), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g436(.A(KEYINPUT101), .B(new_n699), .C1(new_n731), .C2(new_n738), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n752), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n727), .A2(new_n730), .A3(new_n719), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT94), .B1(new_n733), .B2(new_n737), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n699), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n739), .A2(new_n860), .A3(new_n698), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n751), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n490), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n457), .B2(G126), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n494), .B1(new_n871), .B2(new_n458), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n497), .A2(new_n498), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT100), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n494), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n491), .B2(G2105), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n876), .A2(new_n877), .A3(new_n497), .A4(new_n498), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n863), .A2(new_n869), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n863), .B2(new_n869), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n859), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT103), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n886), .B(new_n859), .C1(new_n881), .C2(new_n882), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n863), .A2(new_n869), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n879), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n863), .A2(new_n869), .A3(new_n880), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n892), .A2(new_n859), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n885), .B1(new_n884), .B2(new_n887), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n850), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT105), .B(G37), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n850), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n886), .B1(new_n892), .B2(new_n859), .ZN(new_n900));
  INV_X1    g475(.A(new_n887), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n893), .B(new_n899), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n896), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g479(.A1(new_n844), .A2(new_n614), .ZN(new_n905));
  XOR2_X1   g480(.A(G288), .B(KEYINPUT106), .Z(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(G290), .ZN(new_n907));
  XNOR2_X1  g482(.A(G288), .B(KEYINPUT106), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n587), .A3(new_n586), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(G166), .A2(G305), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n783), .A2(G303), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  OR3_X1    g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(new_n911), .B2(new_n912), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n915), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(new_n909), .A3(new_n907), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n919), .B(KEYINPUT42), .Z(new_n920));
  XOR2_X1   g495(.A(new_n837), .B(new_n613), .Z(new_n921));
  XNOR2_X1  g496(.A(G299), .B(new_n600), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(KEYINPUT41), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n921), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n920), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n905), .B1(new_n926), .B2(new_n614), .ZN(G295));
  OAI21_X1  g502(.A(new_n905), .B1(new_n926), .B2(new_n614), .ZN(G331));
  XNOR2_X1  g503(.A(G168), .B(G301), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n834), .B2(new_n836), .ZN(new_n930));
  XNOR2_X1  g505(.A(G301), .B(G286), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(new_n835), .C1(new_n844), .C2(new_n553), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n932), .A3(KEYINPUT108), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n837), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n924), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n922), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n930), .A2(new_n932), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n919), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT109), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n936), .A2(new_n919), .A3(new_n941), .A4(new_n938), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n919), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n922), .B1(new_n933), .B2(new_n935), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n930), .A2(new_n932), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n946), .A2(new_n924), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AND4_X1   g523(.A1(KEYINPUT43), .A2(new_n943), .A3(new_n898), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n940), .B2(new_n942), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n936), .A2(new_n938), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n944), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT43), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT44), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n943), .A2(new_n948), .A3(new_n955), .A4(new_n898), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n955), .B1(new_n950), .B2(new_n952), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n954), .B1(new_n959), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  INV_X1    g536(.A(new_n873), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n877), .B1(new_n962), .B2(new_n876), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT100), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT110), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n879), .A2(new_n968), .A3(new_n961), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n474), .A2(G2105), .ZN(new_n971));
  INV_X1    g546(.A(new_n465), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(G40), .A3(new_n972), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G2067), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n699), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n797), .A2(new_n799), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT125), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n698), .A2(G2067), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n751), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n977), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n975), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(G290), .A2(G1986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n975), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT48), .Z(new_n989));
  AND2_X1   g564(.A1(new_n797), .A2(new_n799), .ZN(new_n990));
  OR3_X1    g565(.A1(new_n984), .A2(new_n990), .A3(new_n978), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n975), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n986), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n974), .A2(G1996), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n994), .A2(KEYINPUT46), .ZN(new_n995));
  INV_X1    g570(.A(new_n981), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n975), .B1(new_n751), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(KEYINPUT46), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT126), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n1000), .A2(KEYINPUT47), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(KEYINPUT47), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n993), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT124), .ZN(new_n1004));
  INV_X1    g579(.A(G8), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n961), .B1(new_n872), .B2(new_n873), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n499), .A2(KEYINPUT50), .A3(new_n961), .ZN(new_n1009));
  AOI211_X1 g584(.A(G2090), .B(new_n973), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n967), .B(G1384), .C1(new_n874), .C2(new_n878), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1006), .A2(new_n967), .ZN(new_n1012));
  INV_X1    g587(.A(G40), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n1013), .B(new_n465), .C1(new_n474), .C2(G2105), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n775), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1010), .B1(new_n1016), .B2(KEYINPUT111), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n879), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n973), .B1(new_n967), .B2(new_n1006), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1971), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1005), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G303), .A2(G8), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n1024), .B(KEYINPUT55), .Z(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1012), .A2(new_n1014), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1966), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1009), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT50), .B1(new_n499), .B2(new_n961), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n819), .B(new_n1014), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1005), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(G168), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n1035), .B2(G168), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1027), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1020), .A2(new_n1010), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1005), .B1(new_n1041), .B2(KEYINPUT114), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(new_n1020), .B2(new_n1010), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1025), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1026), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n973), .A2(new_n1006), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(new_n1005), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(G288), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT52), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G305), .A2(G1981), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n580), .B2(new_n581), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1052), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT112), .ZN(new_n1057));
  OR3_X1    g632(.A1(new_n1053), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n1052), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1057), .A2(new_n1048), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT52), .B1(G288), .B2(new_n1049), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1048), .B(new_n1062), .C1(new_n1049), .C2(G288), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1051), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1046), .A2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(new_n1048), .B(KEYINPUT113), .Z(new_n1067));
  NAND3_X1  g642(.A1(new_n1061), .A2(new_n1049), .A3(new_n778), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1053), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1966), .B1(new_n1019), .B2(new_n1028), .ZN(new_n1071));
  AOI211_X1 g646(.A(G2084), .B(new_n973), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1072));
  OAI211_X1 g647(.A(G8), .B(G168), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT115), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1037), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1075), .B(new_n1065), .C1(new_n1025), .C2(new_n1023), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1070), .B1(new_n1076), .B2(KEYINPUT63), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1066), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(G2078), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1018), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n970), .A2(new_n1014), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1018), .A2(new_n1019), .A3(new_n744), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1014), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1084), .A2(new_n1080), .B1(new_n712), .B2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1083), .A2(G301), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1019), .A2(new_n1028), .A3(new_n1081), .ZN(new_n1088));
  AOI21_X1  g663(.A(G301), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1079), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G171), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1086), .A2(G301), .A3(new_n1088), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(KEYINPUT54), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1025), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1064), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1090), .A2(new_n1094), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(G168), .A2(new_n1005), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1035), .A2(KEYINPUT51), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1100), .B1(new_n1035), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n973), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n819), .A2(new_n1107), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT122), .B1(new_n1108), .B2(new_n1005), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1103), .B(new_n1104), .C1(new_n1106), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1100), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1105), .B(G8), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT123), .B1(new_n1113), .B2(KEYINPUT51), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1102), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1099), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(G299), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT117), .B1(new_n607), .B2(new_n1121), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n607), .A2(KEYINPUT57), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1107), .A2(G1956), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1018), .A2(new_n1019), .A3(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1119), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1018), .A2(new_n1019), .A3(new_n982), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1018), .A2(new_n1019), .A3(KEYINPUT120), .A4(new_n982), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT58), .B(G1341), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1139), .B(new_n1140), .C1(new_n1047), .C2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1142), .A2(KEYINPUT59), .A3(new_n553), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT59), .B1(new_n1142), .B2(new_n553), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1047), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n1107), .A2(G1348), .B1(new_n1146), .B2(G2067), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n600), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1151));
  INV_X1    g726(.A(G1348), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1085), .A2(new_n1152), .B1(new_n976), .B2(new_n1047), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1153), .A2(KEYINPUT121), .A3(KEYINPUT60), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1149), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1149), .B1(new_n1154), .B2(new_n1151), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1126), .B(KEYINPUT118), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1129), .A2(KEYINPUT119), .A3(new_n1131), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT119), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1161), .A2(KEYINPUT61), .A3(new_n1133), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1136), .A2(new_n1145), .A3(new_n1157), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n600), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1133), .A2(new_n1164), .A3(new_n1147), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1165), .A2(new_n1161), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1078), .B1(new_n1118), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1112), .A2(new_n1111), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1035), .A2(new_n1105), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT51), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1103), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1113), .A2(KEYINPUT123), .A3(KEYINPUT51), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1101), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT62), .B1(new_n1174), .B2(new_n1116), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1115), .A2(new_n1176), .A3(new_n1117), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1175), .A2(new_n1089), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1168), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n791), .B1(new_n586), .B2(new_n587), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n991), .A2(new_n987), .A3(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n974), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1004), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1185));
  AOI211_X1 g760(.A(KEYINPUT124), .B(new_n1183), .C1(new_n1168), .C2(new_n1179), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1003), .B1(new_n1185), .B2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n1189));
  XOR2_X1   g763(.A(new_n662), .B(G2100), .Z(new_n1190));
  NAND3_X1  g764(.A1(new_n903), .A2(new_n1190), .A3(new_n644), .ZN(new_n1191));
  AND3_X1   g765(.A1(new_n683), .A2(G319), .A3(new_n685), .ZN(new_n1192));
  OAI21_X1  g766(.A(new_n1192), .B1(new_n957), .B2(new_n958), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1189), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g768(.A(KEYINPUT104), .B1(new_n900), .B2(new_n901), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n1195), .A2(new_n893), .A3(new_n888), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n897), .B1(new_n1196), .B2(new_n850), .ZN(new_n1197));
  AOI21_X1  g771(.A(G227), .B1(new_n1197), .B2(new_n902), .ZN(new_n1198));
  NAND3_X1  g772(.A1(new_n683), .A2(G319), .A3(new_n685), .ZN(new_n1199));
  INV_X1    g773(.A(G37), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n943), .A2(new_n1200), .A3(new_n952), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1201), .A2(KEYINPUT43), .ZN(new_n1202));
  AOI21_X1  g776(.A(new_n1199), .B1(new_n1202), .B2(new_n956), .ZN(new_n1203));
  NAND4_X1  g777(.A1(new_n1198), .A2(new_n1203), .A3(KEYINPUT127), .A4(new_n644), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n1194), .A2(new_n1204), .ZN(G308));
  NAND3_X1  g779(.A1(new_n1198), .A2(new_n1203), .A3(new_n644), .ZN(G225));
endmodule


