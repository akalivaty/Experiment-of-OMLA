

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593;

  XNOR2_X1 U328 ( .A(n381), .B(n380), .ZN(n406) );
  XNOR2_X1 U329 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U330 ( .A(n369), .B(KEYINPUT73), .ZN(n370) );
  XNOR2_X1 U331 ( .A(n427), .B(n321), .ZN(n322) );
  XNOR2_X1 U332 ( .A(n371), .B(n370), .ZN(n372) );
  INV_X1 U333 ( .A(KEYINPUT23), .ZN(n327) );
  XNOR2_X1 U334 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U335 ( .A(n330), .B(n329), .ZN(n334) );
  XNOR2_X1 U336 ( .A(n379), .B(n378), .ZN(n380) );
  NOR2_X1 U337 ( .A1(n438), .A2(n534), .ZN(n576) );
  XNOR2_X1 U338 ( .A(n581), .B(KEYINPUT41), .ZN(n559) );
  NOR2_X1 U339 ( .A1(n515), .A2(n504), .ZN(n485) );
  INV_X1 U340 ( .A(G15GAT), .ZN(n486) );
  XNOR2_X1 U341 ( .A(n461), .B(G190GAT), .ZN(n462) );
  XNOR2_X1 U342 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U343 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(KEYINPUT69), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n296), .B(G29GAT), .ZN(n297) );
  XOR2_X1 U347 ( .A(n297), .B(KEYINPUT7), .Z(n299) );
  XNOR2_X1 U348 ( .A(KEYINPUT8), .B(KEYINPUT70), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n366) );
  XNOR2_X1 U350 ( .A(G36GAT), .B(G190GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n300), .B(KEYINPUT82), .ZN(n335) );
  XOR2_X1 U352 ( .A(n335), .B(KEYINPUT83), .Z(n302) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n366), .B(n303), .ZN(n316) );
  XOR2_X1 U356 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n305) );
  XNOR2_X1 U357 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U359 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n307) );
  XNOR2_X1 U360 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(n309), .B(n308), .Z(n314) );
  XOR2_X1 U363 ( .A(G99GAT), .B(G85GAT), .Z(n367) );
  XOR2_X1 U364 ( .A(KEYINPUT80), .B(G218GAT), .Z(n311) );
  XOR2_X1 U365 ( .A(G134GAT), .B(KEYINPUT81), .Z(n419) );
  XOR2_X1 U366 ( .A(G50GAT), .B(G162GAT), .Z(n320) );
  XNOR2_X1 U367 ( .A(n419), .B(n320), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n367), .B(n312), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U371 ( .A(n316), .B(n315), .Z(n565) );
  XOR2_X1 U372 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n318) );
  XNOR2_X1 U373 ( .A(G141GAT), .B(KEYINPUT91), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n427) );
  AND2_X1 U375 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XOR2_X1 U376 ( .A(KEYINPUT24), .B(n322), .Z(n326) );
  XOR2_X1 U377 ( .A(G78GAT), .B(G148GAT), .Z(n324) );
  XNOR2_X1 U378 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n368) );
  XNOR2_X1 U380 ( .A(n368), .B(KEYINPUT22), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U382 ( .A(G22GAT), .B(G155GAT), .Z(n384) );
  XNOR2_X1 U383 ( .A(n384), .B(KEYINPUT90), .ZN(n328) );
  XOR2_X1 U384 ( .A(KEYINPUT21), .B(G211GAT), .Z(n332) );
  XNOR2_X1 U385 ( .A(G204GAT), .B(G218GAT), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U387 ( .A(G197GAT), .B(n333), .Z(n340) );
  XOR2_X1 U388 ( .A(n334), .B(n340), .Z(n473) );
  XOR2_X1 U389 ( .A(G8GAT), .B(G183GAT), .Z(n385) );
  XNOR2_X1 U390 ( .A(n335), .B(KEYINPUT98), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n336), .B(KEYINPUT99), .ZN(n337) );
  XOR2_X1 U392 ( .A(n385), .B(n337), .Z(n339) );
  NAND2_X1 U393 ( .A1(G226GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n342) );
  INV_X1 U395 ( .A(n340), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n347) );
  XOR2_X1 U397 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n344) );
  XNOR2_X1 U398 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n445) );
  XNOR2_X1 U400 ( .A(G176GAT), .B(G92GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n345), .B(G64GAT), .ZN(n371) );
  XNOR2_X1 U402 ( .A(n445), .B(n371), .ZN(n346) );
  XOR2_X1 U403 ( .A(n347), .B(n346), .Z(n530) );
  XOR2_X1 U404 ( .A(KEYINPUT121), .B(n530), .Z(n411) );
  INV_X1 U405 ( .A(n565), .ZN(n553) );
  INV_X1 U406 ( .A(KEYINPUT46), .ZN(n383) );
  XOR2_X1 U407 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n349) );
  XNOR2_X1 U408 ( .A(G169GAT), .B(KEYINPUT30), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U410 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n351) );
  XNOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U413 ( .A(n353), .B(n352), .Z(n364) );
  XOR2_X1 U414 ( .A(G15GAT), .B(KEYINPUT71), .Z(n355) );
  XNOR2_X1 U415 ( .A(KEYINPUT72), .B(KEYINPUT68), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n362) );
  XOR2_X1 U417 ( .A(G113GAT), .B(G1GAT), .Z(n423) );
  XOR2_X1 U418 ( .A(G197GAT), .B(G8GAT), .Z(n357) );
  XNOR2_X1 U419 ( .A(G50GAT), .B(G36GAT), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U421 ( .A(n423), .B(n358), .Z(n360) );
  NAND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U426 ( .A(n366), .B(n365), .Z(n543) );
  XOR2_X1 U427 ( .A(n368), .B(n367), .Z(n374) );
  AND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n369) );
  XOR2_X1 U429 ( .A(G120GAT), .B(G71GAT), .Z(n446) );
  XNOR2_X1 U430 ( .A(n372), .B(n446), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U432 ( .A(KEYINPUT13), .B(G57GAT), .Z(n395) );
  XOR2_X1 U433 ( .A(n375), .B(n395), .Z(n381) );
  XOR2_X1 U434 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n377) );
  XNOR2_X1 U435 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n379) );
  XNOR2_X1 U437 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n378) );
  INV_X1 U438 ( .A(n406), .ZN(n581) );
  NAND2_X1 U439 ( .A1(n543), .A2(n559), .ZN(n382) );
  XOR2_X1 U440 ( .A(n383), .B(n382), .Z(n400) );
  XOR2_X1 U441 ( .A(G15GAT), .B(G127GAT), .Z(n441) );
  XNOR2_X1 U442 ( .A(n441), .B(n384), .ZN(n399) );
  XOR2_X1 U443 ( .A(KEYINPUT12), .B(n385), .Z(n387) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U446 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n389) );
  XNOR2_X1 U447 ( .A(G1GAT), .B(KEYINPUT84), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U449 ( .A(n391), .B(n390), .Z(n397) );
  XOR2_X1 U450 ( .A(G211GAT), .B(G78GAT), .Z(n393) );
  XNOR2_X1 U451 ( .A(G71GAT), .B(G64GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n548) );
  INV_X1 U456 ( .A(n548), .ZN(n584) );
  NAND2_X1 U457 ( .A1(n400), .A2(n584), .ZN(n401) );
  NOR2_X1 U458 ( .A1(n553), .A2(n401), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n402), .B(KEYINPUT47), .ZN(n409) );
  XNOR2_X1 U460 ( .A(KEYINPUT36), .B(KEYINPUT108), .ZN(n403) );
  XOR2_X1 U461 ( .A(n403), .B(n553), .Z(n588) );
  NOR2_X1 U462 ( .A1(n584), .A2(n588), .ZN(n404) );
  XOR2_X1 U463 ( .A(KEYINPUT45), .B(n404), .Z(n405) );
  NOR2_X1 U464 ( .A1(n406), .A2(n405), .ZN(n407) );
  INV_X1 U465 ( .A(n543), .ZN(n577) );
  NAND2_X1 U466 ( .A1(n407), .A2(n577), .ZN(n408) );
  NAND2_X1 U467 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U468 ( .A(KEYINPUT48), .B(n410), .ZN(n538) );
  NAND2_X1 U469 ( .A1(n411), .A2(n538), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n412), .B(KEYINPUT54), .ZN(n438) );
  XOR2_X1 U471 ( .A(KEYINPUT6), .B(KEYINPUT97), .Z(n414) );
  XNOR2_X1 U472 ( .A(KEYINPUT96), .B(KEYINPUT4), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U474 ( .A(KEYINPUT95), .B(KEYINPUT92), .Z(n416) );
  XNOR2_X1 U475 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U477 ( .A(n418), .B(n417), .Z(n425) );
  XOR2_X1 U478 ( .A(KEYINPUT0), .B(KEYINPUT85), .Z(n440) );
  XOR2_X1 U479 ( .A(n419), .B(n440), .Z(n421) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U484 ( .A(n426), .B(KEYINPUT93), .Z(n429) );
  XNOR2_X1 U485 ( .A(n427), .B(KEYINPUT94), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n437) );
  XOR2_X1 U487 ( .A(G155GAT), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U488 ( .A(G127GAT), .B(G57GAT), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U490 ( .A(G162GAT), .B(G85GAT), .Z(n433) );
  XNOR2_X1 U491 ( .A(G29GAT), .B(G120GAT), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U493 ( .A(n435), .B(n434), .Z(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n534) );
  NAND2_X1 U495 ( .A1(n473), .A2(n576), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n439), .B(KEYINPUT55), .ZN(n460) );
  XOR2_X1 U497 ( .A(G190GAT), .B(G134GAT), .Z(n443) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U500 ( .A(n444), .B(G99GAT), .Z(n451) );
  XOR2_X1 U501 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(n449), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n459) );
  XOR2_X1 U506 ( .A(KEYINPUT88), .B(G176GAT), .Z(n453) );
  XNOR2_X1 U507 ( .A(G113GAT), .B(G183GAT), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U509 ( .A(KEYINPUT89), .B(KEYINPUT86), .Z(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT20), .B(KEYINPUT87), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U512 ( .A(n457), .B(n456), .Z(n458) );
  XOR2_X1 U513 ( .A(n459), .B(n458), .Z(n466) );
  INV_X1 U514 ( .A(n466), .ZN(n539) );
  NAND2_X1 U515 ( .A1(n460), .A2(n539), .ZN(n573) );
  NOR2_X1 U516 ( .A1(n565), .A2(n573), .ZN(n463) );
  XNOR2_X1 U517 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n461) );
  XOR2_X1 U518 ( .A(n530), .B(KEYINPUT27), .Z(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(KEYINPUT100), .ZN(n536) );
  XOR2_X1 U520 ( .A(n473), .B(KEYINPUT28), .Z(n465) );
  XNOR2_X1 U521 ( .A(KEYINPUT64), .B(n465), .ZN(n542) );
  NOR2_X1 U522 ( .A1(n536), .A2(n542), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n468), .A2(n534), .ZN(n480) );
  AND2_X1 U525 ( .A1(n539), .A2(n530), .ZN(n469) );
  XNOR2_X1 U526 ( .A(KEYINPUT101), .B(n469), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n470), .A2(n473), .ZN(n472) );
  XOR2_X1 U528 ( .A(KEYINPUT102), .B(KEYINPUT25), .Z(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(n478) );
  NOR2_X1 U530 ( .A1(n473), .A2(n539), .ZN(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT26), .B(n474), .ZN(n575) );
  INV_X1 U532 ( .A(n575), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n536), .A2(n475), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n534), .A2(n476), .ZN(n477) );
  NAND2_X1 U535 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(KEYINPUT103), .ZN(n490) );
  NOR2_X1 U538 ( .A1(n553), .A2(n584), .ZN(n482) );
  XNOR2_X1 U539 ( .A(KEYINPUT16), .B(n482), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n490), .A2(n483), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n484), .B(KEYINPUT104), .ZN(n515) );
  NAND2_X1 U542 ( .A1(n543), .A2(n581), .ZN(n504) );
  XOR2_X1 U543 ( .A(KEYINPUT105), .B(n485), .Z(n502) );
  NAND2_X1 U544 ( .A1(n502), .A2(n539), .ZN(n489) );
  XOR2_X1 U545 ( .A(KEYINPUT35), .B(KEYINPUT107), .Z(n487) );
  INV_X1 U546 ( .A(G106GAT), .ZN(n497) );
  NAND2_X1 U547 ( .A1(n584), .A2(n490), .ZN(n491) );
  NOR2_X1 U548 ( .A1(n491), .A2(n588), .ZN(n492) );
  XNOR2_X1 U549 ( .A(n492), .B(KEYINPUT37), .ZN(n505) );
  NAND2_X1 U550 ( .A1(n577), .A2(n559), .ZN(n516) );
  NOR2_X1 U551 ( .A1(n505), .A2(n516), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT115), .B(n493), .Z(n532) );
  NAND2_X1 U553 ( .A1(n532), .A2(n542), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT116), .B(KEYINPUT44), .Z(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(G1339GAT) );
  NAND2_X1 U557 ( .A1(n534), .A2(n502), .ZN(n500) );
  XNOR2_X1 U558 ( .A(G1GAT), .B(KEYINPUT106), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n498), .B(KEYINPUT34), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(G1324GAT) );
  NAND2_X1 U561 ( .A1(n530), .A2(n502), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(G8GAT), .ZN(G1325GAT) );
  NAND2_X1 U563 ( .A1(n542), .A2(n502), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT109), .B(KEYINPUT39), .Z(n508) );
  NOR2_X1 U566 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n506), .B(KEYINPUT38), .ZN(n513) );
  NAND2_X1 U568 ( .A1(n513), .A2(n534), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U570 ( .A(n509), .B(G29GAT), .Z(G1328GAT) );
  NAND2_X1 U571 ( .A1(n513), .A2(n530), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n510), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U573 ( .A1(n513), .A2(n539), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(KEYINPUT40), .ZN(n512) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n542), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U578 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U579 ( .A(n517), .B(KEYINPUT110), .ZN(n525) );
  NAND2_X1 U580 ( .A1(n534), .A2(n525), .ZN(n520) );
  XOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT111), .Z(n518) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(n518), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U584 ( .A1(n525), .A2(n530), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(KEYINPUT112), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(n522), .ZN(G1333GAT) );
  XOR2_X1 U587 ( .A(G71GAT), .B(KEYINPUT113), .Z(n524) );
  NAND2_X1 U588 ( .A1(n525), .A2(n539), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT43), .B(KEYINPUT114), .Z(n527) );
  NAND2_X1 U591 ( .A1(n525), .A2(n542), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G78GAT), .B(n528), .ZN(G1335GAT) );
  NAND2_X1 U594 ( .A1(n532), .A2(n534), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(n529), .ZN(G1336GAT) );
  NAND2_X1 U596 ( .A1(n530), .A2(n532), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n539), .A2(n532), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(G99GAT), .ZN(G1338GAT) );
  INV_X1 U600 ( .A(n534), .ZN(n535) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  AND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n557) );
  NAND2_X1 U603 ( .A1(n557), .A2(n539), .ZN(n540) );
  XOR2_X1 U604 ( .A(KEYINPUT117), .B(n540), .Z(n541) );
  NOR2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n554), .A2(n543), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U609 ( .A1(n554), .A2(n559), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(n547), .ZN(G1341GAT) );
  NAND2_X1 U612 ( .A1(n548), .A2(n554), .ZN(n552) );
  XOR2_X1 U613 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n550) );
  XNOR2_X1 U614 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n556), .B(n555), .ZN(G1343GAT) );
  NAND2_X1 U620 ( .A1(n557), .A2(n575), .ZN(n564) );
  NOR2_X1 U621 ( .A1(n577), .A2(n564), .ZN(n558) );
  XOR2_X1 U622 ( .A(G141GAT), .B(n558), .Z(G1344GAT) );
  INV_X1 U623 ( .A(n559), .ZN(n570) );
  NOR2_X1 U624 ( .A1(n570), .A2(n564), .ZN(n561) );
  XNOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U628 ( .A1(n584), .A2(n564), .ZN(n563) );
  XOR2_X1 U629 ( .A(G155GAT), .B(n563), .Z(G1346GAT) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U631 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  NOR2_X1 U632 ( .A1(n577), .A2(n573), .ZN(n567) );
  XOR2_X1 U633 ( .A(G169GAT), .B(n567), .Z(G1348GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n569) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n570), .A2(n573), .ZN(n571) );
  XOR2_X1 U638 ( .A(n572), .B(n571), .Z(G1349GAT) );
  NOR2_X1 U639 ( .A1(n584), .A2(n573), .ZN(n574) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n587) );
  NOR2_X1 U642 ( .A1(n577), .A2(n587), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n587), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n587), .ZN(n585) );
  XOR2_X1 U650 ( .A(KEYINPUT124), .B(n585), .Z(n586) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n593) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U656 ( .A(KEYINPUT125), .B(n591), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(G1355GAT) );
endmodule

