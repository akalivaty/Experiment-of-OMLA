

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U321 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U322 ( .A(n371), .B(n342), .Z(n515) );
  XNOR2_X1 U323 ( .A(n308), .B(n307), .ZN(n309) );
  NOR2_X1 U324 ( .A1(n393), .A2(n392), .ZN(n483) );
  XNOR2_X1 U325 ( .A(n310), .B(n309), .ZN(n339) );
  XNOR2_X1 U326 ( .A(n428), .B(KEYINPUT33), .ZN(n429) );
  XNOR2_X1 U327 ( .A(n413), .B(KEYINPUT101), .ZN(n414) );
  NOR2_X1 U328 ( .A1(n513), .A2(n472), .ZN(n568) );
  XNOR2_X1 U329 ( .A(n415), .B(n414), .ZN(n512) );
  XOR2_X1 U330 ( .A(n574), .B(KEYINPUT41), .Z(n545) );
  XNOR2_X1 U331 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U332 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U333 ( .A(n479), .B(n478), .ZN(G1349GAT) );
  XNOR2_X1 U334 ( .A(n457), .B(n456), .ZN(G1330GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n290) );
  XNOR2_X1 U336 ( .A(G50GAT), .B(G43GAT), .ZN(n289) );
  XNOR2_X1 U337 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U338 ( .A(KEYINPUT67), .B(n291), .Z(n445) );
  XOR2_X1 U339 ( .A(G99GAT), .B(G85GAT), .Z(n427) );
  XOR2_X1 U340 ( .A(G36GAT), .B(G190GAT), .Z(n334) );
  XOR2_X1 U341 ( .A(n427), .B(n334), .Z(n293) );
  NAND2_X1 U342 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U344 ( .A(KEYINPUT9), .B(G92GAT), .Z(n295) );
  XNOR2_X1 U345 ( .A(G162GAT), .B(G106GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U347 ( .A(n297), .B(n296), .Z(n302) );
  XOR2_X1 U348 ( .A(G29GAT), .B(G134GAT), .Z(n356) );
  XOR2_X1 U349 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n299) );
  XNOR2_X1 U350 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n356), .B(n300), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U354 ( .A(n445), .B(n303), .Z(n562) );
  INV_X1 U355 ( .A(n562), .ZN(n554) );
  XOR2_X1 U356 ( .A(n554), .B(KEYINPUT99), .Z(n304) );
  XNOR2_X1 U357 ( .A(n304), .B(KEYINPUT36), .ZN(n582) );
  INV_X1 U358 ( .A(KEYINPUT100), .ZN(n411) );
  XOR2_X1 U359 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n306) );
  XNOR2_X1 U360 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n310) );
  XNOR2_X1 U362 ( .A(G197GAT), .B(G211GAT), .ZN(n308) );
  INV_X1 U363 ( .A(KEYINPUT81), .ZN(n307) );
  XOR2_X1 U364 ( .A(G78GAT), .B(G148GAT), .Z(n312) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(KEYINPUT69), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n424) );
  XOR2_X1 U367 ( .A(n424), .B(G204GAT), .Z(n318) );
  XOR2_X1 U368 ( .A(KEYINPUT83), .B(KEYINPUT3), .Z(n314) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(G155GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n316) );
  XOR2_X1 U371 ( .A(G162GAT), .B(KEYINPUT2), .Z(n315) );
  XOR2_X1 U372 ( .A(n316), .B(n315), .Z(n359) );
  XNOR2_X1 U373 ( .A(G22GAT), .B(n359), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n339), .B(n319), .ZN(n327) );
  NAND2_X1 U376 ( .A1(G228GAT), .A2(G233GAT), .ZN(n325) );
  XOR2_X1 U377 ( .A(KEYINPUT23), .B(KEYINPUT84), .Z(n321) );
  XNOR2_X1 U378 ( .A(KEYINPUT24), .B(KEYINPUT85), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U380 ( .A(G50GAT), .B(KEYINPUT22), .Z(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n473) );
  XOR2_X1 U384 ( .A(KEYINPUT64), .B(KEYINPUT28), .Z(n328) );
  XNOR2_X1 U385 ( .A(n473), .B(n328), .ZN(n527) );
  XOR2_X1 U386 ( .A(KEYINPUT77), .B(KEYINPUT17), .Z(n330) );
  XNOR2_X1 U387 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U389 ( .A(G169GAT), .B(n331), .Z(n371) );
  XOR2_X1 U390 ( .A(G8GAT), .B(G183GAT), .Z(n395) );
  XOR2_X1 U391 ( .A(KEYINPUT91), .B(n395), .Z(n333) );
  NAND2_X1 U392 ( .A1(G226GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n335) );
  XOR2_X1 U394 ( .A(n335), .B(n334), .Z(n341) );
  XOR2_X1 U395 ( .A(G92GAT), .B(KEYINPUT70), .Z(n337) );
  XNOR2_X1 U396 ( .A(G176GAT), .B(G64GAT), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U398 ( .A(G204GAT), .B(n338), .Z(n431) );
  XNOR2_X1 U399 ( .A(n339), .B(n431), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U401 ( .A(KEYINPUT27), .B(n515), .ZN(n382) );
  XOR2_X1 U402 ( .A(KEYINPUT6), .B(G57GAT), .Z(n344) );
  XNOR2_X1 U403 ( .A(G148GAT), .B(G85GAT), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U405 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n346) );
  XNOR2_X1 U406 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U408 ( .A(n348), .B(n347), .Z(n353) );
  XOR2_X1 U409 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n350) );
  NAND2_X1 U410 ( .A1(G225GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U412 ( .A(KEYINPUT5), .B(n351), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U414 ( .A(G1GAT), .B(G127GAT), .Z(n406) );
  XOR2_X1 U415 ( .A(n354), .B(n406), .Z(n358) );
  XNOR2_X1 U416 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n355), .B(G120GAT), .ZN(n370) );
  XNOR2_X1 U418 ( .A(n370), .B(n356), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n360) );
  XOR2_X1 U420 ( .A(n360), .B(n359), .Z(n391) );
  XNOR2_X1 U421 ( .A(KEYINPUT90), .B(n391), .ZN(n513) );
  NAND2_X1 U422 ( .A1(n382), .A2(n513), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n361), .B(KEYINPUT92), .ZN(n524) );
  NOR2_X1 U424 ( .A1(n527), .A2(n524), .ZN(n378) );
  NAND2_X1 U425 ( .A1(G227GAT), .A2(G233GAT), .ZN(n367) );
  XOR2_X1 U426 ( .A(G183GAT), .B(G99GAT), .Z(n363) );
  XNOR2_X1 U427 ( .A(G43GAT), .B(G15GAT), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U429 ( .A(G134GAT), .B(G190GAT), .Z(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n377) );
  XOR2_X1 U432 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n369) );
  XNOR2_X1 U433 ( .A(G176GAT), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n373) );
  XOR2_X1 U436 ( .A(G71GAT), .B(KEYINPUT78), .Z(n372) );
  XNOR2_X1 U437 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U438 ( .A(n375), .B(n374), .Z(n376) );
  XOR2_X1 U439 ( .A(n377), .B(n376), .Z(n384) );
  NAND2_X1 U440 ( .A1(n378), .A2(n384), .ZN(n379) );
  XNOR2_X1 U441 ( .A(KEYINPUT93), .B(n379), .ZN(n393) );
  INV_X1 U442 ( .A(n384), .ZN(n453) );
  NOR2_X1 U443 ( .A1(n453), .A2(n473), .ZN(n381) );
  XNOR2_X1 U444 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n567) );
  NAND2_X1 U446 ( .A1(n567), .A2(n382), .ZN(n383) );
  XNOR2_X1 U447 ( .A(KEYINPUT95), .B(n383), .ZN(n389) );
  INV_X1 U448 ( .A(n515), .ZN(n470) );
  NOR2_X1 U449 ( .A1(n384), .A2(n470), .ZN(n385) );
  XOR2_X1 U450 ( .A(KEYINPUT96), .B(n385), .Z(n386) );
  NAND2_X1 U451 ( .A1(n386), .A2(n473), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n387), .B(KEYINPUT25), .ZN(n388) );
  NOR2_X1 U453 ( .A1(n389), .A2(n388), .ZN(n390) );
  NOR2_X1 U454 ( .A1(n391), .A2(n390), .ZN(n392) );
  XOR2_X1 U455 ( .A(G15GAT), .B(G22GAT), .Z(n438) );
  XNOR2_X1 U456 ( .A(G71GAT), .B(G57GAT), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n394), .B(KEYINPUT13), .ZN(n423) );
  XNOR2_X1 U458 ( .A(n438), .B(n423), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U460 ( .A(KEYINPUT14), .B(KEYINPUT75), .Z(n398) );
  NAND2_X1 U461 ( .A1(G231GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U463 ( .A(n400), .B(n399), .Z(n405) );
  XOR2_X1 U464 ( .A(KEYINPUT74), .B(KEYINPUT15), .Z(n402) );
  XNOR2_X1 U465 ( .A(G78GAT), .B(G64GAT), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n403), .B(KEYINPUT12), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U469 ( .A(n407), .B(n406), .Z(n409) );
  XNOR2_X1 U470 ( .A(G211GAT), .B(G155GAT), .ZN(n408) );
  XOR2_X1 U471 ( .A(n409), .B(n408), .Z(n480) );
  NOR2_X1 U472 ( .A1(n483), .A2(n480), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n412) );
  NOR2_X1 U474 ( .A1(n582), .A2(n412), .ZN(n415) );
  INV_X1 U475 ( .A(KEYINPUT37), .ZN(n413) );
  INV_X1 U476 ( .A(KEYINPUT32), .ZN(n416) );
  NAND2_X1 U477 ( .A1(KEYINPUT31), .A2(n416), .ZN(n419) );
  INV_X1 U478 ( .A(KEYINPUT31), .ZN(n417) );
  NAND2_X1 U479 ( .A1(n417), .A2(KEYINPUT32), .ZN(n418) );
  NAND2_X1 U480 ( .A1(n419), .A2(n418), .ZN(n421) );
  NAND2_X1 U481 ( .A1(G230GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U483 ( .A(n422), .B(KEYINPUT71), .Z(n426) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U486 ( .A(G120GAT), .B(n427), .Z(n428) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n574) );
  XOR2_X1 U488 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n434) );
  XNOR2_X1 U489 ( .A(G8GAT), .B(G1GAT), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n449) );
  XOR2_X1 U491 ( .A(G141GAT), .B(G197GAT), .Z(n436) );
  XNOR2_X1 U492 ( .A(G29GAT), .B(G36GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U494 ( .A(n437), .B(G113GAT), .Z(n440) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U497 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n442) );
  NAND2_X1 U498 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U500 ( .A(n444), .B(n443), .Z(n447) );
  XNOR2_X1 U501 ( .A(n445), .B(KEYINPUT68), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(n449), .B(n448), .Z(n528) );
  NAND2_X1 U504 ( .A1(n574), .A2(n528), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n450), .B(KEYINPUT72), .ZN(n486) );
  OR2_X1 U506 ( .A1(n512), .A2(n486), .ZN(n452) );
  INV_X1 U507 ( .A(KEYINPUT38), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(n499) );
  AND2_X1 U509 ( .A1(n499), .A2(n453), .ZN(n457) );
  XNOR2_X1 U510 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n455) );
  INV_X1 U511 ( .A(G43GAT), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n480), .B(KEYINPUT108), .ZN(n560) );
  XNOR2_X1 U513 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n459) );
  INV_X1 U514 ( .A(n528), .ZN(n569) );
  NOR2_X1 U515 ( .A1(n569), .A2(n545), .ZN(n458) );
  XOR2_X1 U516 ( .A(n459), .B(n458), .Z(n460) );
  NOR2_X1 U517 ( .A1(n560), .A2(n460), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(KEYINPUT110), .ZN(n462) );
  NAND2_X1 U519 ( .A1(n462), .A2(n554), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n463), .B(KEYINPUT47), .ZN(n468) );
  INV_X1 U521 ( .A(n480), .ZN(n577) );
  NOR2_X1 U522 ( .A1(n582), .A2(n577), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n464), .B(KEYINPUT45), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n465), .A2(n574), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n466), .A2(n528), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U527 ( .A(KEYINPUT48), .B(n469), .ZN(n523) );
  NOR2_X1 U528 ( .A1(n523), .A2(n470), .ZN(n471) );
  XOR2_X1 U529 ( .A(KEYINPUT54), .B(n471), .Z(n472) );
  NAND2_X1 U530 ( .A1(n568), .A2(n473), .ZN(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT55), .B(n474), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n475), .A2(n453), .ZN(n556) );
  INV_X1 U533 ( .A(n556), .ZN(n563) );
  XNOR2_X1 U534 ( .A(KEYINPUT103), .B(n545), .ZN(n532) );
  AND2_X1 U535 ( .A1(n563), .A2(n532), .ZN(n479) );
  XNOR2_X1 U536 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n477) );
  XNOR2_X1 U537 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n476) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n488) );
  XOR2_X1 U539 ( .A(KEYINPUT76), .B(KEYINPUT16), .Z(n482) );
  NAND2_X1 U540 ( .A1(n480), .A2(n554), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(n485) );
  INV_X1 U542 ( .A(n483), .ZN(n484) );
  NAND2_X1 U543 ( .A1(n485), .A2(n484), .ZN(n501) );
  NOR2_X1 U544 ( .A1(n486), .A2(n501), .ZN(n493) );
  NAND2_X1 U545 ( .A1(n493), .A2(n513), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(G1324GAT) );
  NAND2_X1 U547 ( .A1(n493), .A2(n515), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U550 ( .A1(n493), .A2(n453), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U552 ( .A(G15GAT), .B(n492), .Z(G1326GAT) );
  NAND2_X1 U553 ( .A1(n493), .A2(n527), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT98), .B(KEYINPUT39), .Z(n496) );
  NAND2_X1 U556 ( .A1(n499), .A2(n513), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n515), .A2(n499), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n499), .A2(n527), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  NAND2_X1 U564 ( .A1(n532), .A2(n569), .ZN(n511) );
  NOR2_X1 U565 ( .A1(n511), .A2(n501), .ZN(n507) );
  NAND2_X1 U566 ( .A1(n507), .A2(n513), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U568 ( .A1(n507), .A2(n515), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U570 ( .A1(n507), .A2(n453), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n505), .B(KEYINPUT104), .ZN(n506) );
  XNOR2_X1 U572 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U574 ( .A1(n507), .A2(n527), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n510), .Z(G1335GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n513), .A2(n520), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n520), .A2(n515), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(KEYINPUT106), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT107), .Z(n519) );
  NAND2_X1 U584 ( .A1(n520), .A2(n453), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n520), .A2(n527), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n530) );
  NOR2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n543) );
  NAND2_X1 U591 ( .A1(n453), .A2(n543), .ZN(n525) );
  XOR2_X1 U592 ( .A(KEYINPUT111), .B(n525), .Z(n526) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n539), .A2(n528), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  AND2_X1 U597 ( .A1(n532), .A2(n539), .ZN(n534) );
  XNOR2_X1 U598 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n537) );
  NAND2_X1 U602 ( .A1(n539), .A2(n560), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n541) );
  NAND2_X1 U606 ( .A1(n539), .A2(n562), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n543), .A2(n567), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n569), .A2(n553), .ZN(n544) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n545), .A2(n553), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(KEYINPUT52), .B(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n577), .A2(n553), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(G1346GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  NOR2_X1 U623 ( .A1(n569), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(n566), .ZN(G1351GAT) );
  XNOR2_X1 U633 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n581) );
  NOR2_X1 U635 ( .A1(n569), .A2(n581), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n581), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n581), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n580) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(n584), .B(n583), .Z(G1355GAT) );
endmodule

