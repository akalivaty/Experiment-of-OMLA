//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n546, new_n547, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n606, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n460), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n461), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g047(.A(new_n472), .B(KEYINPUT69), .Z(G160));
  NAND2_X1  g048(.A1(new_n462), .A2(new_n464), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n460), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND4_X1  g057(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n460), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n460), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  MUX2_X1   g064(.A(KEYINPUT4), .B(new_n484), .S(KEYINPUT71), .Z(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(new_n483), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n489), .A2(new_n491), .ZN(G164));
  INV_X1    g067(.A(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT6), .B(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n500), .A2(new_n506), .ZN(G303));
  INV_X1    g082(.A(G303), .ZN(G166));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n509));
  NAND3_X1  g084(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(new_n510), .B(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT7), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(KEYINPUT7), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G89), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n513), .B(new_n516), .C1(new_n517), .C2(new_n502), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n497), .A2(new_n501), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n521), .A2(new_n522), .A3(new_n513), .A4(new_n516), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n497), .A2(G63), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n504), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n509), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  AOI211_X1 g104(.A(KEYINPUT74), .B(new_n527), .C1(new_n519), .C2(new_n523), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AOI22_X1  g107(.A1(new_n497), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n499), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n502), .A2(new_n535), .B1(new_n504), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n497), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n499), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n502), .A2(new_n541), .B1(new_n504), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n546), .A2(new_n550), .ZN(G188));
  AND2_X1   g126(.A1(new_n501), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G53), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT9), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n497), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n499), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n520), .A2(KEYINPUT76), .A3(G91), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n502), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n554), .A2(new_n556), .A3(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  NAND2_X1  g138(.A1(new_n520), .A2(G87), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n552), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  AOI22_X1  g142(.A1(new_n520), .A2(G86), .B1(G48), .B2(new_n552), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n497), .A2(G61), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT77), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n499), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT78), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n574));
  AOI211_X1 g149(.A(new_n574), .B(new_n499), .C1(new_n569), .C2(new_n571), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n568), .B1(new_n573), .B2(new_n575), .ZN(G305));
  XNOR2_X1  g151(.A(KEYINPUT79), .B(G85), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n520), .A2(new_n577), .B1(new_n552), .B2(G47), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n499), .B2(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n494), .A2(new_n496), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  INV_X1    g161(.A(G54), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n504), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n586), .B(KEYINPUT80), .C1(new_n587), .C2(new_n504), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n497), .A2(G92), .A3(new_n501), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(KEYINPUT10), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n590), .A2(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n581), .B1(new_n595), .B2(G868), .ZN(G321));
  XNOR2_X1  g171(.A(G321), .B(KEYINPUT81), .ZN(G284));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(G868), .B2(new_n599), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(G868), .B2(new_n599), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT82), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g182(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n608));
  XNOR2_X1  g183(.A(G323), .B(new_n608), .ZN(G282));
  INV_X1    g184(.A(new_n474), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n469), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT13), .Z(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n475), .A2(G123), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n477), .A2(G135), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n460), .A2(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n613), .A2(G2100), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n614), .A2(new_n620), .A3(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2443), .B(G2446), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n635), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(G401));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT85), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2072), .B(G2078), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n640), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n641), .B(KEYINPUT17), .Z(new_n646));
  OAI211_X1 g221(.A(new_n642), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT86), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n643), .A2(new_n639), .A3(new_n641), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n640), .A2(new_n644), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2096), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT87), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n657), .A3(new_n659), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n657), .B2(new_n659), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n657), .B2(new_n659), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G1991), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(G229));
  INV_X1    g252(.A(KEYINPUT24), .ZN(new_n678));
  INV_X1    g253(.A(G34), .ZN(new_n679));
  AOI21_X1  g254(.A(G29), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n678), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G29), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(G160), .B2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(G2084), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(G33), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n469), .A2(G103), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT25), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n610), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(new_n460), .ZN(new_n689));
  AOI211_X1 g264(.A(new_n687), .B(new_n689), .C1(G139), .C2(new_n477), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n685), .B1(new_n690), .B2(new_n682), .ZN(new_n691));
  NOR2_X1   g266(.A1(G5), .A2(G16), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G171), .B2(G16), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n691), .A2(G2072), .B1(G1961), .B2(new_n693), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n684), .B(new_n694), .C1(G2072), .C2(new_n691), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G2084), .B2(new_n683), .ZN(new_n696));
  NOR2_X1   g271(.A1(G16), .A2(G21), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G168), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT93), .B(G1966), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT92), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n700), .ZN(new_n702));
  NOR2_X1   g277(.A1(G29), .A2(G32), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT26), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G105), .B2(new_n469), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n475), .A2(G129), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n477), .A2(G141), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n703), .B1(new_n710), .B2(G29), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT27), .B(G1996), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G164), .A2(new_n682), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G27), .B2(new_n682), .ZN(new_n715));
  INV_X1    g290(.A(G2078), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G28), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n719));
  AOI21_X1  g294(.A(G29), .B1(new_n718), .B2(KEYINPUT30), .ZN(new_n720));
  OR2_X1    g295(.A1(KEYINPUT31), .A2(G11), .ZN(new_n721));
  NAND2_X1  g296(.A1(KEYINPUT31), .A2(G11), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n723), .B1(new_n682), .B2(new_n619), .C1(new_n693), .C2(G1961), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n715), .A2(new_n716), .ZN(new_n725));
  NOR4_X1   g300(.A1(new_n713), .A2(new_n717), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n696), .A2(new_n701), .A3(new_n702), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT94), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G4), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n595), .B2(new_n731), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1348), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT23), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n731), .A2(G20), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n735), .B(new_n736), .C1(G299), .C2(G16), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT95), .B(G1956), .Z(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n739), .B2(new_n738), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n682), .A2(G26), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n475), .A2(G128), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n477), .A2(G140), .ZN(new_n744));
  OR2_X1    g319(.A1(G104), .A2(G2105), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n745), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n742), .B1(new_n747), .B2(G29), .ZN(new_n748));
  MUX2_X1   g323(.A(new_n742), .B(new_n748), .S(KEYINPUT28), .Z(new_n749));
  INV_X1    g324(.A(G2067), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n682), .A2(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n682), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT29), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2090), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n731), .A2(G19), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n544), .B2(new_n731), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(G1341), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n733), .A2(G1348), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n749), .A2(new_n750), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n741), .A2(new_n751), .A3(new_n755), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n729), .A2(new_n730), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT96), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n731), .A2(G22), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G166), .B2(new_n731), .ZN(new_n766));
  INV_X1    g341(.A(G1971), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n731), .A2(G6), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G305), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT32), .B(G1981), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT90), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G23), .ZN(new_n774));
  INV_X1    g349(.A(G288), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT33), .B(G1976), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n768), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n770), .A2(new_n772), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT34), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR3_X1    g356(.A1(new_n779), .A2(KEYINPUT34), .A3(new_n780), .ZN(new_n782));
  MUX2_X1   g357(.A(G24), .B(G290), .S(G16), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1986), .ZN(new_n784));
  AOI22_X1  g359(.A1(G119), .A2(new_n475), .B1(new_n477), .B2(G131), .ZN(new_n785));
  NOR3_X1   g360(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n786));
  OAI21_X1  g361(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n785), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G25), .B(new_n789), .S(G29), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT35), .B(G1991), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n782), .A2(KEYINPUT91), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(KEYINPUT91), .B1(new_n782), .B2(new_n793), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n781), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT36), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n764), .A2(new_n797), .ZN(G150));
  INV_X1    g373(.A(G150), .ZN(G311));
  XNOR2_X1  g374(.A(KEYINPUT98), .B(G93), .ZN(new_n800));
  INV_X1    g375(.A(G55), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n502), .A2(new_n800), .B1(new_n504), .B2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G80), .A2(G543), .ZN(new_n805));
  INV_X1    g380(.A(G67), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n583), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G651), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT97), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n544), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n595), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n813), .A2(new_n816), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n817), .A2(new_n818), .A3(G860), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n810), .A2(G860), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT37), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n819), .A2(new_n821), .ZN(G145));
  NAND2_X1  g397(.A1(new_n690), .A2(KEYINPUT100), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n709), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n612), .B(KEYINPUT102), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(G160), .B(new_n619), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n789), .B(G162), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n826), .B(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n489), .A2(new_n491), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n747), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n477), .A2(G142), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT101), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n475), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n460), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n832), .B(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(G37), .B1(new_n830), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n830), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g417(.A(new_n605), .B(new_n812), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n590), .A2(new_n591), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n593), .A2(new_n594), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n599), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n595), .A2(G299), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT41), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n595), .A2(G299), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n595), .A2(G299), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n847), .A2(KEYINPUT41), .A3(new_n848), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n843), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT42), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR3_X1    g436(.A1(new_n850), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(G303), .B(G290), .Z(new_n863));
  XNOR2_X1  g438(.A(G305), .B(G288), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n859), .B2(new_n860), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n861), .B1(new_n850), .B2(new_n858), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n862), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n862), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g444(.A(G868), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n810), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(G868), .B2(new_n871), .ZN(G295));
  OAI21_X1  g447(.A(new_n870), .B1(G868), .B2(new_n871), .ZN(G331));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n849), .A2(KEYINPUT104), .A3(new_n851), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n856), .B2(KEYINPUT104), .ZN(new_n876));
  NAND2_X1  g451(.A1(G286), .A2(G301), .ZN(new_n877));
  OAI21_X1  g452(.A(G171), .B1(new_n529), .B2(new_n530), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n877), .A2(new_n812), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n812), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n813), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n877), .A2(new_n812), .A3(new_n878), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n883), .A2(new_n884), .B1(new_n847), .B2(new_n848), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n865), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n849), .B1(new_n879), .B2(new_n880), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(new_n856), .A3(new_n884), .ZN(new_n890));
  INV_X1    g465(.A(new_n865), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n895));
  OAI211_X1 g470(.A(KEYINPUT105), .B(new_n865), .C1(new_n881), .C2(new_n885), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n888), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n897), .A2(KEYINPUT106), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n889), .A2(new_n890), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n865), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n897), .B2(KEYINPUT106), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n874), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  AND4_X1   g479(.A1(KEYINPUT43), .A2(new_n888), .A3(new_n894), .A4(new_n896), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT43), .B1(new_n894), .B2(new_n900), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT44), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(G397));
  INV_X1    g483(.A(G1384), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n489), .B2(new_n491), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G40), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n467), .A2(new_n471), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n915));
  NOR3_X1   g490(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n747), .B(new_n750), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT108), .ZN(new_n918));
  INV_X1    g493(.A(G1996), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n709), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n789), .A2(new_n791), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n789), .A2(new_n791), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n918), .A2(new_n920), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G290), .B(G1986), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n916), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(G299), .B(KEYINPUT57), .Z(new_n926));
  OAI211_X1 g501(.A(KEYINPUT45), .B(new_n909), .C1(new_n489), .C2(new_n491), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n927), .A2(new_n472), .ZN(new_n928));
  INV_X1    g503(.A(new_n915), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n912), .B1(new_n910), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(KEYINPUT56), .B(G2072), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n910), .A2(KEYINPUT50), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT114), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT50), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n937), .B(new_n909), .C1(new_n489), .C2(new_n491), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n911), .A2(new_n935), .A3(new_n937), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n913), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1956), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n926), .B1(new_n933), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n943), .A2(new_n926), .A3(new_n933), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n946), .A2(new_n846), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n938), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n914), .B1(new_n949), .B2(new_n934), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n910), .A2(new_n948), .A3(KEYINPUT50), .ZN(new_n951));
  AOI21_X1  g526(.A(G1348), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT116), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n914), .B2(new_n910), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n831), .A2(KEYINPUT116), .A3(new_n909), .A4(new_n913), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(G2067), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT117), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n952), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n952), .B2(new_n957), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n945), .B1(new_n947), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n928), .A2(new_n919), .A3(new_n930), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT58), .B(G1341), .Z(new_n964));
  AOI22_X1  g539(.A1(new_n963), .A2(KEYINPUT118), .B1(new_n956), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT118), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n931), .A2(new_n966), .A3(new_n919), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n544), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT119), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT119), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n971), .A3(new_n544), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(KEYINPUT59), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT59), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n971), .B1(new_n968), .B2(new_n544), .ZN(new_n975));
  AOI211_X1 g550(.A(KEYINPUT119), .B(new_n811), .C1(new_n965), .C2(new_n967), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT120), .B1(new_n946), .B2(new_n944), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(KEYINPUT120), .B(KEYINPUT61), .C1(new_n946), .C2(new_n944), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n961), .A2(KEYINPUT60), .A3(new_n846), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n846), .B1(new_n961), .B2(KEYINPUT60), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n984), .A2(new_n985), .B1(KEYINPUT60), .B2(new_n961), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n962), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n949), .A2(new_n934), .ZN(new_n988));
  INV_X1    g563(.A(G2090), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n988), .A2(new_n989), .A3(new_n913), .A4(new_n951), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n928), .A2(new_n930), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n767), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n950), .A2(KEYINPUT110), .A3(new_n989), .A4(new_n951), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT111), .ZN(new_n997));
  AOI22_X1  g572(.A1(G303), .A2(G8), .B1(KEYINPUT112), .B2(KEYINPUT55), .ZN(new_n998));
  OR2_X1    g573(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n998), .B(new_n999), .Z(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n992), .A2(new_n1001), .A3(new_n994), .A4(new_n995), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n997), .A2(G8), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n994), .B1(new_n941), .B2(G2090), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G8), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1000), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(G305), .A2(G1981), .ZN(new_n1008));
  INV_X1    g583(.A(new_n568), .ZN(new_n1009));
  OAI21_X1  g584(.A(G1981), .B1(new_n1009), .B2(new_n572), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT49), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT113), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n911), .A2(new_n913), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G8), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1016), .ZN(new_n1018));
  INV_X1    g593(.A(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1018), .B(new_n1020), .C1(new_n1019), .C2(G288), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1016), .B1(G1976), .B2(new_n775), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1003), .A2(new_n1007), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT123), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1003), .A2(KEYINPUT123), .A3(new_n1025), .A4(new_n1007), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n931), .B2(new_n716), .ZN(new_n1031));
  INV_X1    g606(.A(G1961), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n950), .A2(new_n951), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G171), .B(KEYINPUT54), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n468), .A2(KEYINPUT121), .A3(new_n470), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT121), .B1(new_n468), .B2(new_n470), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n467), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n930), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(KEYINPUT122), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(KEYINPUT122), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1041), .A2(KEYINPUT53), .A3(new_n716), .A4(new_n927), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1034), .B(new_n1035), .C1(new_n1040), .C2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n911), .A2(KEYINPUT45), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n913), .B1(new_n910), .B2(new_n929), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(KEYINPUT53), .A3(new_n716), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1034), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1043), .B1(new_n1048), .B2(new_n1035), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT115), .B1(new_n1046), .B2(new_n699), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n1052));
  INV_X1    g627(.A(new_n699), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1052), .B(new_n1053), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1051), .B(new_n1054), .C1(G2084), .C2(new_n1033), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1050), .B(G8), .C1(new_n1055), .C2(G286), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G286), .A2(G8), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1050), .B(new_n1058), .C1(new_n1055), .C2(G8), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1049), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1030), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT124), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1030), .A2(new_n1067), .A3(new_n1064), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n987), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1017), .A2(G1976), .A3(G288), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1008), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1018), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1025), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n1003), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT63), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1055), .A2(G8), .A3(G168), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1026), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n997), .A2(G8), .A3(new_n1002), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1006), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1076), .A2(new_n1075), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n1003), .A4(new_n1025), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1074), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT62), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT125), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1060), .A2(new_n1062), .A3(KEYINPUT62), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT125), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1086), .B(KEYINPUT62), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1048), .A2(G301), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1030), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1082), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n925), .B1(new_n1069), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G290), .A2(G1986), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n916), .A2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1094), .B(KEYINPUT48), .Z(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n923), .B2(new_n916), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT126), .B(KEYINPUT46), .Z(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n916), .B2(new_n919), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n919), .B1(KEYINPUT126), .B2(KEYINPUT46), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n918), .A2(new_n710), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1100), .B2(new_n916), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT47), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n918), .A2(new_n920), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1103), .A2(new_n922), .B1(G2067), .B2(new_n747), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n1096), .B(new_n1102), .C1(new_n916), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1092), .A2(new_n1105), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g681(.A1(new_n898), .A2(new_n903), .ZN(new_n1108));
  INV_X1    g682(.A(G319), .ZN(new_n1109));
  NOR3_X1   g683(.A1(G401), .A2(new_n1109), .A3(G227), .ZN(new_n1110));
  NAND4_X1  g684(.A1(new_n841), .A2(new_n675), .A3(new_n676), .A4(new_n1110), .ZN(new_n1111));
  NOR2_X1   g685(.A1(new_n1108), .A2(new_n1111), .ZN(G308));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1113));
  OAI21_X1  g687(.A(new_n1113), .B1(new_n898), .B2(new_n903), .ZN(G225));
endmodule


