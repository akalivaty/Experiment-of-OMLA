//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT79), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n193), .A3(new_n197), .A4(new_n194), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(G101), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n190), .A2(new_n193), .A3(new_n200), .A4(new_n194), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n201), .A2(KEYINPUT4), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT4), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n196), .A2(new_n204), .A3(G101), .A4(new_n198), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT67), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G119), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(G116), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n206), .A2(G116), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n210), .A2(KEYINPUT68), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT68), .B1(new_n210), .B2(new_n211), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT2), .B(G113), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n211), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(new_n214), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n203), .B(new_n205), .C1(new_n216), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n194), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n189), .A2(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n201), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT5), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n210), .A2(KEYINPUT68), .A3(new_n211), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(G113), .B1(new_n210), .B2(KEYINPUT5), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n224), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G110), .B(G122), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n219), .A2(new_n233), .A3(new_n231), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(KEYINPUT6), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n232), .A2(new_n238), .A3(new_n234), .ZN(new_n239));
  INV_X1    g053(.A(G143), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(G146), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  INV_X1    g056(.A(G146), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(G143), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(KEYINPUT66), .A3(G146), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n241), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n240), .A2(G146), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT0), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT64), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(KEYINPUT0), .B2(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n248), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n251), .B2(new_n257), .ZN(new_n261));
  OAI21_X1  g075(.A(G125), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n240), .A2(KEYINPUT66), .A3(G146), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT66), .B1(new_n240), .B2(G146), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n249), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(G143), .B2(new_n243), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n243), .A2(G143), .ZN(new_n269));
  OAI22_X1  g083(.A1(new_n268), .A2(new_n253), .B1(new_n241), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G125), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n262), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G224), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G953), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n237), .A2(new_n239), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT83), .A2(KEYINPUT7), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n262), .A2(new_n274), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT7), .B1(new_n276), .B2(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n283), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n262), .A2(new_n274), .A3(new_n285), .A4(new_n281), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n236), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n233), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n229), .A2(new_n230), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n223), .B1(new_n291), .B2(new_n218), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n217), .A2(new_n225), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n224), .B1(new_n230), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n280), .B1(new_n287), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n188), .B1(new_n279), .B2(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n236), .A2(new_n284), .A3(new_n286), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n292), .A2(new_n294), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n289), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n237), .A2(new_n239), .A3(new_n278), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n187), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n297), .A2(KEYINPUT84), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT84), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n306), .B(new_n188), .C1(new_n279), .C2(new_n296), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G237), .ZN(new_n309));
  INV_X1    g123(.A(G953), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G214), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT85), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G143), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(G237), .A2(G953), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n315), .B(G214), .C1(new_n312), .C2(G143), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G131), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT17), .ZN(new_n319));
  INV_X1    g133(.A(G131), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n314), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT88), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n273), .A2(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n326), .B1(new_n329), .B2(new_n324), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n243), .ZN(new_n331));
  OAI211_X1 g145(.A(G146), .B(new_n326), .C1(new_n329), .C2(new_n324), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT88), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n318), .A2(new_n335), .A3(new_n319), .A4(new_n321), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n317), .A2(KEYINPUT17), .A3(G131), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n323), .A2(new_n334), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n327), .A2(new_n328), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT86), .B1(new_n339), .B2(new_n243), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n243), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT18), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n317), .B1(new_n345), .B2(new_n320), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT18), .A4(G131), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n338), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G113), .B(G122), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(new_n189), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n342), .A2(new_n343), .B1(new_n347), .B2(new_n346), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n337), .A2(new_n331), .A3(new_n332), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(KEYINPUT88), .B2(new_n322), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n357), .B2(new_n336), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT89), .B1(new_n358), .B2(new_n352), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n350), .A2(new_n360), .A3(new_n353), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n354), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT90), .B1(new_n362), .B2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(new_n352), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n350), .B2(new_n353), .ZN(new_n365));
  AOI211_X1 g179(.A(KEYINPUT89), .B(new_n352), .C1(new_n338), .C2(new_n349), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT90), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(new_n280), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(G475), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n240), .A2(G128), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT13), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT91), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n240), .B2(G128), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n253), .A2(KEYINPUT91), .A3(G143), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G134), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G134), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n380), .A3(new_n371), .ZN(new_n381));
  XNOR2_X1  g195(.A(G116), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n192), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G122), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G116), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n192), .B1(new_n388), .B2(KEYINPUT14), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n386), .A2(KEYINPUT92), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT92), .B1(new_n386), .B2(new_n389), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n382), .A2(new_n192), .ZN(new_n393));
  INV_X1    g207(.A(new_n381), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n380), .B1(new_n377), .B2(new_n371), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n384), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT9), .B(G234), .ZN(new_n398));
  INV_X1    g212(.A(G217), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n398), .A2(new_n399), .A3(G953), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n384), .B(new_n400), .C1(new_n392), .C2(new_n396), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n280), .ZN(new_n405));
  INV_X1    g219(.A(G478), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(KEYINPUT15), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(G902), .B1(new_n402), .B2(new_n403), .ZN(new_n409));
  INV_X1    g223(.A(new_n407), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(KEYINPUT93), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT93), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n409), .A2(new_n410), .ZN(new_n414));
  AOI211_X1 g228(.A(G902), .B(new_n407), .C1(new_n402), .C2(new_n403), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(G234), .A2(G237), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n417), .A2(G952), .A3(new_n310), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n417), .A2(G902), .A3(G953), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(G898), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n412), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n318), .A2(new_n321), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n329), .A2(KEYINPUT87), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n425), .B(KEYINPUT19), .Z(new_n426));
  OAI211_X1 g240(.A(new_n332), .B(new_n424), .C1(new_n426), .C2(G146), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n352), .B1(new_n427), .B2(new_n349), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n354), .A2(new_n428), .ZN(new_n429));
  OR2_X1    g243(.A1(G475), .A2(G902), .ZN(new_n430));
  OR3_X1    g244(.A1(new_n429), .A2(KEYINPUT20), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT20), .B1(new_n429), .B2(new_n430), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n370), .A2(new_n423), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT94), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT94), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n370), .A2(new_n423), .A3(new_n433), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n308), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G221), .B1(new_n398), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G469), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(new_n280), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n249), .B1(new_n264), .B2(new_n265), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT80), .ZN(new_n444));
  OAI21_X1  g258(.A(G128), .B1(new_n241), .B2(new_n267), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n253), .B1(new_n249), .B2(KEYINPUT1), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT80), .B1(new_n246), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n448), .A3(new_n266), .ZN(new_n449));
  INV_X1    g263(.A(new_n223), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT10), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n266), .A2(KEYINPUT69), .A3(new_n270), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT69), .B1(new_n266), .B2(new_n270), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n223), .A2(new_n452), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT11), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n380), .B2(G137), .ZN(new_n460));
  INV_X1    g274(.A(G137), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(KEYINPUT11), .A3(G134), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n380), .A2(G137), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G131), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n460), .A2(new_n462), .A3(new_n320), .A4(new_n463), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n260), .A2(new_n261), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n203), .A3(new_n205), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n453), .A2(new_n458), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n472));
  NAND2_X1  g286(.A1(new_n272), .A2(new_n223), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n451), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n474), .B2(new_n467), .ZN(new_n475));
  NOR2_X1   g289(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n468), .B(new_n476), .C1(new_n451), .C2(new_n473), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n471), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n310), .A2(G227), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT78), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G140), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n471), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n451), .A2(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n470), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n467), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n478), .A2(new_n482), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n442), .B1(new_n488), .B2(G469), .ZN(new_n489));
  INV_X1    g303(.A(new_n471), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n468), .B1(new_n485), .B2(new_n470), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n482), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n483), .B(new_n471), .C1(new_n475), .C2(new_n477), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n441), .A3(new_n280), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n440), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n438), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT74), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n280), .B1(new_n498), .B2(KEYINPUT25), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT23), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT67), .B(G119), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(G128), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n206), .A2(new_n253), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n501), .B2(new_n253), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n504), .B2(new_n500), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT24), .B(G110), .Z(new_n506));
  OAI22_X1  g320(.A1(new_n505), .A2(G110), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n339), .A2(new_n243), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n332), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n505), .A2(G110), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(new_n506), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n333), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n310), .A2(G221), .A3(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT73), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n509), .A2(new_n512), .A3(new_n517), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n499), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n498), .A2(KEYINPUT25), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n399), .B1(G234), .B2(new_n280), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n521), .B2(new_n522), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT76), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n519), .A2(new_n520), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n524), .A2(G902), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT75), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n527), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n528), .A2(KEYINPUT76), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n212), .A2(new_n213), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n218), .B1(new_n538), .B2(new_n214), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n271), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n463), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n380), .A2(G137), .ZN(new_n543));
  OAI21_X1  g357(.A(G131), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n544), .A2(new_n466), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n266), .A2(new_n270), .A3(KEYINPUT69), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n251), .A2(new_n257), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT65), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n467), .A2(new_n549), .A3(new_n248), .A4(new_n259), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n539), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT28), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n539), .A2(new_n547), .A3(new_n553), .A4(new_n550), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n539), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n545), .A2(new_n271), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n315), .A2(G210), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT27), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT26), .B(G101), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n560), .A2(KEYINPUT70), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT70), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n552), .A2(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(new_n564), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n547), .B2(new_n550), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n550), .A2(new_n571), .A3(new_n557), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n556), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n564), .A3(new_n551), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT31), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n574), .A2(KEYINPUT31), .A3(new_n564), .A4(new_n551), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(G472), .A2(G902), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(KEYINPUT32), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT32), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n566), .A2(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n584));
  INV_X1    g398(.A(new_n581), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n584), .A2(new_n585), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(KEYINPUT72), .A3(KEYINPUT32), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT71), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n574), .A2(new_n551), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n565), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n568), .A2(new_n564), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT29), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n547), .A2(new_n550), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n539), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n552), .B2(new_n554), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n565), .A2(new_n596), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n592), .B1(new_n603), .B2(G472), .ZN(new_n604));
  INV_X1    g418(.A(G472), .ZN(new_n605));
  AOI211_X1 g419(.A(KEYINPUT71), .B(new_n605), .C1(new_n597), .C2(new_n602), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n537), .B1(new_n591), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT77), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n607), .B1(new_n590), .B2(new_n588), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT77), .B1(new_n612), .B2(new_n537), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n497), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n200), .ZN(G3));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n297), .A2(new_n616), .A3(new_n303), .ZN(new_n617));
  INV_X1    g431(.A(new_n305), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n187), .B1(new_n301), .B2(new_n302), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(KEYINPUT96), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n404), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n404), .A2(new_n622), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n406), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n406), .A2(new_n280), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n409), .B2(new_n406), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT98), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n634));
  INV_X1    g448(.A(new_n628), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n626), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n634), .B(new_n631), .C1(new_n636), .C2(new_n406), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n370), .A2(new_n433), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n621), .A2(new_n638), .A3(KEYINPUT99), .A4(new_n422), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n370), .A2(new_n433), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n633), .A2(new_n637), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n617), .A2(new_n620), .A3(new_n422), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n570), .B2(new_n579), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT95), .B1(new_n647), .B2(new_n605), .ZN(new_n648));
  INV_X1    g462(.A(new_n589), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT95), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(G472), .C1(new_n584), .C2(G902), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n648), .A2(new_n649), .A3(new_n496), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n537), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  AND2_X1   g470(.A1(new_n370), .A2(new_n433), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n412), .A2(new_n416), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n644), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  INV_X1    g477(.A(new_n652), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n517), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n513), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n533), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n523), .B2(new_n525), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT100), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n667), .C1(new_n523), .C2(new_n525), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n438), .A2(new_n664), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT101), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n674), .B(new_n676), .ZN(G12));
  NAND2_X1  g491(.A1(new_n591), .A2(new_n608), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT102), .B(G900), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n419), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n418), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n659), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n496), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n617), .A2(new_n620), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n678), .A2(new_n684), .A3(new_n673), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  NAND2_X1  g503(.A1(new_n593), .A2(new_n564), .ZN(new_n690));
  INV_X1    g504(.A(new_n599), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n551), .A2(new_n565), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(G902), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n605), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n591), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT40), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n682), .B(KEYINPUT39), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n496), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT103), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n698), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n304), .A2(new_n307), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT38), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n641), .A2(new_n658), .ZN(new_n706));
  NOR4_X1   g520(.A1(new_n705), .A2(new_n618), .A3(new_n668), .A4(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n703), .B(new_n707), .C1(new_n699), .C2(new_n702), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  NAND2_X1  g523(.A1(new_n638), .A2(new_n682), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n678), .A2(new_n673), .A3(new_n687), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  AOI21_X1  g527(.A(new_n441), .B1(new_n494), .B2(new_n280), .ZN(new_n714));
  AOI211_X1 g528(.A(G469), .B(G902), .C1(new_n492), .C2(new_n493), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n439), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n646), .A2(new_n609), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  AND3_X1   g535(.A1(new_n609), .A2(new_n660), .A3(new_n718), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(G116), .Z(G18));
  NAND4_X1  g537(.A1(new_n716), .A2(new_n617), .A3(new_n620), .A4(new_n439), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n437), .B2(new_n435), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n678), .A2(new_n725), .A3(new_n673), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NAND4_X1  g541(.A1(new_n641), .A2(new_n658), .A3(new_n617), .A4(new_n620), .ZN(new_n728));
  OAI21_X1  g542(.A(G472), .B1(new_n584), .B2(G902), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n579), .B1(new_n564), .B2(new_n600), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n581), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n536), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n716), .A2(new_n422), .A3(new_n439), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n728), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n387), .ZN(G24));
  NAND3_X1  g549(.A1(new_n729), .A2(new_n731), .A3(new_n668), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n710), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n621), .A3(new_n718), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n704), .B2(new_n305), .ZN(new_n741));
  AOI211_X1 g555(.A(KEYINPUT105), .B(new_n618), .C1(new_n304), .C2(new_n307), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n489), .A2(new_n495), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT104), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n489), .A2(new_n745), .A3(new_n495), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n439), .A3(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n741), .A2(new_n742), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n608), .A2(new_n582), .A3(new_n586), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(KEYINPUT42), .A3(new_n536), .A4(new_n711), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n741), .A2(new_n742), .ZN(new_n754));
  INV_X1    g568(.A(new_n747), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n609), .A2(new_n754), .A3(new_n711), .A4(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n748), .A2(KEYINPUT106), .A3(new_n609), .A4(new_n711), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n753), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  NAND4_X1  g577(.A1(new_n609), .A2(new_n754), .A3(new_n684), .A4(new_n755), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT107), .B(G134), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G36));
  NAND2_X1  g580(.A1(new_n657), .A2(new_n642), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT43), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n668), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT44), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n741), .A2(new_n742), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n771), .B2(KEYINPUT44), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(G469), .B1(new_n488), .B2(KEYINPUT45), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT108), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n776), .A2(KEYINPUT108), .B1(KEYINPUT45), .B2(new_n488), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n442), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT46), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT109), .B1(new_n779), .B2(KEYINPUT46), .ZN(new_n783));
  OAI221_X1 g597(.A(new_n495), .B1(KEYINPUT46), .B2(new_n779), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n439), .A3(new_n700), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n775), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g600(.A(KEYINPUT110), .B(G137), .Z(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(G39));
  NOR4_X1   g602(.A1(new_n773), .A2(new_n678), .A3(new_n536), .A4(new_n710), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n439), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n439), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n325), .ZN(G42));
  NOR4_X1   g610(.A1(new_n767), .A2(new_n537), .A3(new_n618), .A4(new_n440), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n716), .B(KEYINPUT111), .Z(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT112), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n798), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n705), .A3(new_n698), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n768), .A2(new_n681), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n773), .A2(new_n717), .ZN(new_n805));
  INV_X1    g619(.A(new_n736), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n697), .A2(new_n537), .A3(new_n681), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n641), .A2(new_n642), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT43), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n767), .B(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n732), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n418), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n705), .A2(new_n618), .A3(new_n718), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n813), .B1(new_n819), .B2(KEYINPUT50), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  OAI211_X1 g635(.A(KEYINPUT114), .B(new_n821), .C1(new_n817), .C2(new_n818), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n819), .A2(new_n824), .A3(KEYINPUT50), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n705), .A2(new_n618), .A3(new_n718), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n804), .A2(KEYINPUT50), .A3(new_n816), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n812), .B1(new_n823), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n820), .A2(new_n822), .B1(new_n825), .B2(new_n828), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n812), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n799), .A2(new_n440), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n793), .A2(new_n794), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n817), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n754), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n831), .A2(new_n834), .A3(KEYINPUT51), .A4(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(G952), .B(new_n310), .C1(new_n817), .C2(new_n724), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n804), .A2(new_n536), .A3(new_n805), .A4(new_n750), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT48), .Z(new_n842));
  AOI211_X1 g656(.A(new_n840), .B(new_n842), .C1(new_n638), .C2(new_n809), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT51), .B1(new_n838), .B2(new_n830), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI211_X1 g660(.A(KEYINPUT116), .B(KEYINPUT51), .C1(new_n838), .C2(new_n830), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n839), .B(new_n843), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n759), .A2(new_n760), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n756), .A2(new_n757), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n752), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n754), .A2(new_n737), .A3(new_n755), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n672), .B1(new_n591), .B2(new_n608), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n408), .A2(new_n411), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n685), .A2(new_n641), .A3(new_n855), .A4(new_n683), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n754), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n764), .A2(new_n853), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n734), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n304), .A2(new_n422), .A3(new_n305), .A4(new_n307), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n370), .A2(new_n433), .A3(new_n855), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n860), .B1(new_n643), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n653), .A2(new_n862), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n674), .A2(new_n726), .A3(new_n859), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n611), .A2(new_n613), .ZN(new_n865));
  INV_X1    g679(.A(new_n497), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n609), .B(new_n718), .C1(new_n646), .C2(new_n660), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n858), .A2(new_n864), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n852), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n668), .A2(new_n683), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n728), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n697), .A2(new_n755), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n688), .A2(new_n712), .A3(new_n738), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n870), .A2(KEYINPUT53), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n672), .B(new_n308), .C1(new_n435), .C2(new_n437), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n734), .B1(new_n879), .B2(new_n664), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n854), .A2(new_n725), .B1(new_n653), .B2(new_n862), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n868), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n764), .A2(new_n857), .A3(new_n853), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(new_n614), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n762), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n688), .A2(new_n738), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(new_n875), .A3(new_n712), .A4(new_n873), .ZN(new_n887));
  XOR2_X1   g701(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n888));
  NAND2_X1  g702(.A1(new_n874), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n878), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n849), .B1(new_n877), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n874), .A2(KEYINPUT52), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n878), .B1(new_n885), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n887), .A2(new_n889), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(KEYINPUT53), .A3(new_n762), .A4(new_n884), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n895), .A2(new_n849), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n848), .A2(new_n892), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(G952), .A2(G953), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n803), .B1(new_n899), .B2(new_n900), .ZN(G75));
  INV_X1    g715(.A(G952), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(G953), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT118), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n895), .A2(new_n897), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(G210), .A3(G902), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n237), .A2(new_n239), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n278), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n906), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n906), .B2(new_n907), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n904), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g730(.A(KEYINPUT119), .B(new_n904), .C1(new_n912), .C2(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(G51));
  INV_X1    g732(.A(new_n904), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n442), .B(KEYINPUT120), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT57), .Z(new_n921));
  AOI21_X1  g735(.A(new_n849), .B1(new_n895), .B2(new_n897), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n895), .A2(new_n897), .A3(new_n849), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n922), .B2(new_n923), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n921), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n494), .B(KEYINPUT122), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n905), .A2(G902), .A3(new_n777), .A4(new_n778), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n919), .B1(new_n930), .B2(new_n931), .ZN(G54));
  NAND2_X1  g746(.A1(new_n905), .A2(G902), .ZN(new_n933));
  INV_X1    g747(.A(new_n429), .ZN(new_n934));
  NAND2_X1  g748(.A1(KEYINPUT58), .A2(G475), .ZN(new_n935));
  OR3_X1    g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n919), .B1(new_n936), .B2(new_n937), .ZN(G60));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n636), .B(KEYINPUT123), .ZN(new_n940));
  INV_X1    g754(.A(new_n630), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n898), .B1(new_n945), .B2(KEYINPUT121), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n946), .B2(new_n924), .ZN(new_n947));
  INV_X1    g761(.A(new_n943), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT53), .B1(new_n870), .B2(new_n896), .ZN(new_n949));
  AND4_X1   g763(.A1(KEYINPUT53), .A2(new_n876), .A3(new_n762), .A4(new_n884), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT54), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n951), .B2(new_n926), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n904), .B1(new_n952), .B2(new_n940), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n939), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n943), .B(new_n940), .C1(new_n925), .C2(new_n927), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n943), .B1(new_n898), .B2(new_n892), .ZN(new_n956));
  INV_X1    g770(.A(new_n940), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n919), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n958), .A3(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n954), .A2(new_n959), .ZN(G63));
  INV_X1    g774(.A(new_n905), .ZN(new_n961));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n666), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n529), .B1(new_n961), .B2(new_n963), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n904), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n965), .A2(KEYINPUT61), .A3(new_n904), .A4(new_n966), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(G66));
  OAI21_X1  g785(.A(G953), .B1(new_n420), .B2(new_n276), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n882), .A2(new_n614), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(G953), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n908), .B1(G898), .B2(new_n310), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G69));
  NOR2_X1   g790(.A1(new_n572), .A2(new_n573), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(new_n426), .Z(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(G900), .B2(G953), .ZN(new_n979));
  INV_X1    g793(.A(new_n750), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n980), .A2(new_n537), .A3(new_n728), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n785), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n764), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n983), .A2(new_n795), .A3(new_n852), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n886), .A2(new_n712), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  AOI211_X1 g800(.A(KEYINPUT127), .B(new_n986), .C1(new_n775), .C2(new_n785), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n786), .B2(new_n985), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n984), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n979), .B1(new_n990), .B2(G953), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n992));
  INV_X1    g806(.A(new_n795), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n985), .A2(new_n708), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  INV_X1    g809(.A(new_n702), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n773), .B(new_n996), .C1(new_n643), .C2(new_n861), .ZN(new_n997));
  AOI22_X1  g811(.A1(new_n775), .A2(new_n785), .B1(new_n865), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n993), .A2(new_n995), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n310), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n992), .B1(new_n1001), .B2(new_n978), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n991), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n310), .B1(G227), .B2(G900), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G72));
  OR3_X1    g819(.A1(new_n1000), .A2(new_n614), .A3(new_n882), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  AOI21_X1  g822(.A(new_n690), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n693), .A2(new_n574), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n984), .B(new_n973), .C1(new_n987), .C2(new_n989), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n1008), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n594), .A2(new_n575), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n1008), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n877), .B2(new_n891), .ZN(new_n1015));
  NOR4_X1   g829(.A1(new_n1009), .A2(new_n1012), .A3(new_n919), .A4(new_n1015), .ZN(G57));
endmodule


