

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758;

  BUF_X1 U376 ( .A(n673), .Z(n355) );
  XNOR2_X1 U377 ( .A(n551), .B(KEYINPUT1), .ZN(n673) );
  OR2_X1 U378 ( .A1(n718), .A2(G902), .ZN(n409) );
  XNOR2_X2 U379 ( .A(G128), .B(KEYINPUT76), .ZN(n449) );
  XNOR2_X2 U380 ( .A(G116), .B(G119), .ZN(n415) );
  XNOR2_X2 U381 ( .A(n407), .B(G113), .ZN(n416) );
  XNOR2_X1 U382 ( .A(G128), .B(G119), .ZN(n484) );
  INV_X2 U383 ( .A(KEYINPUT3), .ZN(n407) );
  AND2_X2 U384 ( .A1(n425), .A2(n423), .ZN(n422) );
  XNOR2_X2 U385 ( .A(n738), .B(G146), .ZN(n481) );
  XNOR2_X2 U386 ( .A(n526), .B(n451), .ZN(n738) );
  NOR2_X1 U387 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U388 ( .A1(n755), .A2(n756), .ZN(n540) );
  OR2_X1 U389 ( .A1(n639), .A2(G902), .ZN(n394) );
  INV_X1 U390 ( .A(G953), .ZN(n741) );
  AND2_X1 U391 ( .A1(n441), .A2(n442), .ZN(n356) );
  AND2_X2 U392 ( .A1(n441), .A2(n442), .ZN(n357) );
  AND2_X1 U393 ( .A1(n441), .A2(n442), .ZN(n429) );
  NOR2_X1 U394 ( .A1(n753), .A2(n758), .ZN(n358) );
  NOR2_X1 U395 ( .A1(n753), .A2(n758), .ZN(n608) );
  XNOR2_X2 U396 ( .A(n439), .B(n365), .ZN(n588) );
  XNOR2_X2 U397 ( .A(n416), .B(n415), .ZN(n460) );
  XNOR2_X1 U398 ( .A(n555), .B(n408), .ZN(n685) );
  XNOR2_X1 U399 ( .A(KEYINPUT38), .B(KEYINPUT71), .ZN(n408) );
  XNOR2_X1 U400 ( .A(n523), .B(n404), .ZN(n527) );
  XNOR2_X1 U401 ( .A(n525), .B(n524), .ZN(n404) );
  XOR2_X1 U402 ( .A(G131), .B(G140), .Z(n513) );
  XNOR2_X1 U403 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U404 ( .A(G146), .B(G125), .Z(n482) );
  NAND2_X1 U405 ( .A1(n685), .A2(n686), .ZN(n690) );
  AND2_X1 U406 ( .A1(n594), .A2(n533), .ZN(n417) );
  XNOR2_X1 U407 ( .A(n678), .B(n456), .ZN(n598) );
  OR2_X1 U408 ( .A1(n550), .A2(n621), .ZN(n571) );
  OR2_X1 U409 ( .A1(n655), .A2(n549), .ZN(n550) );
  NOR2_X1 U410 ( .A1(n553), .A2(n503), .ZN(n505) );
  XNOR2_X1 U411 ( .A(n571), .B(KEYINPUT105), .ZN(n435) );
  XNOR2_X1 U412 ( .A(n528), .B(G478), .ZN(n544) );
  XNOR2_X1 U413 ( .A(n493), .B(KEYINPUT25), .ZN(n436) );
  OR2_X1 U414 ( .A1(n726), .A2(G902), .ZN(n437) );
  AND2_X1 U415 ( .A1(n720), .A2(KEYINPUT121), .ZN(n380) );
  NAND2_X1 U416 ( .A1(n382), .A2(n720), .ZN(n376) );
  NAND2_X1 U417 ( .A1(n383), .A2(KEYINPUT121), .ZN(n381) );
  XNOR2_X1 U418 ( .A(n448), .B(n447), .ZN(n459) );
  INV_X1 U419 ( .A(KEYINPUT4), .ZN(n447) );
  XNOR2_X1 U420 ( .A(KEYINPUT64), .B(KEYINPUT67), .ZN(n448) );
  XNOR2_X1 U421 ( .A(n449), .B(G143), .ZN(n463) );
  INV_X1 U422 ( .A(KEYINPUT83), .ZN(n462) );
  OR2_X1 U423 ( .A1(G902), .A2(G237), .ZN(n471) );
  XNOR2_X1 U424 ( .A(G116), .B(G107), .ZN(n520) );
  XOR2_X1 U425 ( .A(KEYINPUT9), .B(G122), .Z(n521) );
  XOR2_X1 U426 ( .A(KEYINPUT93), .B(KEYINPUT7), .Z(n524) );
  XNOR2_X1 U427 ( .A(n463), .B(n450), .ZN(n526) );
  INV_X1 U428 ( .A(G134), .ZN(n450) );
  XOR2_X1 U429 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n510) );
  XNOR2_X1 U430 ( .A(G143), .B(G122), .ZN(n506) );
  XNOR2_X1 U431 ( .A(n481), .B(n480), .ZN(n718) );
  XNOR2_X1 U432 ( .A(n570), .B(n569), .ZN(n577) );
  INV_X1 U433 ( .A(KEYINPUT48), .ZN(n569) );
  INV_X1 U434 ( .A(n544), .ZN(n556) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n508) );
  XNOR2_X1 U436 ( .A(n411), .B(n410), .ZN(n478) );
  XNOR2_X1 U437 ( .A(G107), .B(G101), .ZN(n410) );
  XNOR2_X1 U438 ( .A(n412), .B(G110), .ZN(n411) );
  INV_X1 U439 ( .A(G104), .ZN(n412) );
  XNOR2_X1 U440 ( .A(n431), .B(KEYINPUT73), .ZN(n630) );
  XOR2_X1 U441 ( .A(G902), .B(KEYINPUT15), .Z(n637) );
  NOR2_X1 U442 ( .A1(n385), .A2(n728), .ZN(n384) );
  NOR2_X1 U443 ( .A1(n388), .A2(G469), .ZN(n385) );
  NOR2_X1 U444 ( .A1(n690), .A2(n689), .ZN(n531) );
  XNOR2_X1 U445 ( .A(n595), .B(KEYINPUT22), .ZN(n596) );
  INV_X1 U446 ( .A(KEYINPUT69), .ZN(n595) );
  XNOR2_X1 U447 ( .A(n613), .B(KEYINPUT101), .ZN(n501) );
  XNOR2_X1 U448 ( .A(n375), .B(n366), .ZN(n553) );
  NAND2_X1 U449 ( .A1(n458), .A2(n686), .ZN(n375) );
  NOR2_X1 U450 ( .A1(n424), .A2(n364), .ZN(n423) );
  NOR2_X1 U451 ( .A1(n427), .A2(n438), .ZN(n424) );
  INV_X1 U452 ( .A(G472), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n413), .B(n478), .ZN(n406) );
  XNOR2_X1 U454 ( .A(n460), .B(n414), .ZN(n413) );
  XNOR2_X1 U455 ( .A(n443), .B(G122), .ZN(n414) );
  INV_X1 U456 ( .A(KEYINPUT16), .ZN(n443) );
  XNOR2_X1 U457 ( .A(n490), .B(n514), .ZN(n726) );
  INV_X1 U458 ( .A(n395), .ZN(n434) );
  INV_X1 U459 ( .A(KEYINPUT35), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n529), .B(KEYINPUT94), .ZN(n655) );
  INV_X1 U461 ( .A(KEYINPUT122), .ZN(n389) );
  AND2_X1 U462 ( .A1(n381), .A2(n379), .ZN(n378) );
  NAND2_X1 U463 ( .A1(n362), .A2(n376), .ZN(n377) );
  INV_X1 U464 ( .A(KEYINPUT56), .ZN(n398) );
  INV_X1 U465 ( .A(n355), .ZN(n427) );
  AND2_X1 U466 ( .A1(n384), .A2(n430), .ZN(n359) );
  XOR2_X1 U467 ( .A(n484), .B(G140), .Z(n360) );
  AND2_X1 U468 ( .A1(n427), .A2(n438), .ZN(n361) );
  INV_X1 U469 ( .A(n428), .ZN(n421) );
  AND2_X1 U470 ( .A1(n386), .A2(n359), .ZN(n362) );
  AND2_X1 U471 ( .A1(n432), .A2(n667), .ZN(n363) );
  NAND2_X1 U472 ( .A1(n598), .A2(n668), .ZN(n364) );
  INV_X1 U473 ( .A(n431), .ZN(n740) );
  NAND2_X1 U474 ( .A1(n577), .A2(n363), .ZN(n431) );
  XNOR2_X1 U475 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n365) );
  XNOR2_X1 U476 ( .A(KEYINPUT30), .B(KEYINPUT102), .ZN(n366) );
  XNOR2_X1 U477 ( .A(n639), .B(n638), .ZN(n367) );
  XOR2_X1 U478 ( .A(n721), .B(n445), .Z(n368) );
  XOR2_X1 U479 ( .A(n716), .B(n715), .Z(n369) );
  INV_X1 U480 ( .A(n720), .ZN(n388) );
  XNOR2_X1 U481 ( .A(n718), .B(n719), .ZN(n720) );
  AND2_X1 U482 ( .A1(n388), .A2(G469), .ZN(n370) );
  XNOR2_X1 U483 ( .A(KEYINPUT84), .B(n446), .ZN(n728) );
  INV_X1 U484 ( .A(n728), .ZN(n387) );
  XOR2_X1 U485 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n371) );
  INV_X1 U486 ( .A(KEYINPUT121), .ZN(n430) );
  NAND2_X1 U487 ( .A1(n636), .A2(n372), .ZN(n708) );
  XNOR2_X2 U488 ( .A(n629), .B(KEYINPUT45), .ZN(n372) );
  INV_X1 U489 ( .A(n372), .ZN(n733) );
  NAND2_X1 U490 ( .A1(n372), .A2(n630), .ZN(n632) );
  BUF_X1 U491 ( .A(n708), .Z(n373) );
  BUF_X1 U492 ( .A(n588), .Z(n374) );
  NAND2_X1 U493 ( .A1(n356), .A2(G478), .ZN(n723) );
  NAND2_X1 U494 ( .A1(n429), .A2(G472), .ZN(n440) );
  NAND2_X1 U495 ( .A1(n357), .A2(n370), .ZN(n386) );
  INV_X1 U496 ( .A(n600), .ZN(n428) );
  XNOR2_X1 U497 ( .A(n597), .B(n596), .ZN(n600) );
  BUF_X1 U498 ( .A(n593), .Z(n611) );
  XNOR2_X1 U499 ( .A(n505), .B(n504), .ZN(n579) );
  NAND2_X1 U500 ( .A1(n551), .A2(n674), .ZN(n613) );
  INV_X1 U501 ( .A(n554), .ZN(n502) );
  XNOR2_X1 U502 ( .A(n440), .B(n367), .ZN(n400) );
  NAND2_X1 U503 ( .A1(n632), .A2(n631), .ZN(n442) );
  OR2_X1 U504 ( .A1(n733), .A2(n431), .ZN(n707) );
  NAND2_X1 U505 ( .A1(n386), .A2(n384), .ZN(n383) );
  NAND2_X1 U506 ( .A1(n378), .A2(n377), .ZN(G54) );
  NAND2_X1 U507 ( .A1(n382), .A2(n380), .ZN(n379) );
  INV_X1 U508 ( .A(n356), .ZN(n382) );
  XNOR2_X1 U509 ( .A(n390), .B(n389), .ZN(G63) );
  NAND2_X1 U510 ( .A1(n391), .A2(n387), .ZN(n390) );
  XNOR2_X1 U511 ( .A(n723), .B(n392), .ZN(n391) );
  INV_X1 U512 ( .A(n724), .ZN(n392) );
  XNOR2_X2 U513 ( .A(n394), .B(n393), .ZN(n678) );
  NAND2_X1 U514 ( .A1(n541), .A2(n686), .ZN(n439) );
  XNOR2_X1 U515 ( .A(n406), .B(n461), .ZN(n470) );
  BUF_X1 U516 ( .A(n439), .Z(n395) );
  XNOR2_X1 U517 ( .A(n396), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U518 ( .A1(n400), .A2(n387), .ZN(n396) );
  XNOR2_X1 U519 ( .A(n397), .B(n371), .ZN(G60) );
  NAND2_X1 U520 ( .A1(n403), .A2(n387), .ZN(n397) );
  XNOR2_X1 U521 ( .A(n399), .B(n398), .ZN(G51) );
  NAND2_X1 U522 ( .A1(n405), .A2(n387), .ZN(n399) );
  NAND2_X1 U523 ( .A1(n358), .A2(KEYINPUT44), .ZN(n609) );
  XNOR2_X2 U524 ( .A(n402), .B(n401), .ZN(n751) );
  NAND2_X1 U525 ( .A1(n591), .A2(n592), .ZN(n402) );
  XNOR2_X1 U526 ( .A(n722), .B(n368), .ZN(n403) );
  NAND2_X1 U527 ( .A1(n422), .A2(n420), .ZN(n426) );
  XNOR2_X1 U528 ( .A(n419), .B(n589), .ZN(n593) );
  NAND2_X1 U529 ( .A1(n435), .A2(n434), .ZN(n433) );
  XNOR2_X1 U530 ( .A(n433), .B(KEYINPUT36), .ZN(n552) );
  NAND2_X1 U531 ( .A1(n588), .A2(n587), .ZN(n419) );
  INV_X1 U532 ( .A(n593), .ZN(n418) );
  NAND2_X1 U533 ( .A1(n673), .A2(n674), .ZN(n581) );
  XNOR2_X1 U534 ( .A(n717), .B(n369), .ZN(n405) );
  NAND2_X1 U535 ( .A1(n406), .A2(n729), .ZN(n737) );
  XNOR2_X2 U536 ( .A(n409), .B(G469), .ZN(n551) );
  NAND2_X1 U537 ( .A1(n418), .A2(n417), .ZN(n597) );
  NAND2_X1 U538 ( .A1(n428), .A2(n427), .ZN(n619) );
  NAND2_X1 U539 ( .A1(n421), .A2(KEYINPUT98), .ZN(n420) );
  NAND2_X1 U540 ( .A1(n428), .A2(n361), .ZN(n425) );
  XNOR2_X2 U541 ( .A(n426), .B(KEYINPUT99), .ZN(n753) );
  AND2_X2 U542 ( .A1(n708), .A2(n637), .ZN(n441) );
  NAND2_X1 U543 ( .A1(n429), .A2(G210), .ZN(n717) );
  NAND2_X1 U544 ( .A1(n357), .A2(G475), .ZN(n722) );
  NAND2_X1 U545 ( .A1(n357), .A2(G217), .ZN(n725) );
  NAND2_X1 U546 ( .A1(n577), .A2(n667), .ZN(n635) );
  INV_X1 U547 ( .A(n666), .ZN(n432) );
  XNOR2_X2 U548 ( .A(n437), .B(n436), .ZN(n668) );
  INV_X1 U549 ( .A(KEYINPUT98), .ZN(n438) );
  NAND2_X1 U550 ( .A1(n685), .A2(n502), .ZN(n503) );
  XNOR2_X1 U551 ( .A(n475), .B(n474), .ZN(n541) );
  AND2_X1 U552 ( .A1(n508), .A2(G210), .ZN(n444) );
  XNOR2_X1 U553 ( .A(KEYINPUT59), .B(KEYINPUT65), .ZN(n445) );
  XNOR2_X1 U554 ( .A(n464), .B(KEYINPUT17), .ZN(n465) );
  XNOR2_X1 U555 ( .A(n459), .B(G137), .ZN(n451) );
  XNOR2_X1 U556 ( .A(n466), .B(n465), .ZN(n468) );
  XNOR2_X1 U557 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U558 ( .A(KEYINPUT33), .B(KEYINPUT82), .ZN(n582) );
  INV_X1 U559 ( .A(KEYINPUT97), .ZN(n456) );
  XNOR2_X1 U560 ( .A(n454), .B(n444), .ZN(n455) );
  XNOR2_X1 U561 ( .A(n583), .B(n582), .ZN(n703) );
  XNOR2_X1 U562 ( .A(n481), .B(n455), .ZN(n639) );
  NOR2_X1 U563 ( .A1(G952), .A2(n741), .ZN(n446) );
  XOR2_X1 U564 ( .A(G131), .B(KEYINPUT5), .Z(n453) );
  XNOR2_X1 U565 ( .A(n460), .B(G101), .ZN(n452) );
  XNOR2_X1 U566 ( .A(n453), .B(n452), .ZN(n454) );
  INV_X1 U567 ( .A(n598), .ZN(n458) );
  NAND2_X1 U568 ( .A1(n471), .A2(G214), .ZN(n457) );
  XNOR2_X1 U569 ( .A(n457), .B(KEYINPUT86), .ZN(n686) );
  INV_X1 U570 ( .A(n459), .ZN(n461) );
  XNOR2_X1 U571 ( .A(n463), .B(n462), .ZN(n466) );
  NAND2_X1 U572 ( .A1(G224), .A2(n741), .ZN(n464) );
  XOR2_X1 U573 ( .A(n482), .B(KEYINPUT18), .Z(n467) );
  XNOR2_X1 U574 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U575 ( .A(n470), .B(n469), .ZN(n714) );
  NOR2_X1 U576 ( .A1(n637), .A2(n714), .ZN(n475) );
  NAND2_X1 U577 ( .A1(G210), .A2(n471), .ZN(n473) );
  INV_X1 U578 ( .A(KEYINPUT85), .ZN(n472) );
  BUF_X1 U579 ( .A(n541), .Z(n555) );
  XOR2_X1 U580 ( .A(n513), .B(KEYINPUT89), .Z(n477) );
  NAND2_X1 U581 ( .A1(G227), .A2(n741), .ZN(n476) );
  XNOR2_X1 U582 ( .A(n477), .B(n476), .ZN(n479) );
  XOR2_X1 U583 ( .A(KEYINPUT10), .B(n482), .Z(n514) );
  NAND2_X1 U584 ( .A1(G234), .A2(n741), .ZN(n483) );
  XOR2_X1 U585 ( .A(KEYINPUT8), .B(n483), .Z(n522) );
  NAND2_X1 U586 ( .A1(G221), .A2(n522), .ZN(n489) );
  XOR2_X1 U587 ( .A(G110), .B(KEYINPUT24), .Z(n486) );
  XNOR2_X1 U588 ( .A(G137), .B(KEYINPUT23), .ZN(n485) );
  XNOR2_X1 U589 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U590 ( .A(n360), .B(n487), .ZN(n488) );
  XNOR2_X1 U591 ( .A(n489), .B(n488), .ZN(n490) );
  INV_X1 U592 ( .A(n637), .ZN(n491) );
  NAND2_X1 U593 ( .A1(G234), .A2(n491), .ZN(n492) );
  XNOR2_X1 U594 ( .A(KEYINPUT20), .B(n492), .ZN(n494) );
  NAND2_X1 U595 ( .A1(G217), .A2(n494), .ZN(n493) );
  NAND2_X1 U596 ( .A1(n494), .A2(G221), .ZN(n495) );
  XNOR2_X1 U597 ( .A(n495), .B(KEYINPUT21), .ZN(n669) );
  NOR2_X1 U598 ( .A1(n668), .A2(n669), .ZN(n674) );
  NAND2_X1 U599 ( .A1(G237), .A2(G234), .ZN(n496) );
  XNOR2_X1 U600 ( .A(n496), .B(KEYINPUT14), .ZN(n498) );
  NAND2_X1 U601 ( .A1(G952), .A2(n498), .ZN(n701) );
  NOR2_X1 U602 ( .A1(n701), .A2(G953), .ZN(n497) );
  XNOR2_X1 U603 ( .A(n497), .B(KEYINPUT87), .ZN(n586) );
  NAND2_X1 U604 ( .A1(G902), .A2(n498), .ZN(n584) );
  NOR2_X1 U605 ( .A1(G900), .A2(n584), .ZN(n499) );
  NAND2_X1 U606 ( .A1(G953), .A2(n499), .ZN(n500) );
  NAND2_X1 U607 ( .A1(n586), .A2(n500), .ZN(n532) );
  NAND2_X1 U608 ( .A1(n501), .A2(n532), .ZN(n554) );
  XNOR2_X1 U609 ( .A(KEYINPUT78), .B(KEYINPUT39), .ZN(n504) );
  XOR2_X1 U610 ( .A(G104), .B(G113), .Z(n507) );
  XNOR2_X1 U611 ( .A(n507), .B(n506), .ZN(n512) );
  NAND2_X1 U612 ( .A1(G214), .A2(n508), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U614 ( .A(n512), .B(n511), .ZN(n515) );
  XNOR2_X1 U615 ( .A(n514), .B(n513), .ZN(n739) );
  XNOR2_X1 U616 ( .A(n515), .B(n739), .ZN(n721) );
  NOR2_X1 U617 ( .A1(n721), .A2(G902), .ZN(n519) );
  XOR2_X1 U618 ( .A(KEYINPUT13), .B(KEYINPUT92), .Z(n517) );
  XNOR2_X1 U619 ( .A(KEYINPUT91), .B(G475), .ZN(n516) );
  XNOR2_X1 U620 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U621 ( .A(n519), .B(n518), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n521), .B(n520), .ZN(n525) );
  NAND2_X1 U623 ( .A1(G217), .A2(n522), .ZN(n523) );
  XNOR2_X1 U624 ( .A(n526), .B(n527), .ZN(n724) );
  NOR2_X1 U625 ( .A1(n724), .A2(G902), .ZN(n528) );
  NAND2_X1 U626 ( .A1(n557), .A2(n544), .ZN(n529) );
  NOR2_X1 U627 ( .A1(n579), .A2(n655), .ZN(n530) );
  XNOR2_X1 U628 ( .A(n530), .B(KEYINPUT40), .ZN(n755) );
  NOR2_X1 U629 ( .A1(n556), .A2(n557), .ZN(n594) );
  INV_X1 U630 ( .A(n594), .ZN(n689) );
  XNOR2_X1 U631 ( .A(n531), .B(KEYINPUT41), .ZN(n704) );
  INV_X1 U632 ( .A(n669), .ZN(n533) );
  NAND2_X1 U633 ( .A1(n533), .A2(n532), .ZN(n534) );
  INV_X1 U634 ( .A(n668), .ZN(n602) );
  NOR2_X1 U635 ( .A1(n534), .A2(n602), .ZN(n535) );
  XOR2_X1 U636 ( .A(n535), .B(KEYINPUT68), .Z(n549) );
  NOR2_X1 U637 ( .A1(n549), .A2(n598), .ZN(n536) );
  XNOR2_X1 U638 ( .A(KEYINPUT28), .B(n536), .ZN(n538) );
  XNOR2_X1 U639 ( .A(n551), .B(KEYINPUT104), .ZN(n537) );
  NAND2_X1 U640 ( .A1(n538), .A2(n537), .ZN(n542) );
  NOR2_X1 U641 ( .A1(n704), .A2(n542), .ZN(n539) );
  XNOR2_X1 U642 ( .A(KEYINPUT42), .B(n539), .ZN(n756) );
  XNOR2_X1 U643 ( .A(n540), .B(KEYINPUT46), .ZN(n568) );
  INV_X1 U644 ( .A(n374), .ZN(n543) );
  NOR2_X1 U645 ( .A1(n543), .A2(n542), .ZN(n652) );
  NOR2_X1 U646 ( .A1(n544), .A2(n557), .ZN(n649) );
  XNOR2_X1 U647 ( .A(KEYINPUT95), .B(n649), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n655), .A2(n578), .ZN(n617) );
  AND2_X1 U649 ( .A1(n652), .A2(n617), .ZN(n545) );
  NAND2_X1 U650 ( .A1(KEYINPUT70), .A2(n545), .ZN(n546) );
  XNOR2_X1 U651 ( .A(KEYINPUT47), .B(n546), .ZN(n566) );
  XNOR2_X1 U652 ( .A(n678), .B(KEYINPUT96), .ZN(n548) );
  INV_X1 U653 ( .A(KEYINPUT6), .ZN(n547) );
  XNOR2_X1 U654 ( .A(n548), .B(n547), .ZN(n621) );
  OR2_X1 U655 ( .A1(n552), .A2(n427), .ZN(n663) );
  NOR2_X1 U656 ( .A1(n554), .A2(n553), .ZN(n560) );
  INV_X1 U657 ( .A(n555), .ZN(n575) );
  NAND2_X1 U658 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U659 ( .A(n558), .B(KEYINPUT100), .ZN(n580) );
  NOR2_X1 U660 ( .A1(n575), .A2(n580), .ZN(n559) );
  NAND2_X1 U661 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U662 ( .A(KEYINPUT103), .B(n561), .ZN(n752) );
  INV_X1 U663 ( .A(n617), .ZN(n691) );
  NAND2_X1 U664 ( .A1(n652), .A2(n691), .ZN(n562) );
  NOR2_X1 U665 ( .A1(KEYINPUT70), .A2(n562), .ZN(n563) );
  NOR2_X1 U666 ( .A1(n752), .A2(n563), .ZN(n564) );
  NAND2_X1 U667 ( .A1(n663), .A2(n564), .ZN(n565) );
  NOR2_X1 U668 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U669 ( .A1(n568), .A2(n567), .ZN(n570) );
  INV_X1 U670 ( .A(n686), .ZN(n572) );
  NOR2_X1 U671 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U672 ( .A1(n427), .A2(n573), .ZN(n574) );
  XNOR2_X1 U673 ( .A(n574), .B(KEYINPUT43), .ZN(n576) );
  NAND2_X1 U674 ( .A1(n576), .A2(n575), .ZN(n667) );
  NOR2_X1 U675 ( .A1(n579), .A2(n578), .ZN(n666) );
  INV_X1 U676 ( .A(n580), .ZN(n592) );
  XNOR2_X1 U677 ( .A(n581), .B(KEYINPUT72), .ZN(n610) );
  NOR2_X1 U678 ( .A1(n610), .A2(n621), .ZN(n583) );
  OR2_X1 U679 ( .A1(G898), .A2(n741), .ZN(n729) );
  OR2_X1 U680 ( .A1(n729), .A2(n584), .ZN(n585) );
  NAND2_X1 U681 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U682 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n589) );
  XNOR2_X1 U683 ( .A(n611), .B(KEYINPUT88), .ZN(n614) );
  NOR2_X1 U684 ( .A1(n703), .A2(n614), .ZN(n590) );
  XNOR2_X1 U685 ( .A(n590), .B(KEYINPUT34), .ZN(n591) );
  XNOR2_X1 U686 ( .A(KEYINPUT75), .B(n621), .ZN(n599) );
  NOR2_X1 U687 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U688 ( .A1(n601), .A2(n355), .ZN(n603) );
  NOR2_X1 U689 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U690 ( .A(n604), .B(KEYINPUT32), .ZN(n758) );
  NAND2_X1 U691 ( .A1(n751), .A2(n608), .ZN(n605) );
  XNOR2_X1 U692 ( .A(n605), .B(KEYINPUT44), .ZN(n607) );
  INV_X1 U693 ( .A(KEYINPUT79), .ZN(n606) );
  NAND2_X1 U694 ( .A1(n607), .A2(n606), .ZN(n628) );
  NAND2_X1 U695 ( .A1(n609), .A2(KEYINPUT79), .ZN(n624) );
  OR2_X1 U696 ( .A1(n610), .A2(n678), .ZN(n681) );
  NOR2_X1 U697 ( .A1(n681), .A2(n611), .ZN(n612) );
  XNOR2_X1 U698 ( .A(n612), .B(KEYINPUT31), .ZN(n659) );
  NOR2_X1 U699 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U700 ( .A1(n615), .A2(n678), .ZN(n643) );
  NAND2_X1 U701 ( .A1(n659), .A2(n643), .ZN(n616) );
  XNOR2_X1 U702 ( .A(n616), .B(KEYINPUT90), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n618), .A2(n617), .ZN(n622) );
  NOR2_X1 U704 ( .A1(n668), .A2(n619), .ZN(n620) );
  NAND2_X1 U705 ( .A1(n621), .A2(n620), .ZN(n640) );
  AND2_X1 U706 ( .A1(n622), .A2(n640), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n626) );
  AND2_X1 U708 ( .A1(n751), .A2(KEYINPUT79), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  INV_X1 U710 ( .A(KEYINPUT2), .ZN(n631) );
  OR2_X1 U711 ( .A1(n631), .A2(n666), .ZN(n633) );
  XOR2_X1 U712 ( .A(KEYINPUT77), .B(n633), .Z(n634) );
  NOR2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U714 ( .A(KEYINPUT106), .B(KEYINPUT62), .Z(n638) );
  XNOR2_X1 U715 ( .A(G101), .B(n640), .ZN(G3) );
  NOR2_X1 U716 ( .A1(n655), .A2(n643), .ZN(n642) );
  XNOR2_X1 U717 ( .A(G104), .B(KEYINPUT107), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n642), .B(n641), .ZN(G6) );
  INV_X1 U719 ( .A(n649), .ZN(n660) );
  NOR2_X1 U720 ( .A1(n660), .A2(n643), .ZN(n648) );
  XOR2_X1 U721 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n645) );
  XNOR2_X1 U722 ( .A(G107), .B(KEYINPUT26), .ZN(n644) );
  XNOR2_X1 U723 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U724 ( .A(KEYINPUT108), .B(n646), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n648), .B(n647), .ZN(G9) );
  XOR2_X1 U726 ( .A(G128), .B(KEYINPUT29), .Z(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n649), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n651), .B(n650), .ZN(G30) );
  INV_X1 U729 ( .A(n655), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n654), .B(G146), .ZN(G48) );
  NOR2_X1 U732 ( .A1(n655), .A2(n659), .ZN(n657) );
  XNOR2_X1 U733 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n656) );
  XNOR2_X1 U734 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U735 ( .A(G113), .B(n658), .ZN(G15) );
  NOR2_X1 U736 ( .A1(n660), .A2(n659), .ZN(n662) );
  XNOR2_X1 U737 ( .A(G116), .B(KEYINPUT113), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n662), .B(n661), .ZN(G18) );
  INV_X1 U739 ( .A(n663), .ZN(n664) );
  XNOR2_X1 U740 ( .A(G125), .B(n664), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U742 ( .A(G134), .B(n666), .Z(G36) );
  XNOR2_X1 U743 ( .A(G140), .B(n667), .ZN(G42) );
  XOR2_X1 U744 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n671) );
  NAND2_X1 U745 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U746 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U747 ( .A(KEYINPUT114), .B(n672), .ZN(n677) );
  NOR2_X1 U748 ( .A1(n674), .A2(n355), .ZN(n675) );
  XNOR2_X1 U749 ( .A(KEYINPUT50), .B(n675), .ZN(n676) );
  NOR2_X1 U750 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U753 ( .A(KEYINPUT51), .B(n682), .ZN(n683) );
  NOR2_X1 U754 ( .A1(n704), .A2(n683), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n684), .B(KEYINPUT116), .ZN(n697) );
  NOR2_X1 U756 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U757 ( .A(KEYINPUT117), .B(n687), .Z(n688) );
  NOR2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n692), .B(KEYINPUT118), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U762 ( .A1(n703), .A2(n695), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U764 ( .A(n698), .B(KEYINPUT119), .Z(n699) );
  XNOR2_X1 U765 ( .A(KEYINPUT52), .B(n699), .ZN(n700) );
  NOR2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U767 ( .A(n702), .B(KEYINPUT120), .ZN(n706) );
  NOR2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n711) );
  NAND2_X1 U770 ( .A1(n707), .A2(n631), .ZN(n709) );
  NAND2_X1 U771 ( .A1(n709), .A2(n373), .ZN(n710) );
  NAND2_X1 U772 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U773 ( .A1(n712), .A2(G953), .ZN(n713) );
  XNOR2_X1 U774 ( .A(n713), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U775 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n716) );
  XNOR2_X1 U776 ( .A(n714), .B(KEYINPUT80), .ZN(n715) );
  XOR2_X1 U777 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n719) );
  XNOR2_X1 U778 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U779 ( .A1(n728), .A2(n727), .ZN(G66) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U782 ( .A1(n731), .A2(G898), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n732), .B(KEYINPUT123), .ZN(n735) );
  NOR2_X1 U784 ( .A1(n733), .A2(G953), .ZN(n734) );
  NOR2_X1 U785 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n737), .B(n736), .ZN(G69) );
  XOR2_X1 U787 ( .A(n738), .B(n739), .Z(n744) );
  XOR2_X1 U788 ( .A(n744), .B(n740), .Z(n742) );
  NAND2_X1 U789 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n743), .B(KEYINPUT124), .ZN(n749) );
  XNOR2_X1 U791 ( .A(G227), .B(n744), .ZN(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U793 ( .A1(n746), .A2(G953), .ZN(n747) );
  XOR2_X1 U794 ( .A(KEYINPUT125), .B(n747), .Z(n748) );
  NAND2_X1 U795 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U796 ( .A(n750), .B(KEYINPUT126), .ZN(G72) );
  XNOR2_X1 U797 ( .A(n751), .B(G122), .ZN(G24) );
  XOR2_X1 U798 ( .A(G143), .B(n752), .Z(G45) );
  XOR2_X1 U799 ( .A(n753), .B(G110), .Z(n754) );
  XNOR2_X1 U800 ( .A(KEYINPUT110), .B(n754), .ZN(G12) );
  XOR2_X1 U801 ( .A(n755), .B(G131), .Z(G33) );
  XNOR2_X1 U802 ( .A(G137), .B(KEYINPUT127), .ZN(n757) );
  XNOR2_X1 U803 ( .A(n757), .B(n756), .ZN(G39) );
  XOR2_X1 U804 ( .A(G119), .B(n758), .Z(G21) );
endmodule

