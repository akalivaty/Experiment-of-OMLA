//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n215), .B(new_n216), .C1(new_n202), .C2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n207), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n201), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n214), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT0), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n214), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n212), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n206), .A2(new_n207), .ZN(new_n235));
  AOI22_X1  g0035(.A1(new_n228), .A2(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n236), .B1(new_n228), .B2(new_n230), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n227), .A2(new_n238), .ZN(G361));
  XOR2_X1   g0039(.A(G238), .B(G244), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G264), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n247), .B(G270), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G358));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n207), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n201), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n252), .B(new_n255), .Z(G351));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n217), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT3), .B(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(G232), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G226), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G97), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n258), .ZN(new_n271));
  AOI211_X1 g0071(.A(new_n261), .B(new_n263), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT13), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT75), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n273), .A2(G179), .B1(new_n274), .B2(KEYINPUT14), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n273), .A2(new_n276), .B1(new_n274), .B2(KEYINPUT14), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n272), .B(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n274), .A2(KEYINPUT14), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G169), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n275), .A2(new_n277), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n283), .A2(new_n231), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT72), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n286), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(new_n231), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT72), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n211), .A2(G20), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G68), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n296), .A2(new_n207), .B1(new_n212), .B2(G68), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n212), .A2(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n221), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n289), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT11), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n288), .A2(new_n202), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT12), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n294), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT74), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n282), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n279), .A2(G200), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n273), .A2(G190), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n310), .B(new_n311), .C1(new_n306), .C2(new_n307), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n293), .A2(G77), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n288), .A2(new_n221), .ZN(new_n314));
  XOR2_X1   g0114(.A(KEYINPUT15), .B(G87), .Z(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(new_n298), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n318), .A2(new_n296), .B1(new_n212), .B2(new_n221), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n289), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n313), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT73), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n260), .A2(new_n222), .ZN(new_n324));
  OR3_X1    g0124(.A1(new_n324), .A2(KEYINPUT71), .A3(new_n263), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n265), .A2(G232), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n264), .B(new_n326), .C1(new_n217), .C2(new_n265), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n271), .C1(G107), .C2(new_n264), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT71), .B1(new_n324), .B2(new_n263), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G200), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n313), .A2(KEYINPUT73), .A3(new_n314), .A4(new_n320), .ZN(new_n332));
  INV_X1    g0132(.A(G190), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n323), .A2(new_n331), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n309), .A2(new_n312), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n288), .A2(new_n289), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G50), .A3(new_n292), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n318), .B(KEYINPUT69), .ZN(new_n339));
  INV_X1    g0139(.A(G150), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n339), .A2(new_n298), .B1(new_n340), .B2(new_n296), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(G20), .B2(new_n208), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n338), .B1(G50), .B2(new_n286), .C1(new_n342), .C2(new_n284), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n265), .A2(G222), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G223), .A2(G1698), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n264), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(new_n271), .C1(G77), .C2(new_n264), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n259), .A2(new_n262), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n347), .B(new_n348), .C1(new_n220), .C2(new_n260), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT70), .B(G179), .Z(new_n350));
  OR2_X1    g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n276), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n343), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(G200), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT9), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n355), .B1(new_n333), .B2(new_n349), .C1(new_n343), .C2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n343), .A2(new_n356), .ZN(new_n358));
  OR3_X1    g0158(.A1(new_n357), .A2(KEYINPUT10), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT10), .B1(new_n357), .B2(new_n358), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n354), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(KEYINPUT3), .A2(G33), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT7), .B1(new_n364), .B2(new_n212), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NOR4_X1   g0166(.A1(new_n362), .A2(new_n363), .A3(new_n366), .A4(G20), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n295), .A2(G159), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n203), .A2(new_n205), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G20), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT76), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n374), .A3(G20), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n368), .A2(new_n369), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT16), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n371), .A2(new_n374), .A3(G20), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n374), .B1(new_n371), .B2(G20), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n368), .A4(new_n369), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(new_n382), .A3(new_n289), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n220), .A2(G1698), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n384), .B1(G223), .B2(G1698), .C1(new_n362), .C2(new_n363), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G87), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n271), .ZN(new_n388));
  INV_X1    g0188(.A(new_n260), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n263), .B1(new_n389), .B2(G232), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n333), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT77), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n390), .ZN(new_n393));
  INV_X1    g0193(.A(G200), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n258), .B1(new_n385), .B2(new_n386), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n348), .B1(new_n260), .B2(new_n224), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT77), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n399), .A3(new_n333), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n392), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n339), .A2(new_n288), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n339), .B1(new_n211), .B2(G20), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n337), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n383), .A2(new_n401), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n383), .A2(new_n402), .A3(new_n404), .ZN(new_n408));
  INV_X1    g0208(.A(new_n350), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n398), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n393), .A2(new_n276), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n408), .A2(KEYINPUT18), .A3(new_n410), .A4(new_n411), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n407), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT78), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n415), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n405), .B(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT78), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n330), .A2(new_n350), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n323), .A2(new_n332), .B1(new_n276), .B2(new_n330), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n420), .A2(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AND4_X1   g0224(.A1(new_n336), .A2(new_n361), .A3(new_n417), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT90), .ZN(new_n427));
  INV_X1    g0227(.A(G45), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G1), .ZN(new_n429));
  AND2_X1   g0229(.A1(KEYINPUT5), .A2(G41), .ZN(new_n430));
  NOR2_X1   g0230(.A1(KEYINPUT5), .A2(G41), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G264), .A3(new_n258), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G250), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(G1698), .ZN(new_n436));
  AND2_X1   g0236(.A1(G257), .A2(G1698), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n436), .A2(new_n437), .B1(new_n362), .B2(new_n363), .ZN(new_n438));
  INV_X1    g0238(.A(G294), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n268), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n258), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n427), .B1(new_n434), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G257), .A2(G1698), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n435), .B2(G1698), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n440), .B1(new_n264), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n433), .B(KEYINPUT90), .C1(new_n446), .C2(new_n258), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT5), .B(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(G274), .A3(new_n429), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n448), .A2(KEYINPUT91), .A3(G179), .A4(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n443), .A2(G179), .A3(new_n450), .A4(new_n447), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT91), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n433), .B(new_n450), .C1(new_n446), .C2(new_n258), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G169), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n211), .A2(G33), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n337), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G107), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT25), .B1(new_n288), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n461), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n460), .A2(G107), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(KEYINPUT89), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n212), .B(G87), .C1(new_n362), .C2(new_n363), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT22), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT22), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n264), .A2(new_n470), .A3(new_n212), .A4(G87), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G116), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G20), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n212), .A2(G107), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT23), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n472), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(KEYINPUT89), .A3(new_n466), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n474), .B1(new_n469), .B2(new_n471), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n466), .A2(KEYINPUT89), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n477), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n467), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n465), .B1(new_n483), .B2(new_n284), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n457), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n465), .ZN(new_n486));
  INV_X1    g0286(.A(new_n467), .ZN(new_n487));
  AND4_X1   g0287(.A1(new_n481), .A2(new_n472), .A3(new_n475), .A4(new_n477), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n481), .B1(new_n480), .B2(new_n477), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n486), .B1(new_n490), .B2(new_n289), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n443), .A2(new_n450), .A3(new_n447), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n394), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(G190), .B2(new_n455), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n485), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(new_n212), .C1(G33), .C2(new_n269), .ZN(new_n498));
  INV_X1    g0298(.A(G116), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G20), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n289), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT88), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(KEYINPUT20), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(KEYINPUT20), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n498), .A2(new_n503), .A3(new_n289), .A4(new_n500), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n288), .A2(new_n499), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n458), .A2(G116), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n510), .B1(new_n291), .B2(new_n512), .ZN(new_n513));
  AOI211_X1 g0313(.A(KEYINPUT87), .B(new_n511), .C1(new_n287), .C2(new_n290), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n265), .A2(G257), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G264), .A2(G1698), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n264), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G303), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n364), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n520), .A3(new_n271), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n432), .A2(G270), .A3(new_n258), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n450), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n515), .A2(G169), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n513), .A2(new_n514), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n523), .A2(G200), .ZN(new_n528));
  INV_X1    g0328(.A(new_n523), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G190), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n527), .A2(new_n509), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n515), .A2(G179), .A3(new_n529), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n515), .A2(KEYINPUT21), .A3(G169), .A4(new_n523), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n526), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n298), .B2(new_n269), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT86), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n264), .A2(new_n212), .A3(G68), .ZN(new_n539));
  NAND3_X1  g0339(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n212), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  INV_X1    g0342(.A(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(KEYINPUT86), .B(new_n535), .C1(new_n298), .C2(new_n269), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n538), .A2(new_n539), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n289), .B1(new_n288), .B2(new_n316), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n460), .A2(new_n315), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n435), .B1(new_n428), .B2(G1), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n211), .A2(new_n262), .A3(G45), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n258), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n222), .A2(G1698), .ZN(new_n553));
  OAI221_X1 g0353(.A(new_n553), .B1(G238), .B2(G1698), .C1(new_n362), .C2(new_n363), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n473), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n555), .B2(new_n271), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n548), .A2(new_n549), .B1(new_n557), .B2(new_n276), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT85), .B1(new_n556), .B2(new_n409), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n258), .B1(new_n554), .B2(new_n473), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT85), .ZN(new_n561));
  NOR4_X1   g0361(.A1(new_n560), .A2(new_n561), .A3(new_n552), .A4(new_n350), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(G200), .B1(new_n560), .B2(new_n552), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n460), .A2(G87), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n547), .A2(new_n289), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n316), .A2(new_n288), .ZN(new_n567));
  AND4_X1   g0367(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n556), .A2(G190), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n558), .A2(new_n563), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n534), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(G244), .B(new_n265), .C1(new_n362), .C2(new_n363), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT4), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .A4(new_n265), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(G250), .A2(G1698), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n362), .B2(new_n363), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT81), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(KEYINPUT81), .B(new_n578), .C1(new_n362), .C2(new_n363), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n581), .A2(new_n582), .B1(G33), .B2(G283), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n258), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n231), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n449), .A2(new_n429), .B1(new_n585), .B2(new_n257), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT82), .B1(new_n586), .B2(G257), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n432), .A2(KEYINPUT82), .A3(G257), .A4(new_n258), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n450), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT83), .B1(new_n591), .B2(new_n394), .ZN(new_n592));
  OR3_X1    g0392(.A1(new_n286), .A2(KEYINPUT80), .A3(G97), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT80), .B1(new_n286), .B2(G97), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n459), .B2(new_n269), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n269), .A2(new_n461), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(new_n542), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n597), .A2(new_n269), .A3(G107), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n212), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n296), .A2(new_n221), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT79), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(G107), .B1(new_n365), .B2(new_n367), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT79), .ZN(new_n606));
  INV_X1    g0406(.A(new_n603), .ZN(new_n607));
  XNOR2_X1  g0407(.A(G97), .B(G107), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n600), .B1(new_n597), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n606), .B(new_n607), .C1(new_n609), .C2(new_n212), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n604), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n596), .B1(new_n611), .B2(new_n289), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT81), .B1(new_n264), .B2(new_n578), .ZN(new_n613));
  INV_X1    g0413(.A(new_n582), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n497), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n575), .A2(new_n576), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n271), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n450), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n432), .A2(G257), .A3(new_n258), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT82), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n621), .B2(new_n588), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(G190), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n617), .A2(new_n622), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT83), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n625), .A3(G200), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n592), .A2(new_n612), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT84), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n611), .A2(new_n289), .ZN(new_n629));
  INV_X1    g0429(.A(new_n596), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n617), .A2(new_n409), .A3(new_n622), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n624), .A2(new_n276), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n628), .B1(new_n627), .B2(new_n634), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n496), .B(new_n572), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n426), .A2(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n312), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n423), .A2(new_n422), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n309), .B2(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n641), .A2(new_n419), .B1(new_n414), .B2(new_n415), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n359), .A2(new_n360), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n353), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n548), .A2(new_n549), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n557), .A2(new_n276), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n556), .A2(new_n409), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n569), .A2(new_n548), .A3(new_n564), .A4(new_n565), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n650), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n452), .B(KEYINPUT91), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n491), .B1(new_n656), .B2(new_n456), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n526), .A2(new_n532), .A3(new_n533), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n627), .A2(new_n495), .A3(new_n652), .A4(new_n634), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n649), .B(new_n655), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n651), .B1(new_n650), .B2(new_n570), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n645), .B1(new_n426), .B2(new_n663), .ZN(G369));
  INV_X1    g0464(.A(G13), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G20), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n231), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT92), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT27), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(G213), .B1(new_n667), .B2(KEYINPUT27), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT92), .B1(new_n667), .B2(KEYINPUT27), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G343), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n515), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT93), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n658), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n534), .B2(new_n678), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n681), .A2(KEYINPUT94), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT94), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n680), .B2(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n496), .B1(new_n491), .B2(new_n675), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n657), .A2(new_n676), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n658), .A2(new_n675), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n496), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n657), .A2(new_n675), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n691), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n229), .ZN(new_n697));
  OR3_X1    g0497(.A1(new_n697), .A2(KEYINPUT95), .A3(G41), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT95), .B1(new_n697), .B2(G41), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n544), .A2(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n235), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(new_n700), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n612), .A2(new_n623), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n625), .B1(new_n624), .B2(G200), .ZN(new_n707));
  AOI211_X1 g0507(.A(KEYINPUT83), .B(new_n394), .C1(new_n617), .C2(new_n622), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT84), .B1(new_n709), .B2(new_n650), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n572), .A3(new_n496), .A4(new_n675), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n617), .A2(new_n443), .A3(new_n622), .A4(new_n447), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n529), .A2(G179), .A3(new_n556), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n521), .A2(G179), .A3(new_n450), .A4(new_n522), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n557), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n591), .A2(KEYINPUT30), .A3(new_n719), .A4(new_n448), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n529), .A2(new_n350), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n624), .A3(new_n557), .A4(new_n492), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n723), .B2(new_n676), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT97), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n717), .A2(KEYINPUT96), .A3(new_n722), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n720), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT96), .B1(new_n717), .B2(new_n722), .ZN(new_n729));
  OAI211_X1 g0529(.A(KEYINPUT31), .B(new_n676), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n713), .A2(new_n726), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n734), .B(new_n675), .C1(new_n661), .C2(new_n662), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT26), .B1(new_n634), .B2(new_n653), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n629), .A2(new_n630), .B1(new_n624), .B2(new_n276), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n570), .A2(new_n651), .A3(new_n632), .A4(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n739), .B(new_n649), .C1(new_n659), .C2(new_n660), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n740), .A2(new_n675), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n735), .B1(new_n741), .B2(new_n734), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n733), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n705), .B1(new_n743), .B2(G1), .ZN(G364));
  OR3_X1    g0544(.A1(KEYINPUT98), .A2(G13), .A3(G33), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT98), .B1(G13), .B2(G33), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n231), .B1(G20), .B2(new_n276), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n252), .A2(G45), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n697), .A2(new_n264), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n235), .B2(new_n428), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n751), .A2(new_n754), .B1(new_n499), .B2(new_n697), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n229), .A2(G355), .A3(new_n264), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n749), .B(new_n750), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n700), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n211), .B1(new_n666), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n212), .A2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(G179), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(new_n764), .A3(new_n394), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT100), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n264), .B1(new_n770), .B2(G329), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n333), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n212), .ZN(new_n773));
  INV_X1    g0573(.A(G326), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n212), .A2(new_n333), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n350), .A2(G200), .A3(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n771), .B1(new_n439), .B2(new_n773), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n350), .A2(new_n763), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n394), .A2(G179), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n775), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n519), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n763), .A2(new_n783), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR4_X1   g0588(.A1(new_n777), .A2(new_n782), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G322), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n350), .A2(new_n394), .A3(new_n775), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(KEYINPUT99), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT99), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n350), .A2(new_n793), .A3(new_n394), .A4(new_n775), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n778), .A2(new_n394), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT33), .B(G317), .Z(new_n798));
  OAI221_X1 g0598(.A(new_n789), .B1(new_n790), .B2(new_n795), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT103), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n780), .A2(new_n221), .B1(new_n461), .B2(new_n786), .ZN(new_n801));
  INV_X1    g0601(.A(new_n773), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n796), .A2(G68), .B1(G97), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT102), .ZN(new_n804));
  INV_X1    g0604(.A(new_n795), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n801), .B(new_n804), .C1(G58), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n769), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n806), .B(new_n809), .C1(new_n207), .C2(new_n776), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n264), .B1(new_n784), .B2(new_n543), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT101), .Z(new_n812));
  OAI21_X1  g0612(.A(new_n800), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n757), .B(new_n762), .C1(new_n813), .C2(new_n750), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n749), .B(KEYINPUT104), .Z(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n680), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n686), .B(new_n762), .C1(G330), .C2(new_n680), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  OAI22_X1  g0620(.A1(new_n795), .A2(new_n439), .B1(new_n269), .B2(new_n773), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT105), .Z(new_n822));
  OAI21_X1  g0622(.A(new_n364), .B1(new_n769), .B2(new_n781), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n784), .A2(new_n461), .B1(new_n786), .B2(new_n543), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n825), .B1(new_n499), .B2(new_n780), .C1(new_n519), .C2(new_n776), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G283), .B2(new_n796), .ZN(new_n827));
  INV_X1    g0627(.A(new_n776), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G150), .A2(new_n796), .B1(new_n828), .B2(G137), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n807), .B2(new_n780), .C1(new_n795), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT106), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT34), .Z(new_n833));
  NOR2_X1   g0633(.A1(new_n784), .A2(new_n207), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n773), .A2(new_n201), .B1(new_n202), .B2(new_n786), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n264), .B1(new_n769), .B2(new_n836), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n750), .B1(new_n827), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n761), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n747), .A2(new_n750), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n221), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n323), .A2(new_n332), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n676), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(new_n335), .B1(new_n423), .B2(new_n422), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n423), .A2(new_n422), .A3(new_n675), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n842), .B1(new_n748), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n848), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n663), .B2(new_n676), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n675), .B(new_n848), .C1(new_n661), .C2(new_n662), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(new_n733), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n762), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n849), .A2(new_n855), .ZN(G384));
  INV_X1    g0656(.A(KEYINPUT39), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n408), .A2(new_n674), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n418), .B2(new_n419), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n412), .A2(new_n858), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  INV_X1    g0661(.A(new_n405), .ZN(new_n862));
  NOR4_X1   g0662(.A1(new_n860), .A2(KEYINPUT108), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT108), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT37), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n412), .A2(new_n405), .A3(new_n858), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n860), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n861), .B1(new_n858), .B2(KEYINPUT107), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n405), .A3(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n408), .A2(new_n674), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT107), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n867), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n877), .A2(new_n859), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n857), .B1(new_n869), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n309), .A2(new_n676), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n877), .B2(new_n859), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n420), .A2(new_n873), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n876), .A4(new_n872), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT39), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n880), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n308), .A2(new_n676), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n309), .A2(new_n312), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n282), .A2(new_n308), .A3(new_n676), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n846), .B2(new_n852), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n882), .A2(new_n884), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n418), .A2(new_n674), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n886), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n644), .B1(new_n742), .B2(new_n425), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n850), .B1(new_n888), .B2(new_n889), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT109), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n724), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI211_X1 g0703(.A(KEYINPUT109), .B(KEYINPUT31), .C1(new_n723), .C2(new_n676), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT110), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n905), .A2(new_n713), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(new_n905), .B2(new_n713), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n900), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n882), .A2(new_n884), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n899), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n870), .A2(new_n865), .A3(KEYINPUT37), .A4(new_n405), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n868), .B(new_n912), .C1(new_n416), .C2(new_n858), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n878), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n899), .B1(new_n914), .B2(new_n884), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n890), .A2(new_n848), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n637), .A2(new_n676), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n902), .A2(new_n901), .ZN(new_n918));
  INV_X1    g0718(.A(new_n724), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n904), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT110), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n905), .A2(new_n713), .A3(new_n906), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n916), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n915), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n911), .A2(new_n926), .A3(G330), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n924), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n425), .A2(new_n928), .A3(G330), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n893), .A3(new_n900), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(new_n899), .B1(new_n915), .B2(new_n925), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n425), .A3(new_n928), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n898), .B(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n211), .B2(new_n666), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT35), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n233), .B1(new_n937), .B2(new_n609), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(G116), .C1(new_n937), .C2(new_n609), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT36), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n235), .A2(G77), .A3(new_n370), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(G50), .B2(new_n202), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(G1), .A3(new_n665), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n936), .A2(new_n940), .A3(new_n943), .ZN(G367));
  OAI211_X1 g0744(.A(new_n627), .B(new_n634), .C1(new_n612), .C2(new_n675), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n650), .A2(new_n676), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n693), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT111), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n634), .B1(new_n945), .B2(new_n485), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n949), .A2(KEYINPUT42), .B1(new_n675), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n548), .A2(new_n565), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n676), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n654), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n649), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n954), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n961), .B1(new_n954), .B2(new_n962), .ZN(new_n965));
  INV_X1    g0765(.A(new_n691), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n964), .A2(new_n965), .B1(new_n966), .B2(new_n947), .ZN(new_n967));
  INV_X1    g0767(.A(new_n965), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n966), .A2(new_n947), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n963), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n695), .A2(new_n947), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT44), .Z(new_n973));
  NOR2_X1   g0773(.A1(new_n695), .A2(new_n947), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n691), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n683), .A2(KEYINPUT112), .A3(new_n685), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n689), .A2(new_n692), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT112), .B1(new_n683), .B2(new_n685), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n978), .A2(new_n693), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n693), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n982), .B(KEYINPUT112), .C1(new_n683), .C2(new_n685), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n743), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n743), .B1(new_n977), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n700), .B(KEYINPUT41), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n760), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n959), .A2(new_n816), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n802), .A2(G68), .ZN(new_n991));
  INV_X1    g0791(.A(G137), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n991), .B1(new_n201), .B2(new_n784), .C1(new_n769), .C2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n786), .A2(new_n221), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n780), .A2(new_n207), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n797), .A2(new_n807), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n264), .B1(new_n776), .B2(new_n830), .ZN(new_n997));
  OR4_X1    g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n993), .B(new_n998), .C1(G150), .C2(new_n805), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n805), .A2(G303), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n784), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n780), .B2(new_n787), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT46), .B1(new_n1001), .B2(G116), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n364), .B1(new_n786), .B2(new_n269), .C1(new_n773), .C2(new_n461), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(G311), .C2(new_n828), .ZN(new_n1006));
  INV_X1    g0806(.A(G317), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n769), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1003), .B(new_n1008), .C1(G294), .C2(new_n796), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n999), .B1(new_n1000), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT47), .Z(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n750), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n749), .A2(new_n750), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n229), .B2(new_n316), .C1(new_n248), .C2(new_n753), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n761), .A3(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n971), .A2(new_n989), .B1(new_n990), .B2(new_n1015), .ZN(G387));
  OAI21_X1  g0816(.A(KEYINPUT116), .B1(new_n984), .B2(new_n743), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n743), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT116), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1018), .A2(new_n981), .A3(new_n1019), .A4(new_n983), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n758), .A3(new_n985), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n690), .A2(new_n815), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n697), .A2(new_n461), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n229), .A2(new_n264), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n245), .A2(G45), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT113), .Z(new_n1026));
  OR3_X1    g0826(.A1(new_n318), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT50), .B1(new_n318), .B2(G50), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1027), .A2(new_n1028), .A3(new_n428), .A4(new_n701), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n202), .A2(new_n221), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n752), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT114), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1023), .B1(new_n701), .B2(new_n1024), .C1(new_n1026), .C2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n762), .B1(new_n1033), .B2(new_n1013), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G303), .A2(new_n779), .B1(new_n796), .B2(G311), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n790), .B2(new_n776), .C1(new_n795), .C2(new_n1007), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT115), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT48), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n787), .B2(new_n773), .C1(new_n439), .C2(new_n784), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT49), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n786), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n264), .B1(new_n1041), .B2(G116), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(new_n774), .C2(new_n769), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n264), .B1(new_n797), .B2(new_n339), .C1(new_n202), .C2(new_n780), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G150), .B2(new_n770), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n776), .A2(new_n807), .B1(new_n269), .B2(new_n786), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n316), .A2(new_n773), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1001), .A2(G77), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n805), .A2(G50), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1045), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n750), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1022), .B(new_n1034), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n984), .A2(new_n760), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1021), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(KEYINPUT117), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT117), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1021), .A2(new_n1054), .A3(new_n1058), .A4(new_n1055), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(G393));
  XOR2_X1   g0860(.A(new_n977), .B(KEYINPUT118), .Z(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n760), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n795), .A2(new_n781), .B1(new_n1007), .B2(new_n776), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT52), .Z(new_n1064));
  AOI211_X1 g0864(.A(new_n264), .B(new_n1064), .C1(G294), .C2(new_n779), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n519), .B2(new_n797), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n784), .A2(new_n787), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n773), .A2(new_n499), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n769), .A2(new_n790), .B1(new_n461), .B2(new_n786), .ZN(new_n1069));
  NOR4_X1   g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n795), .A2(new_n807), .B1(new_n340), .B2(new_n776), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT51), .Z(new_n1072));
  AOI211_X1 g0872(.A(new_n364), .B(new_n1072), .C1(G143), .C2(new_n770), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n221), .B2(new_n773), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n784), .A2(new_n202), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n780), .A2(new_n318), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n797), .A2(new_n207), .B1(new_n543), .B2(new_n786), .ZN(new_n1077));
  NOR4_X1   g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n750), .B1(new_n1070), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1013), .B1(new_n269), .B2(new_n229), .C1(new_n753), .C2(new_n255), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n762), .B1(new_n947), .B2(new_n749), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n700), .B1(new_n977), .B2(new_n985), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n977), .B2(new_n985), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1062), .A2(new_n1082), .A3(new_n1084), .ZN(G390));
  OAI211_X1 g0885(.A(G330), .B(new_n848), .C1(new_n907), .C2(new_n908), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n891), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n845), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n740), .A2(new_n675), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n846), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  AND4_X1   g0891(.A1(G330), .A2(new_n731), .A3(new_n848), .A4(new_n890), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1087), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n891), .B1(new_n732), .B2(new_n850), .ZN(new_n1095));
  OAI211_X1 g0895(.A(G330), .B(new_n900), .C1(new_n907), .C2(new_n908), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n852), .A2(new_n846), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n897), .A2(new_n929), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n881), .B1(new_n1098), .B2(new_n890), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n880), .B2(new_n885), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n914), .A2(new_n884), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1090), .A2(new_n890), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n881), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1096), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT39), .B1(new_n914), .B2(new_n884), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT39), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1111), .A2(new_n1112), .B1(new_n892), .B2(new_n881), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n1092), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1103), .A2(new_n1110), .A3(new_n1115), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1105), .A2(new_n1109), .A3(new_n1093), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1096), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1102), .B(new_n1100), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1116), .A2(new_n758), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n760), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n747), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  INV_X1    g0925(.A(G125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n264), .B1(new_n776), .B2(new_n1125), .C1(new_n769), .C2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n802), .A2(G159), .B1(new_n1041), .B2(G50), .ZN(new_n1128));
  XOR2_X1   g0928(.A(KEYINPUT54), .B(G143), .Z(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1128), .B1(new_n797), .B2(new_n992), .C1(new_n780), .C2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1127), .B(new_n1131), .C1(G132), .C2(new_n805), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n784), .A2(new_n340), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT53), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n364), .B1(new_n784), .B2(new_n543), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT119), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n202), .B2(new_n786), .C1(new_n439), .C2(new_n769), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n780), .A2(new_n269), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n795), .A2(new_n499), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n776), .A2(new_n787), .B1(new_n221), .B2(new_n773), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n796), .A2(G107), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1132), .A2(new_n1134), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n761), .B1(new_n1143), .B2(new_n1053), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n339), .B2(new_n841), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1124), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1121), .A2(new_n1123), .A3(new_n1146), .ZN(G378));
  INV_X1    g0947(.A(new_n896), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1149));
  XNOR2_X1  g0949(.A(new_n361), .B(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n343), .A2(new_n674), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT120), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n927), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n932), .A2(KEYINPUT120), .A3(G330), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1153), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND4_X1   g0957(.A1(KEYINPUT120), .A2(new_n911), .A3(G330), .A4(new_n926), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1158), .A2(new_n1152), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1148), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT120), .B1(new_n932), .B2(G330), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1152), .B1(new_n1161), .B2(new_n1158), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1156), .A2(new_n1153), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n896), .A3(new_n1163), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1120), .A2(new_n1102), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT121), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT121), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1120), .A2(new_n1168), .A3(new_n1102), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1165), .A2(new_n1170), .A3(KEYINPUT57), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1168), .B1(new_n1120), .B2(new_n1102), .ZN(new_n1173));
  AOI211_X1 g0973(.A(KEYINPUT121), .B(new_n1101), .C1(new_n1122), .C2(new_n1100), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1172), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1171), .A2(new_n1177), .A3(new_n758), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n207), .B1(new_n362), .B2(G41), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1130), .A2(new_n784), .B1(new_n773), .B2(new_n340), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n776), .A2(new_n1126), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G137), .C2(new_n779), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n836), .B2(new_n797), .C1(new_n1125), .C2(new_n795), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT59), .ZN(new_n1185));
  AOI21_X1  g0985(.A(G33), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(G41), .B1(new_n770), .B2(G124), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n807), .C2(new_n786), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1179), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n786), .A2(new_n201), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n796), .A2(G97), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n828), .A2(G116), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n264), .A2(G41), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n991), .A4(new_n1194), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1191), .B(new_n1195), .C1(new_n315), .C2(new_n779), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n770), .A2(G283), .B1(G77), .B2(new_n1001), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n461), .C2(new_n795), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT58), .Z(new_n1199));
  OAI21_X1  g0999(.A(new_n750), .B1(new_n1190), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n762), .B1(new_n207), .B2(new_n841), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n1152), .C2(new_n748), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1165), .B2(new_n760), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1178), .A2(new_n1204), .ZN(G375));
  NAND3_X1  g1005(.A1(new_n1101), .A2(new_n1094), .A3(new_n1099), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1103), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(new_n987), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT122), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n759), .B(KEYINPUT123), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n891), .A2(new_n747), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n773), .A2(new_n207), .B1(new_n201), .B2(new_n786), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n364), .B1(new_n796), .B2(new_n1129), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n1125), .B2(new_n769), .C1(new_n836), .C2(new_n776), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1212), .B(new_n1214), .C1(G137), .C2(new_n805), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n340), .B2(new_n780), .C1(new_n807), .C2(new_n784), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n994), .B1(G97), .B2(new_n1001), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n316), .B2(new_n773), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n364), .B1(new_n439), .B2(new_n776), .C1(new_n780), .C2(new_n461), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G283), .C2(new_n805), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n499), .B2(new_n797), .C1(new_n519), .C2(new_n769), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1053), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n762), .B(new_n1222), .C1(new_n202), .C2(new_n841), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1100), .A2(new_n1210), .B1(new_n1211), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1209), .A2(new_n1224), .ZN(G381));
  NAND3_X1  g1025(.A1(new_n1057), .A2(new_n819), .A3(new_n1059), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(G384), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT124), .ZN(new_n1228));
  INV_X1    g1028(.A(G378), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1178), .A2(new_n1229), .A3(new_n1204), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1228), .A2(new_n1230), .A3(G387), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(G381), .A2(G390), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(G407));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1230), .ZN(G409));
  INV_X1    g1034(.A(KEYINPUT126), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G387), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1226), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n819), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(G393), .A2(G396), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(G387), .A3(new_n1226), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1239), .A2(G390), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G390), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1229), .B1(new_n1178), .B2(new_n1204), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT125), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n700), .B1(new_n1207), .B2(KEYINPUT60), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1092), .B1(new_n1086), .B2(new_n891), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1248), .A2(new_n1091), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT60), .B1(new_n1249), .B2(new_n1101), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1246), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1103), .B2(new_n1206), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(new_n1254), .A2(KEYINPUT125), .A3(new_n700), .A4(new_n1250), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1224), .B1(new_n1252), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G384), .B(new_n1224), .C1(new_n1252), .C2(new_n1255), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n988), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1210), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1176), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1263), .A2(G378), .A3(new_n1203), .ZN(new_n1264));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G343), .ZN(new_n1266));
  NOR4_X1   g1066(.A1(new_n1245), .A2(new_n1260), .A3(new_n1264), .A4(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1245), .A2(new_n1266), .A3(new_n1264), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(G2897), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1260), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1258), .A2(new_n1259), .A3(new_n1270), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n1267), .A2(new_n1268), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1266), .B1(G375), .B2(G378), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1264), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1276), .A2(new_n1268), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1244), .B1(new_n1275), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1280), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1267), .B2(KEYINPUT63), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G375), .A2(G378), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1266), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1288), .A3(new_n1278), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1285), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1284), .B1(new_n1290), .B2(new_n1267), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1282), .A2(new_n1291), .ZN(G405));
  INV_X1    g1092(.A(new_n1230), .ZN(new_n1293));
  OAI211_X1 g1093(.A(KEYINPUT127), .B(new_n1277), .C1(new_n1293), .C2(new_n1245), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1287), .B(new_n1230), .C1(new_n1295), .C2(new_n1260), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1244), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1297), .B(new_n1298), .ZN(G402));
endmodule


