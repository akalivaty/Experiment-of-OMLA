//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n206), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT1), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n209), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT64), .Z(new_n231));
  AOI21_X1  g0031(.A(new_n225), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  AND3_X1   g0032(.A1(new_n221), .A2(new_n222), .A3(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT67), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G68), .ZN(new_n247));
  INV_X1    g0047(.A(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n246), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n254), .A2(new_n227), .A3(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n226), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(G50), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n255), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(G50), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g0063(.A(KEYINPUT8), .B(G58), .Z(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n264), .A2(new_n266), .B1(G150), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n268), .A2(KEYINPUT69), .B1(G20), .B2(new_n203), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n263), .B1(new_n271), .B2(new_n257), .ZN(new_n272));
  XOR2_X1   g0072(.A(new_n272), .B(KEYINPUT9), .Z(new_n273));
  AND2_X1   g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT68), .B1(new_n274), .B2(new_n226), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(G1), .A4(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G226), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n274), .A2(new_n226), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(new_n211), .B2(new_n289), .ZN(new_n290));
  MUX2_X1   g0090(.A(G222), .B(G223), .S(G1698), .Z(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n275), .A2(new_n281), .A3(G274), .A4(new_n278), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n283), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(G200), .B2(new_n294), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n273), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n273), .A2(new_n300), .A3(new_n297), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT3), .B(G33), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(G238), .A3(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(G232), .A3(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n306), .C1(new_n206), .C2(new_n303), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n284), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n282), .A2(G244), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n308), .A2(new_n293), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n257), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n264), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  INV_X1    g0115(.A(new_n266), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n313), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n258), .A2(G77), .A3(new_n260), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n211), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT70), .B1(new_n255), .B2(new_n211), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n312), .B1(G169), .B2(new_n310), .C1(new_n319), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n310), .A2(G190), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n319), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n327), .C1(new_n328), .C2(new_n310), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n272), .B1(new_n332), .B2(new_n294), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n294), .A2(G179), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n302), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n258), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n264), .A2(new_n260), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n338), .A2(new_n339), .B1(new_n262), .B2(new_n264), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G58), .A2(G68), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n229), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(G20), .B1(G159), .B2(new_n267), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT74), .ZN(new_n344));
  AOI21_X1  g0144(.A(G20), .B1(new_n287), .B2(new_n288), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(KEYINPUT7), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT7), .ZN(new_n347));
  OAI211_X1 g0147(.A(KEYINPUT74), .B(new_n347), .C1(new_n303), .C2(G20), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(G20), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n287), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n286), .A2(KEYINPUT75), .A3(G33), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n288), .A3(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n346), .A2(new_n348), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n343), .B1(new_n354), .B2(new_n248), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n313), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n265), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT72), .B1(new_n265), .B2(KEYINPUT3), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n287), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT73), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(new_n349), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT72), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n286), .B2(G33), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n265), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n347), .B1(new_n367), .B2(G20), .ZN(new_n368));
  INV_X1    g0168(.A(new_n349), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT73), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n362), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G68), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(KEYINPUT16), .A3(new_n343), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n340), .B1(new_n357), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  INV_X1    g0175(.A(G226), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G1698), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G223), .B2(G1698), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n375), .B1(new_n360), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n284), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n275), .A2(G232), .A3(new_n280), .A4(new_n278), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n293), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT76), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G223), .A2(G1698), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n376), .B2(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n367), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n285), .B1(new_n387), .B2(new_n375), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n388), .A2(new_n382), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n328), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n388), .A2(new_n382), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n295), .A2(KEYINPUT77), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n295), .A2(KEYINPUT77), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n391), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n374), .A2(new_n397), .A3(KEYINPUT17), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT17), .B1(new_n374), .B2(new_n397), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n346), .A2(new_n348), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n353), .A2(new_n349), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n248), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n343), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n356), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n373), .A2(new_n405), .A3(new_n257), .ZN(new_n406));
  INV_X1    g0206(.A(new_n340), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n332), .B1(new_n384), .B2(new_n390), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n392), .A2(new_n311), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT18), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n409), .A2(new_n410), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n413), .B1(new_n374), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n400), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT71), .B1(new_n262), .B2(G68), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT12), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT11), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n266), .A2(G77), .B1(G20), .B2(new_n248), .ZN(new_n421));
  INV_X1    g0221(.A(new_n267), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n202), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n257), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n419), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n258), .A2(G68), .A3(new_n260), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n282), .A2(G238), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G97), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n376), .A2(new_n305), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(G232), .B2(new_n305), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n432), .B2(new_n289), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n284), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n293), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(KEYINPUT13), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(G169), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n311), .B2(new_n438), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n438), .B2(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n428), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n438), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n428), .B1(new_n444), .B2(G190), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n328), .B2(new_n444), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n337), .A2(new_n417), .A3(new_n447), .ZN(new_n448));
  MUX2_X1   g0248(.A(G250), .B(G257), .S(G1698), .Z(new_n449));
  AOI22_X1  g0249(.A1(new_n367), .A2(new_n449), .B1(G33), .B2(G294), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n450), .A2(new_n285), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n259), .A2(G45), .ZN(new_n452));
  OR2_X1    g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(G274), .A3(new_n275), .A4(new_n278), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n279), .A2(new_n455), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G264), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n451), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n295), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(KEYINPUT86), .C1(G200), .C2(new_n460), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n367), .A2(KEYINPUT22), .A3(new_n227), .A4(G87), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n464));
  OR3_X1    g0264(.A1(new_n227), .A2(KEYINPUT23), .A3(G107), .ZN(new_n465));
  NAND2_X1  g0265(.A1(KEYINPUT84), .A2(KEYINPUT24), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT23), .B1(new_n227), .B2(G107), .ZN(new_n467));
  AND4_X1   g0267(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n227), .A2(G87), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n289), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n463), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT84), .A2(KEYINPUT24), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n313), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n258), .B1(G1), .B2(new_n265), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT25), .B1(new_n255), .B2(new_n206), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n255), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n476), .A2(new_n206), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n462), .B(new_n480), .C1(KEYINPUT86), .C2(new_n461), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n460), .A2(G179), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n459), .A2(KEYINPUT85), .A3(G169), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT85), .B1(new_n459), .B2(G169), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n484), .A2(new_n485), .B1(new_n475), .B2(new_n479), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  XOR2_X1   g0288(.A(new_n488), .B(KEYINPUT80), .Z(new_n489));
  NAND4_X1  g0289(.A1(new_n303), .A2(KEYINPUT4), .A3(G244), .A4(new_n305), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n303), .A2(G250), .A3(G1698), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n305), .A2(G244), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n360), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT81), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n492), .A2(new_n495), .A3(KEYINPUT81), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n284), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n457), .A2(G257), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n501), .A2(new_n456), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G200), .ZN(new_n504));
  XOR2_X1   g0304(.A(KEYINPUT78), .B(G97), .Z(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n506), .A2(KEYINPUT6), .A3(new_n206), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT6), .B1(new_n207), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n510), .A2(new_n227), .B1(new_n211), .B2(new_n422), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n354), .A2(new_n206), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n257), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n255), .A2(new_n205), .ZN(new_n514));
  XOR2_X1   g0314(.A(new_n514), .B(KEYINPUT79), .Z(new_n515));
  INV_X1    g0315(.A(new_n476), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(G97), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n500), .A2(G190), .A3(new_n502), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n504), .A2(new_n513), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n503), .A2(new_n332), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n500), .A2(new_n311), .A3(new_n502), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n513), .A2(new_n517), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n262), .A2(G116), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n516), .B2(G116), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n489), .B(new_n227), .C1(G33), .C2(new_n505), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n313), .B1(G20), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT20), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n455), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(G270), .A3(new_n275), .A4(new_n278), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G257), .A2(G1698), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n213), .B2(G1698), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n367), .A2(new_n539), .B1(G303), .B2(new_n289), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n456), .B(new_n537), .C1(new_n540), .C2(new_n285), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G200), .ZN(new_n542));
  INV_X1    g0342(.A(new_n396), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n535), .B(new_n542), .C1(new_n543), .C2(new_n541), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT21), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n541), .A2(G169), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n535), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n533), .A2(new_n534), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n526), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n541), .A2(new_n311), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n549), .A2(KEYINPUT21), .A3(G169), .A4(new_n541), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n544), .A2(new_n547), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n476), .A2(new_n315), .ZN(new_n554));
  XNOR2_X1  g0354(.A(new_n554), .B(KEYINPUT83), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n367), .A2(new_n227), .A3(G68), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n505), .B2(new_n316), .ZN(new_n558));
  INV_X1    g0358(.A(G87), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n505), .A2(new_n559), .A3(new_n206), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n227), .B1(new_n430), .B2(new_n557), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n561), .A2(new_n562), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n556), .B(new_n558), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(new_n257), .B1(new_n255), .B2(new_n315), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n555), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(G250), .B1(new_n259), .B2(G45), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n452), .A2(G274), .ZN(new_n570));
  OR3_X1    g0370(.A1(new_n279), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G238), .A2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n212), .B2(G1698), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n367), .A2(new_n573), .B1(G33), .B2(G116), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n571), .B1(new_n285), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G169), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n311), .B2(new_n575), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n568), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n575), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G190), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n575), .A2(G200), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n516), .A2(G87), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n567), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n553), .A2(new_n584), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n448), .A2(new_n487), .A3(new_n524), .A4(new_n585), .ZN(G372));
  OR2_X1    g0386(.A1(new_n325), .A2(KEYINPUT89), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n325), .A2(KEYINPUT89), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n443), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(new_n400), .A3(new_n446), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT88), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT18), .B1(new_n408), .B2(new_n411), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n374), .A2(new_n414), .A3(new_n413), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n412), .A2(new_n415), .A3(KEYINPUT88), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT90), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n302), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n299), .A2(KEYINPUT90), .A3(new_n301), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n335), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n486), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n547), .A2(new_n552), .A3(new_n551), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n481), .A2(new_n523), .A3(new_n519), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT87), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n584), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n578), .A2(KEYINPUT87), .A3(new_n583), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n605), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT26), .B1(new_n523), .B2(new_n584), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n608), .A3(new_n609), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n578), .B(new_n612), .C1(new_n614), .C2(KEYINPUT26), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n448), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n602), .A2(new_n617), .ZN(G369));
  NAND3_X1  g0418(.A1(new_n259), .A2(new_n227), .A3(G13), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(G213), .ZN(new_n622));
  INV_X1    g0422(.A(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n487), .B1(new_n480), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n486), .B2(new_n625), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n535), .A2(new_n625), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n604), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n553), .B2(new_n628), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(G330), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n486), .A2(new_n481), .A3(new_n604), .A4(new_n625), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n603), .B2(new_n625), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(G399));
  OR2_X1    g0436(.A1(new_n560), .A2(G116), .ZN(new_n637));
  INV_X1    g0437(.A(new_n223), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(G41), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G1), .ZN(new_n641));
  OAI22_X1  g0441(.A1(new_n637), .A2(new_n641), .B1(new_n230), .B2(new_n640), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n642), .B(KEYINPUT28), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n616), .A2(new_n625), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT29), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n614), .A2(KEYINPUT26), .ZN(new_n647));
  OR3_X1    g0447(.A1(new_n523), .A2(new_n584), .A3(KEYINPUT26), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n578), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT93), .B1(new_n603), .B2(new_n604), .ZN(new_n651));
  INV_X1    g0451(.A(new_n604), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT93), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n486), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n606), .A2(new_n610), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n624), .B1(new_n650), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT29), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n646), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n487), .A2(new_n524), .A3(new_n585), .A4(new_n625), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n460), .B1(new_n500), .B2(new_n502), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT91), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n579), .A2(G179), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n541), .B(new_n666), .C1(new_n662), .C2(new_n663), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT30), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n451), .A2(new_n458), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n575), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n500), .A2(new_n670), .A3(new_n502), .A4(new_n550), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n665), .A2(new_n667), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n668), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI211_X1 g0474(.A(KEYINPUT31), .B(new_n624), .C1(new_n672), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n666), .A2(new_n541), .ZN(new_n676));
  INV_X1    g0476(.A(new_n662), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(KEYINPUT91), .ZN(new_n678));
  INV_X1    g0478(.A(new_n671), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n678), .A2(new_n664), .B1(KEYINPUT30), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n673), .B(KEYINPUT92), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n625), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n661), .B(new_n675), .C1(new_n682), .C2(KEYINPUT31), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n660), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n643), .B1(new_n685), .B2(G1), .ZN(G364));
  NOR2_X1   g0486(.A1(new_n254), .A2(G20), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n259), .B1(new_n687), .B2(G45), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n639), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(G355), .A2(KEYINPUT94), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n638), .A2(new_n289), .ZN(new_n693));
  NAND2_X1  g0493(.A1(G355), .A2(KEYINPUT94), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n367), .A2(new_n638), .ZN(new_n696));
  INV_X1    g0496(.A(new_n231), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(G45), .ZN(new_n698));
  INV_X1    g0498(.A(G45), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n252), .A2(new_n699), .ZN(new_n700));
  OAI221_X1 g0500(.A(new_n695), .B1(G116), .B2(new_n223), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n254), .A2(new_n265), .A3(KEYINPUT95), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT95), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(G13), .B2(G33), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G20), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n226), .B1(G20), .B2(new_n332), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n691), .B1(new_n701), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n328), .A2(G179), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n712), .A2(new_n227), .A3(new_n295), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n289), .B1(new_n713), .B2(G87), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n227), .A2(new_n311), .A3(G200), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n715), .A2(new_n295), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n295), .A2(G20), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT96), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n712), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI221_X1 g0521(.A(new_n714), .B1(new_n717), .B2(new_n211), .C1(new_n721), .C2(new_n206), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n227), .A2(new_n311), .A3(new_n328), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n396), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n227), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n725), .A2(G50), .B1(new_n728), .B2(G97), .ZN(new_n729));
  INV_X1    g0529(.A(G58), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n396), .A2(new_n715), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n723), .A2(KEYINPUT97), .A3(new_n295), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT97), .B1(new_n723), .B2(new_n295), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n722), .B(new_n733), .C1(G68), .C2(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n719), .A2(G179), .A3(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G159), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT32), .Z(new_n741));
  XOR2_X1   g0541(.A(KEYINPUT33), .B(G317), .Z(new_n742));
  NOR2_X1   g0542(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G322), .ZN(new_n744));
  INV_X1    g0544(.A(G294), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n732), .A2(new_n744), .B1(new_n745), .B2(new_n727), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n743), .B(new_n746), .C1(G311), .C2(new_n716), .ZN(new_n747));
  INV_X1    g0547(.A(G283), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n721), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G326), .ZN(new_n750));
  INV_X1    g0550(.A(G303), .ZN(new_n751));
  INV_X1    g0551(.A(new_n713), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n289), .B1(new_n724), .B2(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n749), .B(new_n753), .C1(G329), .C2(new_n739), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n738), .A2(new_n741), .B1(new_n747), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n708), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n710), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT98), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n707), .B(KEYINPUT99), .Z(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n630), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n630), .A2(G330), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n631), .A2(new_n691), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(G396));
  NOR2_X1   g0563(.A1(new_n327), .A2(new_n625), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n587), .B2(new_n588), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n331), .A2(KEYINPUT102), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n330), .A2(KEYINPUT102), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n765), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n644), .A2(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n766), .A2(new_n767), .B1(new_n769), .B2(new_n765), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n625), .B(new_n773), .C1(new_n611), .C2(new_n615), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n691), .B1(new_n775), .B2(new_n684), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(KEYINPUT103), .B1(new_n684), .B2(new_n775), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(KEYINPUT103), .B2(new_n776), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n705), .A2(new_n708), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n691), .B1(new_n211), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n725), .A2(G137), .B1(new_n716), .B2(G159), .ZN(new_n781));
  INV_X1    g0581(.A(G143), .ZN(new_n782));
  INV_X1    g0582(.A(G150), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n781), .B1(new_n782), .B2(new_n732), .C1(new_n736), .C2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT34), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n367), .B1(new_n730), .B2(new_n727), .C1(new_n752), .C2(new_n202), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n721), .A2(new_n248), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(G132), .C2(new_n739), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n720), .A2(G87), .ZN(new_n790));
  INV_X1    g0590(.A(new_n739), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT100), .Z(new_n794));
  OAI221_X1 g0594(.A(new_n289), .B1(new_n205), .B2(new_n727), .C1(new_n752), .C2(new_n206), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n732), .A2(new_n745), .B1(new_n751), .B2(new_n724), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n795), .B(new_n796), .C1(G116), .C2(new_n716), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n748), .B2(new_n736), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n789), .B1(new_n794), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n800), .A2(KEYINPUT101), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n708), .B1(new_n800), .B2(KEYINPUT101), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n780), .B1(new_n773), .B2(new_n706), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n778), .A2(new_n803), .ZN(G384));
  INV_X1    g0604(.A(new_n510), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT35), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT35), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n806), .A2(G116), .A3(new_n228), .A4(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT36), .Z(new_n809));
  NAND4_X1  g0609(.A1(new_n229), .A2(G50), .A3(G77), .A4(new_n341), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n259), .B(G13), .C1(new_n810), .C2(new_n247), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n443), .A2(new_n624), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT107), .ZN(new_n815));
  INV_X1    g0615(.A(new_n622), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n408), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n374), .A2(new_n397), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n817), .A2(new_n818), .A3(new_n592), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n622), .B1(new_n406), .B2(new_n407), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n374), .B2(new_n397), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n374), .A2(new_n414), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(KEYINPUT37), .A2(new_n819), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n817), .A2(new_n818), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT37), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n825), .A2(new_n592), .A3(new_n826), .A4(new_n822), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n595), .A2(new_n400), .A3(new_n596), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n820), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT106), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n831), .A2(KEYINPUT106), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n826), .B1(new_n825), .B2(new_n822), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n373), .A2(new_n257), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT16), .B1(new_n372), .B2(new_n343), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n407), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n816), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n411), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT37), .A4(new_n818), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n843), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n417), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n846), .A2(new_n848), .A3(KEYINPUT38), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n815), .B1(new_n838), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT106), .B1(new_n831), .B2(new_n833), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n835), .B(new_n832), .C1(new_n828), .C2(new_n830), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n815), .B(new_n850), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT38), .B1(new_n846), .B2(new_n848), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n814), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n816), .B1(new_n595), .B2(new_n596), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n325), .A2(new_n624), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n774), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n428), .A2(new_n624), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT104), .Z(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n447), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n866), .A2(new_n443), .A3(new_n446), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n861), .B1(new_n857), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n860), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n646), .A2(new_n659), .A3(new_n448), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n602), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n874), .B(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n849), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n852), .B2(new_n853), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT92), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n673), .B(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT31), .B(new_n624), .C1(new_n881), .C2(new_n672), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n882), .B(new_n661), .C1(new_n682), .C2(KEYINPUT31), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n771), .B1(new_n869), .B2(new_n868), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n879), .A2(KEYINPUT40), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n883), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n856), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n448), .A2(new_n883), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(G330), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n877), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT108), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n895), .B1(new_n259), .B2(new_n687), .C1(new_n877), .C2(new_n893), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(KEYINPUT108), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n812), .B1(new_n896), .B2(new_n897), .ZN(G367));
  OAI21_X1  g0698(.A(new_n709), .B1(new_n223), .B2(new_n315), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n242), .B2(new_n696), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n731), .A2(G150), .B1(G68), .B2(new_n728), .ZN(new_n901));
  INV_X1    g0701(.A(G159), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n901), .B1(new_n202), .B2(new_n717), .C1(new_n902), .C2(new_n736), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n739), .A2(G137), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n725), .A2(G143), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n720), .A2(G77), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n289), .B1(new_n713), .B2(G58), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n713), .A2(G116), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT46), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n367), .B1(new_n731), .B2(G303), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n739), .A2(G317), .B1(new_n720), .B2(new_n506), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(G107), .A2(new_n728), .B1(new_n716), .B2(G283), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n914), .B1(new_n792), .B2(new_n724), .C1(new_n736), .C2(new_n745), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n903), .A2(new_n908), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT47), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n691), .B(new_n900), .C1(new_n917), .C2(new_n708), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n567), .A2(new_n582), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n624), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n608), .A2(new_n609), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n578), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n918), .B1(new_n922), .B2(new_n759), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT110), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n522), .A2(new_n624), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n524), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n613), .A2(new_n624), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n930), .A2(new_n634), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT42), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n524), .A2(new_n603), .A3(new_n927), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n624), .B1(new_n935), .B2(new_n523), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT109), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n926), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n633), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n930), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n924), .A2(new_n925), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n635), .A2(new_n930), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n635), .A2(new_n930), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n941), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT111), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT111), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n955), .A3(new_n941), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n948), .A2(new_n633), .A3(new_n951), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT112), .ZN(new_n959));
  INV_X1    g0759(.A(new_n634), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n604), .A2(new_n625), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n960), .B1(new_n627), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(new_n631), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n685), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n660), .A2(new_n684), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT112), .B1(new_n966), .B2(new_n963), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n685), .B1(new_n958), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n639), .B(KEYINPUT41), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n689), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n923), .B1(new_n946), .B2(new_n972), .ZN(G387));
  OAI211_X1 g0773(.A(new_n968), .B(new_n639), .C1(new_n685), .C2(new_n964), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n360), .B1(new_n791), .B2(new_n750), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G283), .A2(new_n728), .B1(new_n713), .B2(G294), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n731), .A2(G317), .B1(G303), .B2(new_n716), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n744), .B2(new_n724), .C1(new_n792), .C2(new_n736), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT113), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n976), .B1(new_n979), .B2(KEYINPUT48), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(KEYINPUT48), .B2(new_n979), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT49), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n975), .B(new_n982), .C1(G116), .C2(new_n720), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n713), .A2(G77), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n367), .B(new_n984), .C1(new_n791), .C2(new_n783), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G159), .A2(new_n725), .B1(new_n731), .B2(G50), .ZN(new_n986));
  INV_X1    g0786(.A(new_n315), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n987), .A2(new_n728), .B1(new_n716), .B2(G68), .ZN(new_n988));
  INV_X1    g0788(.A(new_n264), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n986), .B(new_n988), .C1(new_n989), .C2(new_n736), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n985), .B(new_n990), .C1(G97), .C2(new_n720), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n708), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n696), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n239), .B2(G45), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n637), .B2(new_n693), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n264), .A2(new_n202), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT50), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n699), .B1(new_n248), .B2(new_n211), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n997), .A2(new_n637), .A3(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n995), .A2(new_n999), .B1(G107), .B2(new_n223), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n691), .B1(new_n1000), .B2(new_n709), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n992), .B(new_n1001), .C1(new_n627), .C2(new_n759), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n974), .B(new_n1002), .C1(new_n688), .C2(new_n963), .ZN(G393));
  NAND2_X1  g0803(.A1(new_n953), .A2(new_n957), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n968), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1005), .B(new_n639), .C1(new_n968), .C2(new_n958), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1004), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n928), .A2(new_n707), .A3(new_n929), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n709), .B1(new_n223), .B2(new_n505), .C1(new_n246), .C2(new_n993), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n690), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n732), .A2(new_n902), .B1(new_n783), .B2(new_n724), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT114), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT51), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n790), .B1(new_n791), .B2(new_n782), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n367), .B1(new_n752), .B2(new_n248), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n728), .A2(G77), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n717), .B2(new_n989), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n202), .B2(new_n736), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G317), .A2(new_n725), .B1(new_n731), .B2(G311), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT115), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT52), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n303), .B1(new_n713), .B2(G283), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n529), .B2(new_n727), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G294), .B2(new_n716), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n739), .A2(G322), .B1(new_n720), .B2(G107), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n751), .C2(new_n736), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1013), .A2(new_n1019), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1010), .B1(new_n1028), .B2(new_n708), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1007), .A2(new_n689), .B1(new_n1008), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1006), .A2(new_n1030), .ZN(G390));
  NAND3_X1  g0831(.A1(new_n884), .A2(G330), .A3(new_n883), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT107), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n871), .A2(new_n813), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1034), .A2(new_n858), .A3(new_n854), .A4(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n655), .A2(new_n656), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n625), .B(new_n773), .C1(new_n1037), .C2(new_n649), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n863), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n814), .B1(new_n1039), .B2(new_n870), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n879), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1032), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n683), .A2(G330), .A3(new_n773), .A4(new_n870), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n1040), .B2(new_n879), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1036), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT116), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1036), .A2(new_n1045), .A3(KEYINPUT116), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1042), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1034), .A2(new_n705), .A3(new_n858), .A4(new_n854), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n691), .B1(new_n989), .B2(new_n779), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT119), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n303), .B1(new_n713), .B2(G87), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n1016), .C1(new_n721), .C2(new_n248), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n731), .A2(G116), .B1(new_n506), .B2(new_n716), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n748), .B2(new_n724), .C1(new_n206), .C2(new_n736), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1055), .B(new_n1057), .C1(G294), .C2(new_n739), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT121), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n727), .A2(new_n902), .ZN(new_n1062));
  INV_X1    g0862(.A(G128), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n303), .B1(new_n724), .B2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1062), .B(new_n1064), .C1(G132), .C2(new_n731), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT54), .B(G143), .Z(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT120), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1067), .A2(new_n716), .B1(new_n720), .B2(G50), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT53), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n752), .B2(new_n783), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n713), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1070), .A2(new_n1071), .B1(G125), .B2(new_n739), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n737), .A2(G137), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1065), .A2(new_n1068), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1060), .A2(new_n1061), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1053), .B1(new_n1075), .B2(new_n708), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1050), .A2(new_n689), .B1(new_n1051), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1032), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1036), .A2(new_n1045), .A3(KEYINPUT116), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT116), .B1(new_n1036), .B2(new_n1045), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT117), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n883), .A2(G330), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n870), .B1(new_n1085), .B2(new_n773), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1043), .A2(new_n863), .A3(new_n1038), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n870), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n883), .A2(G330), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n771), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n862), .B1(new_n658), .B2(new_n773), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT117), .A4(new_n1043), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n683), .A2(G330), .A3(new_n773), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1089), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1032), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n864), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1088), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1085), .A2(new_n448), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n875), .A2(new_n602), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(KEYINPUT118), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n639), .B1(new_n1083), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1050), .A2(new_n1103), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1077), .B1(new_n1105), .B2(new_n1106), .ZN(G378));
  AOI21_X1  g0907(.A(new_n1100), .B1(new_n1050), .B2(new_n1098), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n601), .A2(new_n336), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n272), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n1110), .A3(new_n816), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n601), .B(new_n336), .C1(new_n272), .C2(new_n622), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n849), .B1(new_n836), .B2(new_n837), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n884), .A2(KEYINPUT40), .A3(new_n883), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n888), .B(G330), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1118), .A2(new_n885), .A3(G330), .A4(new_n888), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n874), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1123), .A2(new_n1124), .B1(new_n860), .B2(new_n873), .ZN(new_n1127));
  OAI21_X1  g0927(.A(KEYINPUT57), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n639), .B1(new_n1108), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1080), .B(new_n1098), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1101), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1125), .B(new_n874), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT57), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n689), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G116), .A2(new_n725), .B1(new_n731), .B2(G107), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n315), .B2(new_n717), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n721), .A2(new_n730), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G283), .B2(new_n739), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n728), .A2(G68), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n367), .A2(G41), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n984), .A4(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1137), .B(new_n1142), .C1(G97), .C2(new_n737), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1143), .A2(KEYINPUT58), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(KEYINPUT58), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1145), .C1(new_n1141), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n737), .A2(G132), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n725), .A2(G125), .B1(new_n716), .B2(G137), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1067), .A2(new_n713), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n731), .A2(G128), .B1(G150), .B2(new_n728), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(G33), .A2(G41), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n721), .B2(new_n902), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G124), .B2(new_n739), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1153), .A2(new_n1154), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n708), .B1(new_n1147), .B2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT122), .Z(new_n1160));
  AOI21_X1  g0960(.A(new_n691), .B1(new_n202), .B2(new_n779), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n1118), .C2(new_n706), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1135), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1134), .A2(new_n1164), .ZN(G375));
  NOR2_X1   g0965(.A1(new_n870), .A2(new_n706), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n360), .B(new_n1138), .C1(G159), .C2(new_n713), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1063), .B2(new_n791), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n737), .A2(new_n1067), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G132), .A2(new_n725), .B1(new_n731), .B2(G137), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G50), .A2(new_n728), .B1(new_n716), .B2(G150), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n731), .A2(G283), .B1(G107), .B2(new_n716), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n745), .B2(new_n724), .C1(new_n529), .C2(new_n736), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n739), .A2(G303), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n728), .A2(new_n987), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n303), .B1(new_n713), .B2(G97), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1175), .A2(new_n906), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1168), .A2(new_n1172), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n756), .B1(new_n1179), .B2(KEYINPUT123), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(KEYINPUT123), .B2(new_n1179), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n779), .A2(new_n248), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n690), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1166), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1098), .B2(new_n689), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT124), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1091), .A2(new_n1092), .A3(new_n1043), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1187), .A2(new_n1084), .B1(new_n1096), .B2(new_n864), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n1093), .A3(new_n1100), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1102), .A2(new_n1189), .A3(new_n971), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT125), .ZN(G381));
  OR4_X1    g0992(.A1(G396), .A2(G390), .A3(G393), .A4(G384), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1193), .A2(G381), .A3(G387), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1051), .A2(new_n1076), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1083), .B2(new_n688), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n640), .B1(new_n1050), .B2(new_n1103), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1083), .A2(new_n1104), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G375), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1194), .A2(new_n1199), .A3(new_n1200), .ZN(G407));
  INV_X1    g1001(.A(G213), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(G343), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1199), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT126), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G213), .B(G407), .C1(new_n1206), .C2(new_n1207), .ZN(G409));
  NAND2_X1  g1008(.A1(new_n1203), .A2(G2897), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(KEYINPUT60), .B2(new_n1102), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1188), .A2(KEYINPUT60), .A3(new_n1093), .A4(new_n1100), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n639), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1098), .A2(new_n689), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1184), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT124), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT124), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1217), .B(new_n1184), .C1(new_n1098), .C2(new_n689), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1211), .A2(new_n1213), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(G384), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1100), .B1(new_n1188), .B2(new_n1093), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT60), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1189), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n639), .A3(new_n1212), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G384), .B1(new_n1186), .B2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1209), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1186), .A2(new_n1225), .A3(G384), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(G2897), .A4(new_n1203), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1227), .A2(KEYINPUT127), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT127), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1164), .C1(new_n1129), .C2(new_n1133), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1131), .A2(new_n1132), .A3(new_n971), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1199), .B1(new_n1235), .B2(new_n1163), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1203), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1233), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT63), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1221), .A2(new_n1226), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1241), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1203), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(KEYINPUT63), .A3(new_n1242), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(G393), .B(G396), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n969), .A2(new_n971), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n945), .B1(new_n1248), .B2(new_n689), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G390), .B1(new_n1249), .B2(new_n923), .ZN(new_n1250));
  INV_X1    g1050(.A(G390), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G387), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1247), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  XOR2_X1   g1054(.A(G393), .B(G396), .Z(new_n1255));
  NAND3_X1  g1055(.A1(new_n1249), .A2(new_n923), .A3(G390), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(new_n1251), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1253), .A2(new_n1254), .A3(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1240), .A2(new_n1244), .A3(new_n1246), .A4(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1245), .A2(new_n1261), .A3(new_n1242), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1254), .B1(new_n1245), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1261), .B1(new_n1245), .B2(new_n1242), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1262), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1253), .A2(new_n1258), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1260), .B1(new_n1266), .B2(new_n1268), .ZN(G405));
  NAND2_X1  g1069(.A1(G375), .A2(new_n1199), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n1234), .A3(new_n1243), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1243), .B1(new_n1270), .B2(new_n1234), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1267), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1273), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(G402));
endmodule


