//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n204), .B2(KEYINPUT84), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n208), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n220));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n220), .A2(new_n221), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n223), .B1(new_n222), .B2(new_n224), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n211), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n228), .B(KEYINPUT85), .Z(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n210), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n222), .A2(new_n224), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n227), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  INV_X1    g036(.A(G197gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT11), .B(G169gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT12), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n227), .A2(KEYINPUT18), .A3(new_n230), .A4(new_n233), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n222), .A2(new_n224), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n211), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n233), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT86), .B(KEYINPUT13), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n229), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n236), .A2(new_n242), .A3(new_n243), .A4(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT87), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n234), .A2(new_n235), .B1(new_n246), .B2(new_n249), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(KEYINPUT87), .A3(new_n242), .A4(new_n243), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n243), .ZN(new_n256));
  INV_X1    g055(.A(new_n242), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n253), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259));
  INV_X1    g058(.A(G211gat), .ZN(new_n260));
  INV_X1    g059(.A(G218gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n259), .B1(KEYINPUT22), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(G169gat), .ZN(new_n267));
  INV_X1    g066(.A(G176gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT26), .ZN(new_n270));
  NAND2_X1  g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT26), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n277));
  OR2_X1    g076(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G183gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT27), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G183gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n277), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n279), .ZN(new_n287));
  NOR2_X1   g086(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT28), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n276), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT64), .B1(new_n274), .B2(KEYINPUT23), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n294), .B(new_n295), .C1(G169gat), .C2(G176gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(KEYINPUT23), .B2(new_n274), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n278), .A2(new_n281), .A3(new_n279), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n273), .A2(KEYINPUT24), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n278), .A2(KEYINPUT66), .A3(new_n281), .A4(new_n279), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n300), .A2(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(new_n297), .A3(new_n299), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n292), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n266), .B1(new_n316), .B2(KEYINPUT29), .ZN(new_n317));
  INV_X1    g116(.A(new_n292), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n294), .B1(new_n269), .B2(new_n295), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n274), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n320));
  OAI211_X1 g119(.A(KEYINPUT25), .B(new_n299), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n301), .A2(new_n302), .B1(new_n304), .B2(new_n306), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n321), .B1(new_n308), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n271), .B1(new_n269), .B2(new_n295), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n324), .B1(new_n293), .B2(new_n296), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT25), .B1(new_n325), .B2(new_n312), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n318), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n266), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT70), .B1(new_n317), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n331), .B1(new_n333), .B2(new_n266), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n265), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G8gat), .B(G36gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT71), .ZN(new_n337));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n328), .B1(new_n327), .B2(new_n332), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n316), .A2(new_n266), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n341), .A2(new_n342), .A3(new_n265), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n335), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT72), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT72), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n335), .A2(new_n347), .A3(new_n340), .A4(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(G1gat), .B(G29gat), .Z(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G57gat), .B(G85gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G134gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G127gat), .ZN(new_n358));
  INV_X1    g157(.A(G127gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G134gat), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G120gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G113gat), .ZN(new_n363));
  INV_X1    g162(.A(G113gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G120gat), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT1), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT67), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n359), .B2(G134gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n361), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n358), .A2(new_n360), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n360), .A2(KEYINPUT67), .ZN(new_n371));
  XNOR2_X1  g170(.A(G113gat), .B(G120gat), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(KEYINPUT1), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n376));
  INV_X1    g175(.A(G155gat), .ZN(new_n377));
  INV_X1    g176(.A(G162gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G141gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G148gat), .ZN(new_n383));
  INV_X1    g182(.A(G148gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G141gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n385), .A3(KEYINPUT73), .ZN(new_n386));
  OR3_X1    g185(.A1(new_n384), .A2(KEYINPUT73), .A3(G141gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n377), .A2(new_n378), .ZN(new_n389));
  XNOR2_X1  g188(.A(G141gat), .B(G148gat), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n380), .B(new_n389), .C1(new_n390), .C2(KEYINPUT2), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n369), .A2(new_n373), .A3(new_n388), .A4(new_n391), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n356), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n388), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n388), .A2(new_n391), .A3(KEYINPUT74), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n388), .A2(new_n391), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n403), .A2(KEYINPUT3), .B1(new_n369), .B2(new_n373), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n369), .A2(new_n373), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n403), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n355), .B1(new_n408), .B2(new_n394), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n409), .A2(KEYINPUT75), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT75), .ZN(new_n412));
  AND4_X1   g211(.A1(new_n369), .A2(new_n373), .A3(new_n388), .A4(new_n391), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n369), .A2(new_n373), .B1(new_n388), .B2(new_n391), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n356), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n415), .B2(KEYINPUT5), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n406), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT77), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n394), .B2(KEYINPUT4), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n395), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n394), .A2(new_n418), .A3(KEYINPUT4), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n422), .A2(new_n410), .A3(new_n355), .A4(new_n405), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n354), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT6), .ZN(new_n426));
  INV_X1    g225(.A(new_n354), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT75), .B1(new_n409), .B2(new_n410), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n415), .A2(new_n412), .A3(KEYINPUT5), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n428), .A2(new_n429), .B1(new_n405), .B2(new_n396), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n355), .A2(new_n410), .ZN(new_n431));
  AOI221_X4 g230(.A(new_n431), .B1(new_n402), .B2(new_n404), .C1(new_n420), .C2(new_n421), .ZN(new_n432));
  OAI211_X1 g231(.A(KEYINPUT6), .B(new_n427), .C1(new_n430), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT83), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n427), .B1(new_n430), .B2(new_n432), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n354), .A3(new_n423), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n426), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n349), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n265), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n331), .B1(new_n341), .B2(new_n342), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n317), .A2(KEYINPUT70), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT37), .B1(new_n444), .B2(new_n343), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n335), .A2(new_n446), .A3(new_n344), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n445), .A2(KEYINPUT38), .A3(new_n339), .A4(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n441), .B1(new_n330), .B2(new_n334), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n341), .A2(new_n342), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n446), .B1(new_n450), .B2(new_n265), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n447), .A2(new_n339), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n448), .B1(new_n453), .B2(KEYINPUT38), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n440), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n346), .A2(new_n456), .A3(new_n348), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n340), .B1(new_n335), .B2(new_n344), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n444), .A2(new_n339), .A3(new_n343), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(KEYINPUT30), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n422), .A2(new_n405), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n356), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n413), .A2(new_n414), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n465), .B2(new_n355), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n420), .A2(new_n421), .B1(new_n402), .B2(new_n404), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(new_n355), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n468), .A3(new_n354), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n435), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n473));
  OR3_X1    g272(.A1(new_n469), .A2(new_n473), .A3(new_n470), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n473), .B1(new_n469), .B2(new_n470), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G228gat), .A2(G233gat), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT29), .B1(new_n400), .B2(new_n401), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n479), .A2(new_n441), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G22gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n397), .B1(new_n265), .B2(KEYINPUT29), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n403), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n480), .A2(new_n484), .A3(new_n486), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n489), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n482), .B1(new_n491), .B2(new_n487), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G78gat), .B(G106gat), .ZN(new_n494));
  INV_X1    g293(.A(G50gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT81), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT81), .A4(new_n498), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n455), .A2(new_n477), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n438), .A2(KEYINPUT78), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT78), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n435), .A2(new_n437), .A3(new_n506), .A4(new_n436), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n507), .A3(new_n433), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n457), .A3(new_n460), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n501), .A2(new_n502), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n300), .A2(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n407), .B1(new_n512), .B2(new_n292), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT34), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n374), .B(new_n318), .C1(new_n323), .C2(new_n326), .ZN(new_n515));
  NAND2_X1  g314(.A1(G227gat), .A2(G233gat), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT69), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n513), .A2(new_n516), .A3(new_n515), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT34), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n518), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G43gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(G71gat), .B(G99gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n516), .B1(new_n513), .B2(new_n515), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT32), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n516), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n310), .A2(new_n315), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n374), .B1(new_n532), .B2(new_n318), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n512), .A2(new_n407), .A3(new_n292), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT33), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(KEYINPUT68), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n528), .B2(KEYINPUT33), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n530), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(KEYINPUT32), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n526), .A2(new_n536), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n523), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n526), .B1(new_n535), .B2(KEYINPUT32), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT68), .B1(new_n535), .B2(new_n536), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n528), .A2(new_n538), .A3(KEYINPUT33), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n522), .A2(new_n521), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n517), .A2(new_n518), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n541), .A2(new_n542), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n544), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n554), .B1(new_n544), .B2(new_n553), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n504), .A2(new_n511), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n501), .A2(new_n502), .A3(new_n544), .A4(new_n553), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT35), .B1(new_n509), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n457), .A2(new_n460), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT35), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n439), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n540), .A2(new_n523), .A3(new_n543), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n551), .B1(new_n548), .B2(new_n552), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n561), .A2(new_n563), .A3(new_n503), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n258), .B1(new_n558), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571));
  INV_X1    g370(.A(G71gat), .ZN(new_n572));
  INV_X1    g371(.A(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT88), .ZN(new_n575));
  XOR2_X1   g374(.A(G57gat), .B(G64gat), .Z(new_n576));
  INV_X1    g375(.A(KEYINPUT88), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G71gat), .B(G78gat), .Z(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT8), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(KEYINPUT92), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(KEYINPUT92), .B2(new_n585), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT93), .B(G92gat), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n591));
  INV_X1    g390(.A(G92gat), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n591), .B(KEYINPUT7), .C1(new_n589), .C2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  OAI211_X1 g393(.A(G85gat), .B(G92gat), .C1(new_n594), .C2(KEYINPUT91), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n587), .A2(new_n590), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G99gat), .B(G106gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n587), .A2(new_n590), .A3(new_n596), .A4(new_n598), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n581), .A2(new_n600), .A3(new_n582), .A4(new_n601), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n605), .A2(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G230gat), .ZN(new_n609));
  INV_X1    g408(.A(G233gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n603), .A2(new_n605), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n611), .ZN(new_n615));
  XOR2_X1   g414(.A(G120gat), .B(G148gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT96), .ZN(new_n617));
  XOR2_X1   g416(.A(G176gat), .B(G204gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n613), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT98), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n620), .B1(new_n613), .B2(new_n615), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n625), .B1(new_n624), .B2(new_n627), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n583), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G127gat), .B(G155gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n211), .B1(new_n632), .B2(new_n583), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT89), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G183gat), .B(G211gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n637), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G232gat), .A2(G233gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT90), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n244), .B2(new_n602), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT94), .Z(new_n651));
  XNOR2_X1  g450(.A(G190gat), .B(G218gat), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT95), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n225), .A2(new_n226), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n656), .A2(new_n602), .B1(KEYINPUT95), .B2(new_n652), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n651), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n650), .B(KEYINPUT94), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n656), .A2(new_n602), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n654), .B(new_n653), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n662));
  XOR2_X1   g461(.A(G134gat), .B(G162gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n658), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n658), .B2(new_n661), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n645), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n570), .B1(new_n631), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n668), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n629), .A2(new_n630), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(KEYINPUT99), .A3(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n569), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n508), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g477(.A1(new_n674), .A2(new_n561), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n202), .B2(new_n679), .ZN(new_n682));
  MUX2_X1   g481(.A(new_n681), .B(new_n682), .S(KEYINPUT42), .Z(G1325gat));
  AOI21_X1  g482(.A(G15gat), .B1(new_n675), .B2(new_n566), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT100), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n555), .B2(new_n556), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT36), .B1(new_n564), .B2(new_n565), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n544), .A2(new_n553), .A3(new_n554), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(KEYINPUT101), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n687), .A2(new_n690), .A3(KEYINPUT102), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(G15gat), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n685), .B1(new_n675), .B2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n674), .A2(new_n503), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT43), .B(G22gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NOR2_X1   g500(.A1(new_n666), .A2(new_n667), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n558), .B2(new_n568), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n687), .A2(new_n690), .B1(new_n510), .B2(new_n509), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n706), .A2(new_n504), .B1(new_n560), .B2(new_n567), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n702), .A2(new_n705), .ZN(new_n708));
  OAI22_X1  g507(.A1(new_n704), .A2(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n644), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n253), .A2(new_n255), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n256), .A2(new_n257), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(new_n671), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT105), .Z(new_n717));
  NOR2_X1   g516(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT106), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT106), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n721), .B2(new_n508), .ZN(new_n722));
  AND4_X1   g521(.A1(new_n569), .A2(new_n644), .A3(new_n702), .A4(new_n671), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n216), .A3(new_n676), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(G1328gat));
  OAI21_X1  g526(.A(G36gat), .B1(new_n721), .B2(new_n561), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n723), .A2(new_n212), .A3(new_n461), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(KEYINPUT107), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n730), .A2(KEYINPUT107), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n728), .B(new_n733), .C1(new_n731), .C2(new_n729), .ZN(G1329gat));
  INV_X1    g533(.A(G43gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n723), .A2(new_n735), .A3(new_n566), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n710), .A2(new_n691), .A3(new_n717), .ZN(new_n737));
  NAND2_X1  g536(.A1(KEYINPUT47), .A2(G43gat), .ZN(new_n738));
  OAI221_X1 g537(.A(new_n736), .B1(KEYINPUT108), .B2(KEYINPUT47), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n736), .A2(KEYINPUT108), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n719), .A2(new_n696), .A3(new_n720), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(G43gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n742), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g542(.A1(new_n503), .A2(G50gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n723), .A2(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n710), .A2(new_n503), .A3(new_n717), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT48), .B(new_n745), .C1(new_n746), .C2(new_n495), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n719), .A2(new_n510), .A3(new_n720), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n748), .A2(G50gat), .B1(new_n723), .B2(new_n744), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g549(.A1(new_n504), .A2(new_n691), .A3(new_n511), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n568), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n671), .A2(new_n668), .A3(new_n715), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n508), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n561), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n754), .B2(new_n695), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n566), .A2(new_n572), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n754), .B2(new_n763), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g564(.A1(new_n754), .A2(new_n503), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(new_n573), .ZN(G1335gat));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n258), .A2(new_n768), .A3(new_n644), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n768), .B1(new_n258), .B2(new_n644), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n671), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n709), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774), .B2(new_n508), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n702), .B1(new_n769), .B2(new_n771), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT51), .B1(new_n752), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  AOI211_X1 g578(.A(new_n779), .B(new_n776), .C1(new_n751), .C2(new_n568), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n631), .A2(new_n589), .A3(new_n676), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n775), .B1(new_n781), .B2(new_n782), .ZN(G1336gat));
  INV_X1    g582(.A(new_n774), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n588), .B1(new_n784), .B2(new_n461), .ZN(new_n785));
  INV_X1    g584(.A(new_n781), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n671), .A2(G92gat), .A3(new_n561), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1337gat));
  INV_X1    g589(.A(G99gat), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n786), .A2(new_n791), .A3(new_n566), .A4(new_n631), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n784), .A2(new_n696), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT111), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G99gat), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(KEYINPUT111), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n792), .B1(new_n795), .B2(new_n796), .ZN(G1338gat));
  AND3_X1   g596(.A1(new_n455), .A2(new_n477), .A3(new_n503), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n511), .A2(new_n557), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n568), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n705), .B1(new_n800), .B2(new_n702), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n707), .A2(new_n708), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n510), .B(new_n773), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  XOR2_X1   g602(.A(KEYINPUT112), .B(G106gat), .Z(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n671), .A2(G106gat), .A3(new_n503), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n778), .B2(new_n780), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT53), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n804), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n709), .A2(KEYINPUT113), .A3(new_n510), .A4(new_n773), .ZN(new_n816));
  AOI211_X1 g615(.A(new_n811), .B(new_n813), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n803), .A2(new_n814), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n805), .A3(new_n816), .ZN(new_n819));
  INV_X1    g618(.A(new_n813), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT114), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n810), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g623(.A(KEYINPUT115), .B(new_n810), .C1(new_n817), .C2(new_n821), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1339gat));
  NAND3_X1  g625(.A1(new_n670), .A2(new_n258), .A3(new_n671), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT116), .B1(new_n608), .B2(new_n612), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n606), .A2(new_n607), .A3(new_n831), .A4(new_n611), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n830), .A2(new_n613), .A3(KEYINPUT54), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n611), .B1(new_n606), .B2(new_n607), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n620), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n621), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n833), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n829), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n839), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n841), .A2(KEYINPUT117), .A3(new_n621), .A4(new_n837), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n842), .A3(new_n715), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n227), .A2(new_n233), .ZN(new_n844));
  OAI22_X1  g643(.A1(new_n844), .A2(new_n230), .B1(new_n246), .B2(new_n249), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n253), .A2(new_n255), .B1(new_n845), .B2(new_n241), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n629), .B2(new_n630), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n702), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  AND4_X1   g647(.A1(new_n702), .A2(new_n846), .A3(new_n840), .A4(new_n842), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n828), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n712), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n848), .A2(new_n849), .A3(new_n828), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n827), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n853), .A2(new_n503), .A3(new_n566), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n461), .A2(new_n508), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n258), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(new_n364), .ZN(G1340gat));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n671), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(new_n362), .ZN(G1341gat));
  OAI21_X1  g659(.A(G127gat), .B1(new_n856), .B2(new_n712), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n645), .A2(new_n359), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n856), .B2(new_n862), .ZN(G1342gat));
  NAND2_X1  g662(.A1(new_n702), .A2(new_n561), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(G134gat), .A3(new_n508), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT56), .Z(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n856), .B2(new_n703), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1343gat));
  NAND2_X1  g668(.A1(new_n691), .A2(new_n855), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n258), .A2(new_n382), .ZN(new_n872));
  XOR2_X1   g671(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(new_n853), .B2(new_n510), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n838), .A2(new_n839), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n715), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n702), .B1(new_n847), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n644), .B1(new_n879), .B2(new_n849), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n876), .B(new_n503), .C1(new_n880), .C2(new_n827), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n871), .B(new_n872), .C1(new_n875), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n696), .A2(new_n508), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n853), .A2(new_n510), .A3(new_n561), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n382), .B1(new_n884), .B2(new_n258), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(KEYINPUT58), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT58), .B1(new_n882), .B2(new_n885), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT121), .B(KEYINPUT58), .C1(new_n882), .C2(new_n885), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n888), .A2(new_n889), .B1(new_n892), .B2(new_n893), .ZN(G1344gat));
  INV_X1    g693(.A(new_n884), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n384), .A3(new_n631), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n871), .B1(new_n875), .B2(new_n881), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n671), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(KEYINPUT59), .A3(new_n384), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n853), .A2(new_n510), .A3(new_n874), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n669), .A2(new_n672), .A3(new_n258), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n702), .A2(new_n846), .A3(new_n877), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n644), .B1(new_n879), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n503), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n906), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT122), .B1(new_n906), .B2(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n631), .B(new_n871), .C1(new_n902), .C2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n900), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n896), .B1(new_n899), .B2(new_n911), .ZN(G1345gat));
  OAI21_X1  g711(.A(G155gat), .B1(new_n897), .B2(new_n712), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n377), .A3(new_n645), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n897), .B2(new_n703), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n853), .A2(new_n510), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n864), .A2(G162gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n883), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n561), .A2(new_n676), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n854), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n715), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n921), .B(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n566), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n510), .B1(new_n925), .B2(KEYINPUT124), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n853), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n258), .A2(new_n267), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(G1348gat));
  NAND3_X1  g729(.A1(new_n928), .A2(G176gat), .A3(new_n631), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT125), .ZN(new_n932));
  AOI21_X1  g731(.A(G176gat), .B1(new_n922), .B2(new_n631), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n922), .A2(new_n290), .A3(new_n645), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n853), .A2(new_n926), .A3(new_n927), .ZN(new_n936));
  OAI21_X1  g735(.A(G183gat), .B1(new_n936), .B2(new_n712), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT60), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n935), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n922), .A2(new_n289), .A3(new_n702), .ZN(new_n943));
  OAI21_X1  g742(.A(G190gat), .B1(new_n936), .B2(new_n703), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1351gat));
  OR3_X1    g746(.A1(new_n902), .A2(new_n909), .A3(KEYINPUT126), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n924), .A2(new_n695), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT126), .B1(new_n902), .B2(new_n909), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n258), .A2(new_n238), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n695), .A2(new_n921), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n917), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n238), .B1(new_n954), .B2(new_n258), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n952), .A2(new_n955), .ZN(G1352gat));
  NAND4_X1  g755(.A1(new_n948), .A2(new_n631), .A3(new_n949), .A4(new_n950), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G204gat), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n954), .A2(G204gat), .A3(new_n671), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1353gat));
  NAND4_X1  g760(.A1(new_n917), .A2(new_n260), .A3(new_n645), .A4(new_n953), .ZN(new_n962));
  NOR2_X1   g761(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n949), .A2(new_n645), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n907), .A2(new_n908), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n901), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n966), .B2(new_n260), .ZN(new_n967));
  NAND2_X1  g766(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n966), .A2(new_n260), .A3(new_n963), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n962), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  NOR2_X1   g770(.A1(new_n703), .A2(new_n261), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n261), .B1(new_n954), .B2(new_n703), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(G1355gat));
endmodule


