//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n445, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1116, new_n1117, new_n1118,
    new_n1119;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g031(.A1(new_n439), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(G567), .A2(new_n459), .B1(new_n456), .B2(G2106), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n470), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n472), .B1(G2105), .B2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n470), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n470), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n480), .B1(new_n483), .B2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n481), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT69), .Z(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT70), .Z(G162));
  NAND4_X1  g064(.A1(new_n468), .A2(G138), .A3(new_n481), .A4(new_n469), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR4_X1   g070(.A1(new_n475), .A2(KEYINPUT4), .A3(new_n495), .A4(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n468), .A2(new_n469), .ZN(new_n500));
  INV_X1    g075(.A(G126), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n463), .A2(G2105), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n502), .A2(G2105), .B1(G102), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT72), .B(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(new_n508), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G75), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n507), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(G62), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(G166));
  NAND2_X1  g097(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n509), .A2(new_n511), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n523), .A2(G543), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n512), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n528), .B(new_n530), .C1(new_n518), .C2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(new_n527), .A2(G52), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n524), .A2(new_n518), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n518), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n537), .A2(G90), .B1(new_n514), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n536), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n527), .A2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n537), .A2(G81), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT75), .Z(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(new_n514), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT76), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(new_n554));
  XOR2_X1   g129(.A(new_n554), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(new_n527), .A2(G53), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n537), .A2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT78), .B(G65), .Z(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n518), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n560), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n566), .B(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n527), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n537), .A2(G87), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(new_n514), .A2(G73), .ZN(new_n575));
  INV_X1    g150(.A(G48), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n524), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n514), .A2(G61), .ZN(new_n579));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n524), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(new_n517), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  XNOR2_X1  g159(.A(KEYINPUT81), .B(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n527), .A2(G47), .B1(new_n537), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT82), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n508), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n537), .A2(G92), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT10), .Z(new_n594));
  NAND2_X1  g169(.A1(new_n527), .A2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT83), .B(G66), .Z(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n518), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n566), .B(KEYINPUT79), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  XNOR2_X1  g181(.A(G297), .B(KEYINPUT84), .ZN(G280));
  NOR2_X1   g182(.A1(new_n600), .A2(G559), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G860), .B2(new_n601), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT85), .ZN(G148));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n549), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n608), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g189(.A(G135), .ZN(new_n615));
  OR3_X1    g190(.A1(new_n482), .A2(KEYINPUT87), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n480), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n481), .A2(G111), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT88), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n620));
  OAI21_X1  g195(.A(KEYINPUT87), .B1(new_n482), .B2(new_n615), .ZN(new_n621));
  NAND4_X1  g196(.A1(new_n616), .A2(new_n617), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n481), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT86), .B(G2100), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n624), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2435), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2438), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G14), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2067), .B(G2678), .Z(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  AOI21_X1  g227(.A(new_n648), .B1(KEYINPUT17), .B2(new_n650), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n646), .A2(new_n647), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n653), .B(new_n654), .C1(KEYINPUT17), .C2(new_n650), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n649), .B(KEYINPUT89), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n652), .B(new_n655), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(new_n623), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(G227));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n671), .C1(new_n669), .C2(new_n668), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(G1986), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT90), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT22), .B(G1981), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(G229));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n680), .A2(KEYINPUT23), .A3(G20), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT23), .ZN(new_n682));
  INV_X1    g257(.A(G20), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G16), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n681), .B(new_n684), .C1(new_n605), .C2(new_n680), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1956), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT31), .B(G11), .ZN(new_n687));
  INV_X1    g262(.A(G2084), .ZN(new_n688));
  INV_X1    g263(.A(G160), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT91), .B(G29), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT24), .B(G34), .Z(new_n692));
  OAI22_X1  g267(.A1(new_n689), .A2(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(G16), .A2(G19), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n550), .B2(G16), .ZN(new_n695));
  OAI221_X1 g270(.A(new_n687), .B1(new_n688), .B2(new_n693), .C1(new_n695), .C2(G1341), .ZN(new_n696));
  NOR2_X1   g271(.A1(G4), .A2(G16), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n601), .B2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G1961), .ZN(new_n699));
  OAI21_X1  g274(.A(KEYINPUT99), .B1(G5), .B2(G16), .ZN(new_n700));
  OR3_X1    g275(.A1(KEYINPUT99), .A2(G5), .A3(G16), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n700), .B(new_n701), .C1(G301), .C2(new_n680), .ZN(new_n702));
  OAI22_X1  g277(.A1(new_n698), .A2(G1348), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G29), .A2(G32), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n503), .A2(G105), .ZN(new_n705));
  INV_X1    g280(.A(G129), .ZN(new_n706));
  INV_X1    g281(.A(G141), .ZN(new_n707));
  OAI221_X1 g282(.A(new_n705), .B1(new_n479), .B2(new_n706), .C1(new_n707), .C2(new_n482), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT97), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT26), .Z(new_n711));
  NOR2_X1   g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n704), .B1(new_n712), .B2(G29), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G1996), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n480), .A2(G128), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n483), .A2(G140), .ZN(new_n717));
  NOR2_X1   g292(.A1(G104), .A2(G2105), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(new_n481), .B2(G116), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n691), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n721), .A2(G26), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n720), .A2(G29), .B1(KEYINPUT28), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(KEYINPUT28), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2067), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n715), .B(new_n725), .C1(new_n688), .C2(new_n693), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n698), .A2(G1348), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n690), .A2(G33), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n483), .A2(G139), .ZN(new_n729));
  NAND2_X1  g304(.A1(G115), .A2(G2104), .ZN(new_n730));
  INV_X1    g305(.A(G127), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n475), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G2105), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n503), .A2(G103), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  NAND3_X1  g310(.A1(new_n729), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n728), .B1(new_n737), .B2(new_n690), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G2072), .Z(new_n739));
  OR2_X1    g314(.A1(new_n622), .A2(new_n721), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT30), .B(G28), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n702), .A2(new_n699), .B1(new_n690), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n721), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n721), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n695), .A2(G1341), .B1(G2078), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n726), .A2(new_n727), .A3(new_n743), .A4(new_n746), .ZN(new_n747));
  NOR4_X1   g322(.A1(new_n686), .A2(new_n696), .A3(new_n703), .A4(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G16), .A2(G23), .ZN(new_n749));
  INV_X1    g324(.A(G288), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT33), .B(G1976), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n680), .A2(G22), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G166), .B2(new_n680), .ZN(new_n755));
  INV_X1    g330(.A(G1971), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n680), .A2(G6), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n583), .B2(new_n680), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT32), .B(G1981), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n753), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT34), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n680), .A2(G24), .ZN(new_n764));
  INV_X1    g339(.A(G290), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n680), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT95), .B(G1986), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n480), .A2(G119), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n483), .A2(G131), .ZN(new_n770));
  NOR2_X1   g345(.A1(G95), .A2(G2105), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(new_n481), .B2(G107), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n769), .B(new_n770), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT93), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(new_n691), .ZN(new_n775));
  INV_X1    g350(.A(G25), .ZN(new_n776));
  OAI21_X1  g351(.A(KEYINPUT92), .B1(new_n691), .B2(new_n776), .ZN(new_n777));
  OR3_X1    g352(.A1(new_n691), .A2(KEYINPUT92), .A3(new_n776), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT35), .B(G1991), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT94), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n779), .B(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n763), .A2(new_n768), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(KEYINPUT36), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(KEYINPUT36), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n748), .B(new_n787), .C1(new_n785), .C2(new_n783), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n745), .A2(G2078), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n691), .A2(G35), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G162), .B2(new_n691), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT29), .B(G2090), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G21), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G168), .B2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT98), .B(G1966), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n788), .A2(new_n789), .A3(new_n793), .A4(new_n797), .ZN(G311));
  INV_X1    g373(.A(G311), .ZN(G150));
  NAND2_X1  g374(.A1(new_n527), .A2(G55), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n537), .A2(G93), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n800), .B(new_n801), .C1(new_n508), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G860), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT37), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n601), .A2(G559), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT38), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT39), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n803), .B1(new_n550), .B2(KEYINPUT100), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n550), .A2(KEYINPUT100), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n809), .B(new_n810), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n808), .B(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n805), .B1(new_n812), .B2(G860), .ZN(G145));
  XNOR2_X1  g388(.A(new_n712), .B(new_n720), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT101), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n505), .B(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT102), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(KEYINPUT102), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n818), .A2(new_n737), .A3(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT103), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(KEYINPUT103), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n817), .B(KEYINPUT104), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n821), .A2(new_n822), .B1(new_n736), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(G142), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n481), .A2(G118), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT105), .Z(new_n828));
  OAI22_X1  g403(.A1(new_n482), .A2(new_n825), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G130), .B2(new_n480), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n626), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n774), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT106), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n824), .B(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n622), .B(G160), .Z(new_n835));
  XNOR2_X1  g410(.A(G162), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(G37), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n824), .A2(new_n833), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n839), .B(new_n836), .C1(new_n832), .C2(new_n824), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g417(.A1(new_n803), .A2(new_n611), .ZN(new_n843));
  XNOR2_X1  g418(.A(G290), .B(new_n750), .ZN(new_n844));
  XNOR2_X1  g419(.A(G166), .B(new_n583), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT108), .Z(new_n848));
  AND2_X1   g423(.A1(new_n844), .A2(new_n846), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(KEYINPUT109), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(KEYINPUT109), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT42), .Z(new_n853));
  AOI21_X1  g428(.A(new_n601), .B1(G299), .B2(KEYINPUT107), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT107), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n605), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n854), .B(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n811), .B(new_n608), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(KEYINPUT41), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n860), .B2(new_n858), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n853), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n843), .B1(new_n862), .B2(new_n611), .ZN(G295));
  OAI21_X1  g438(.A(new_n843), .B1(new_n862), .B2(new_n611), .ZN(G331));
  XNOR2_X1  g439(.A(G168), .B(G301), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n811), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n857), .A2(new_n867), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n852), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n868), .A2(new_n852), .A3(new_n870), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT43), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n868), .A2(KEYINPUT110), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(new_n878), .A3(new_n872), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n868), .B(new_n870), .C1(KEYINPUT110), .C2(new_n852), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n874), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(new_n880), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n879), .A2(KEYINPUT43), .A3(new_n874), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  MUX2_X1   g461(.A(new_n883), .B(new_n886), .S(KEYINPUT44), .Z(G397));
  INV_X1    g462(.A(G1384), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT45), .B1(new_n816), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(G160), .A2(G40), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G1996), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT111), .Z(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT46), .Z(new_n896));
  INV_X1    g471(.A(new_n892), .ZN(new_n897));
  INV_X1    g472(.A(G2067), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n720), .B(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n899), .A2(new_n712), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n896), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT47), .Z(new_n902));
  AOI21_X1  g477(.A(KEYINPUT112), .B1(new_n895), .B2(new_n712), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n895), .A2(KEYINPUT112), .A3(new_n712), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n899), .B1(new_n893), .B2(new_n712), .ZN(new_n905));
  AOI211_X1 g480(.A(new_n903), .B(new_n904), .C1(new_n892), .C2(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n774), .B(new_n780), .Z(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(new_n897), .B2(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(G290), .A2(G1986), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n897), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT48), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n774), .A2(new_n780), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n720), .A2(G2067), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n897), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n902), .A2(new_n912), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT127), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT53), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n816), .A2(KEYINPUT45), .A3(new_n888), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n920), .A2(new_n891), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n493), .B1(new_n490), .B2(KEYINPUT4), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n922), .A2(new_n923), .A3(new_n496), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n502), .A2(G2105), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n503), .A2(G102), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n888), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n921), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n919), .B1(new_n931), .B2(G2078), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT126), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(KEYINPUT113), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT113), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n505), .A2(new_n936), .A3(new_n888), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n890), .B1(KEYINPUT50), .B2(new_n928), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n699), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n932), .A2(new_n933), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n938), .A2(KEYINPUT45), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n891), .B1(new_n929), .B2(new_n928), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n919), .A2(G2078), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n934), .A2(new_n944), .A3(new_n945), .A4(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1966), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n942), .A2(new_n688), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(G168), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(G8), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT51), .ZN(new_n958));
  AOI21_X1  g533(.A(G168), .B1(new_n954), .B2(new_n955), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n960));
  OAI211_X1 g535(.A(G8), .B(new_n956), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n958), .A2(new_n961), .A3(KEYINPUT62), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT62), .B1(new_n958), .B2(new_n961), .ZN(new_n963));
  OAI211_X1 g538(.A(G171), .B(new_n952), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n931), .A2(new_n756), .ZN(new_n966));
  INV_X1    g541(.A(G2090), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n942), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n965), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(G166), .A2(new_n965), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT55), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n935), .A2(KEYINPUT50), .A3(new_n937), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n974), .A2(KEYINPUT117), .A3(new_n891), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT117), .B1(new_n974), .B2(new_n891), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n928), .A2(KEYINPUT50), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n967), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n965), .B1(new_n979), .B2(new_n966), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(new_n971), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n982));
  NAND2_X1  g557(.A1(G305), .A2(G1981), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n583), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(KEYINPUT114), .A3(new_n985), .ZN(new_n986));
  OR3_X1    g561(.A1(new_n583), .A2(KEYINPUT114), .A3(new_n984), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n982), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n938), .A2(new_n891), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(new_n965), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n986), .A2(new_n982), .A3(new_n987), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n990), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n750), .A2(G1976), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT52), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(G288), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n993), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n981), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n973), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n997), .A2(new_n1001), .A3(new_n750), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n985), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n993), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n997), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1011), .B(new_n972), .C1(new_n971), .C2(new_n980), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n954), .A2(new_n955), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1013), .A2(new_n965), .A3(G286), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1010), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1005), .A2(KEYINPUT118), .A3(new_n972), .A4(new_n1014), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT63), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n971), .A2(KEYINPUT119), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n969), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1018), .B1(new_n969), .B2(new_n1021), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n1011), .A4(new_n1014), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1006), .A2(new_n1009), .A3(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT122), .B(G2072), .Z(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT56), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n921), .A2(new_n930), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n936), .B1(new_n505), .B2(new_n888), .ZN(new_n1031));
  AOI211_X1 g606(.A(KEYINPUT113), .B(G1384), .C1(new_n498), .C2(new_n504), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n939), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1030), .B1(new_n1033), .B2(new_n890), .ZN(new_n1034));
  INV_X1    g609(.A(new_n977), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n974), .A2(KEYINPUT117), .A3(new_n891), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n1038));
  INV_X1    g613(.A(G1956), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1029), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n560), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(new_n566), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1348), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n943), .A2(new_n1049), .B1(new_n898), .B2(new_n992), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n600), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT120), .B1(new_n978), .B2(G1956), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1047), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n1029), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1055), .B1(new_n1054), .B2(new_n1029), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1029), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1047), .B(new_n1060), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT61), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT61), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1048), .A2(new_n1056), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n920), .A2(new_n893), .A3(new_n930), .A4(new_n891), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT58), .B(G1341), .Z(new_n1068));
  NAND2_X1  g643(.A1(new_n991), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n549), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1066), .B1(new_n1071), .B2(KEYINPUT59), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1070), .A2(KEYINPUT123), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1071), .B2(KEYINPUT59), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1070), .A2(KEYINPUT124), .A3(new_n1073), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT125), .B1(new_n1065), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT125), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1083), .B(new_n1080), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1050), .A2(KEYINPUT60), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(new_n601), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(KEYINPUT60), .B2(new_n1050), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1058), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1012), .ZN(new_n1090));
  XNOR2_X1  g665(.A(G301), .B(KEYINPUT54), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n952), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n921), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(new_n889), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1094), .B2(new_n950), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n934), .A2(new_n944), .A3(new_n945), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n958), .A2(new_n961), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1090), .A2(new_n1092), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1026), .B1(new_n1089), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(G290), .A2(G1986), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n897), .B1(new_n909), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n908), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n918), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1048), .A2(new_n1056), .A3(new_n1063), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1063), .B1(new_n1048), .B2(new_n1056), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1081), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1083), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1065), .A2(KEYINPUT125), .A3(new_n1081), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n1088), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1098), .B1(new_n1109), .B2(new_n1057), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1006), .A2(new_n1025), .A3(new_n1009), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1102), .B(new_n918), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n917), .B1(new_n1103), .B2(new_n1113), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g689(.A(G319), .B1(new_n642), .B2(new_n643), .ZN(new_n1116));
  AOI21_X1  g690(.A(new_n1116), .B1(new_n877), .B2(new_n882), .ZN(new_n1117));
  INV_X1    g691(.A(G229), .ZN(new_n1118));
  NOR2_X1   g692(.A1(new_n841), .A2(G227), .ZN(new_n1119));
  AND3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(G308));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(G225));
endmodule


