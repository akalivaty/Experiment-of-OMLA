

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n736), .A2(n697), .ZN(n699) );
  OR2_X1 U553 ( .A1(n686), .A2(n685), .ZN(n758) );
  NOR2_X1 U554 ( .A1(G651), .A2(n638), .ZN(n645) );
  XOR2_X1 U555 ( .A(G543), .B(KEYINPUT0), .Z(n638) );
  INV_X1 U556 ( .A(G651), .ZN(n520) );
  NOR2_X1 U557 ( .A1(n638), .A2(n520), .ZN(n641) );
  NAND2_X1 U558 ( .A1(G77), .A2(n641), .ZN(n517) );
  NOR2_X1 U559 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U560 ( .A1(G90), .A2(n642), .ZN(n516) );
  NAND2_X1 U561 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U562 ( .A(KEYINPUT9), .B(n518), .ZN(n526) );
  NAND2_X1 U563 ( .A1(G52), .A2(n645), .ZN(n519) );
  XOR2_X1 U564 ( .A(KEYINPUT72), .B(n519), .Z(n524) );
  NOR2_X1 U565 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U566 ( .A(KEYINPUT1), .B(n521), .Z(n646) );
  NAND2_X1 U567 ( .A1(G64), .A2(n646), .ZN(n522) );
  XNOR2_X1 U568 ( .A(KEYINPUT71), .B(n522), .ZN(n523) );
  NOR2_X1 U569 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n526), .A2(n525), .ZN(G301) );
  INV_X1 U571 ( .A(G301), .ZN(G171) );
  XOR2_X1 U572 ( .A(KEYINPUT104), .B(G2435), .Z(n528) );
  XNOR2_X1 U573 ( .A(G2454), .B(G2438), .ZN(n527) );
  XNOR2_X1 U574 ( .A(n528), .B(n527), .ZN(n532) );
  XOR2_X1 U575 ( .A(G2427), .B(G2443), .Z(n530) );
  XNOR2_X1 U576 ( .A(KEYINPUT103), .B(G2446), .ZN(n529) );
  XNOR2_X1 U577 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U578 ( .A(n532), .B(n531), .Z(n534) );
  XNOR2_X1 U579 ( .A(KEYINPUT102), .B(G2451), .ZN(n533) );
  XNOR2_X1 U580 ( .A(n534), .B(n533), .ZN(n537) );
  XOR2_X1 U581 ( .A(G1348), .B(G1341), .Z(n535) );
  XNOR2_X1 U582 ( .A(G2430), .B(n535), .ZN(n536) );
  XOR2_X1 U583 ( .A(n537), .B(n536), .Z(n538) );
  AND2_X1 U584 ( .A1(G14), .A2(n538), .ZN(G401) );
  AND2_X1 U585 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U586 ( .A(G860), .B(KEYINPUT76), .Z(n591) );
  NAND2_X1 U587 ( .A1(G56), .A2(n646), .ZN(n539) );
  XOR2_X1 U588 ( .A(KEYINPUT14), .B(n539), .Z(n545) );
  NAND2_X1 U589 ( .A1(n642), .A2(G81), .ZN(n540) );
  XNOR2_X1 U590 ( .A(n540), .B(KEYINPUT12), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G68), .A2(n641), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U593 ( .A(KEYINPUT13), .B(n543), .Z(n544) );
  NOR2_X1 U594 ( .A1(n545), .A2(n544), .ZN(n547) );
  NAND2_X1 U595 ( .A1(n645), .A2(G43), .ZN(n546) );
  NAND2_X1 U596 ( .A1(n547), .A2(n546), .ZN(n938) );
  OR2_X1 U597 ( .A1(n591), .A2(n938), .ZN(G153) );
  INV_X1 U598 ( .A(G57), .ZN(G237) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  INV_X1 U601 ( .A(G2105), .ZN(n550) );
  NOR2_X1 U602 ( .A1(G2104), .A2(n550), .ZN(n883) );
  NAND2_X1 U603 ( .A1(G125), .A2(n883), .ZN(n549) );
  AND2_X1 U604 ( .A1(G2105), .A2(G2104), .ZN(n884) );
  NAND2_X1 U605 ( .A1(G113), .A2(n884), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n684) );
  AND2_X1 U607 ( .A1(n550), .A2(G2104), .ZN(n888) );
  NAND2_X1 U608 ( .A1(G101), .A2(n888), .ZN(n551) );
  XNOR2_X1 U609 ( .A(n551), .B(KEYINPUT65), .ZN(n552) );
  XNOR2_X1 U610 ( .A(KEYINPUT23), .B(n552), .ZN(n558) );
  XNOR2_X1 U611 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n554) );
  NOR2_X1 U612 ( .A1(G2105), .A2(G2104), .ZN(n553) );
  XNOR2_X1 U613 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X2 U614 ( .A(KEYINPUT66), .B(n555), .ZN(n891) );
  NAND2_X1 U615 ( .A1(n891), .A2(G137), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n556), .B(KEYINPUT68), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n686) );
  NOR2_X1 U618 ( .A1(n684), .A2(n686), .ZN(G160) );
  NAND2_X1 U619 ( .A1(G51), .A2(n645), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G63), .A2(n646), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U622 ( .A(KEYINPUT6), .B(n561), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n642), .A2(G89), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U625 ( .A1(G76), .A2(n641), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U627 ( .A(n565), .B(KEYINPUT5), .Z(n566) );
  NOR2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT77), .B(n568), .Z(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT7), .B(n569), .Z(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n831) );
  NAND2_X1 U635 ( .A1(n831), .A2(G567), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT75), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT11), .B(n572), .ZN(G234) );
  NAND2_X1 U638 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G92), .A2(n642), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G66), .A2(n646), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G79), .A2(n641), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G54), .A2(n645), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT15), .B(n579), .Z(n922) );
  OR2_X1 U647 ( .A1(n922), .A2(G868), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U649 ( .A1(G91), .A2(n642), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G65), .A2(n646), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G78), .A2(n641), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G53), .A2(n645), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT73), .B(n588), .Z(n928) );
  XOR2_X1 U657 ( .A(KEYINPUT74), .B(n928), .Z(G299) );
  NOR2_X1 U658 ( .A1(G299), .A2(G868), .ZN(n590) );
  INV_X1 U659 ( .A(G868), .ZN(n658) );
  NOR2_X1 U660 ( .A1(G286), .A2(n658), .ZN(n589) );
  NOR2_X1 U661 ( .A1(n590), .A2(n589), .ZN(G297) );
  NAND2_X1 U662 ( .A1(G559), .A2(n591), .ZN(n592) );
  XNOR2_X1 U663 ( .A(KEYINPUT78), .B(n592), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n593), .A2(n922), .ZN(n594) );
  XNOR2_X1 U665 ( .A(KEYINPUT16), .B(n594), .ZN(G148) );
  NOR2_X1 U666 ( .A1(G868), .A2(n938), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G868), .A2(n922), .ZN(n595) );
  NOR2_X1 U668 ( .A1(G559), .A2(n595), .ZN(n596) );
  NOR2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U670 ( .A(KEYINPUT79), .B(n598), .Z(G282) );
  NAND2_X1 U671 ( .A1(G123), .A2(n883), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n599), .B(KEYINPUT18), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n888), .A2(G99), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U675 ( .A1(n884), .A2(G111), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G135), .A2(n891), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n977) );
  XNOR2_X1 U679 ( .A(n977), .B(G2096), .ZN(n607) );
  INV_X1 U680 ( .A(G2100), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(G156) );
  NAND2_X1 U682 ( .A1(G93), .A2(n642), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G67), .A2(n646), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n641), .A2(G80), .ZN(n610) );
  XOR2_X1 U686 ( .A(KEYINPUT80), .B(n610), .Z(n611) );
  NOR2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n645), .A2(G55), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n659) );
  NAND2_X1 U690 ( .A1(G559), .A2(n922), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n938), .B(n615), .ZN(n656) );
  NOR2_X1 U692 ( .A1(G860), .A2(n656), .ZN(n616) );
  XOR2_X1 U693 ( .A(n659), .B(n616), .Z(G145) );
  NAND2_X1 U694 ( .A1(n641), .A2(G73), .ZN(n617) );
  XNOR2_X1 U695 ( .A(KEYINPUT2), .B(n617), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n642), .A2(G86), .ZN(n618) );
  XOR2_X1 U697 ( .A(KEYINPUT81), .B(n618), .Z(n620) );
  NAND2_X1 U698 ( .A1(n646), .A2(G61), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U700 ( .A(KEYINPUT82), .B(n621), .Z(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U702 ( .A(n624), .B(KEYINPUT83), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G48), .A2(n645), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U705 ( .A1(G60), .A2(n646), .ZN(n627) );
  XNOR2_X1 U706 ( .A(n627), .B(KEYINPUT70), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n641), .A2(G72), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G85), .A2(n642), .ZN(n630) );
  XNOR2_X1 U710 ( .A(KEYINPUT69), .B(n630), .ZN(n631) );
  NOR2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n645), .A2(G47), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(G290) );
  NAND2_X1 U714 ( .A1(G49), .A2(n645), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U717 ( .A1(n646), .A2(n637), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n638), .A2(G87), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G75), .A2(n641), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G88), .A2(n642), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G50), .A2(n645), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G62), .A2(n646), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(G166) );
  XNOR2_X1 U727 ( .A(G299), .B(G305), .ZN(n655) );
  XNOR2_X1 U728 ( .A(G290), .B(G288), .ZN(n653) );
  XNOR2_X1 U729 ( .A(G166), .B(KEYINPUT19), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(n659), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n655), .B(n654), .ZN(n836) );
  XNOR2_X1 U733 ( .A(n836), .B(n656), .ZN(n657) );
  NOR2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n661) );
  NOR2_X1 U735 ( .A1(G868), .A2(n659), .ZN(n660) );
  NOR2_X1 U736 ( .A1(n661), .A2(n660), .ZN(G295) );
  XOR2_X1 U737 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n663) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n666), .A2(G2072), .ZN(n667) );
  XOR2_X1 U743 ( .A(KEYINPUT85), .B(n667), .Z(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U745 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U748 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U749 ( .A1(G96), .A2(n670), .ZN(n916) );
  NAND2_X1 U750 ( .A1(n916), .A2(G2106), .ZN(n674) );
  NAND2_X1 U751 ( .A1(G108), .A2(G120), .ZN(n671) );
  NOR2_X1 U752 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G69), .A2(n672), .ZN(n917) );
  NAND2_X1 U754 ( .A1(n917), .A2(G567), .ZN(n673) );
  NAND2_X1 U755 ( .A1(n674), .A2(n673), .ZN(n918) );
  NOR2_X1 U756 ( .A1(n675), .A2(n918), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n676), .B(KEYINPUT86), .ZN(n833) );
  NAND2_X1 U758 ( .A1(G36), .A2(n833), .ZN(G176) );
  NAND2_X1 U759 ( .A1(n888), .A2(G102), .ZN(n678) );
  NAND2_X1 U760 ( .A1(G138), .A2(n891), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G126), .A2(n883), .ZN(n680) );
  NAND2_X1 U763 ( .A1(G114), .A2(n884), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U765 ( .A1(n682), .A2(n681), .ZN(G164) );
  INV_X1 U766 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U767 ( .A(KEYINPUT31), .B(KEYINPUT96), .ZN(n696) );
  INV_X1 U768 ( .A(G40), .ZN(n683) );
  OR2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n685) );
  INV_X1 U770 ( .A(n758), .ZN(n687) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n759) );
  NAND2_X1 U772 ( .A1(n687), .A2(n759), .ZN(n736) );
  NAND2_X1 U773 ( .A1(G8), .A2(n736), .ZN(n805) );
  NOR2_X1 U774 ( .A1(G1966), .A2(n805), .ZN(n750) );
  NOR2_X1 U775 ( .A1(G2084), .A2(n736), .ZN(n746) );
  NOR2_X1 U776 ( .A1(n750), .A2(n746), .ZN(n688) );
  NAND2_X1 U777 ( .A1(G8), .A2(n688), .ZN(n689) );
  XNOR2_X1 U778 ( .A(KEYINPUT30), .B(n689), .ZN(n690) );
  NOR2_X1 U779 ( .A1(G168), .A2(n690), .ZN(n694) );
  INV_X1 U780 ( .A(G1961), .ZN(n945) );
  NAND2_X1 U781 ( .A1(n736), .A2(n945), .ZN(n692) );
  INV_X1 U782 ( .A(n736), .ZN(n716) );
  XNOR2_X1 U783 ( .A(G2078), .B(KEYINPUT25), .ZN(n1009) );
  NAND2_X1 U784 ( .A1(n716), .A2(n1009), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n727) );
  NOR2_X1 U786 ( .A1(G171), .A2(n727), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U788 ( .A(n696), .B(n695), .ZN(n732) );
  INV_X1 U789 ( .A(G1996), .ZN(n697) );
  XOR2_X1 U790 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n698) );
  XNOR2_X1 U791 ( .A(n699), .B(n698), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n736), .A2(G1341), .ZN(n704) );
  INV_X1 U793 ( .A(n704), .ZN(n700) );
  NOR2_X1 U794 ( .A1(n938), .A2(n700), .ZN(n701) );
  AND2_X1 U795 ( .A1(n705), .A2(n701), .ZN(n702) );
  NOR2_X1 U796 ( .A1(n702), .A2(n922), .ZN(n703) );
  XNOR2_X1 U797 ( .A(n703), .B(KEYINPUT93), .ZN(n714) );
  NAND2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U799 ( .A1(n938), .A2(n706), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n707), .A2(n922), .ZN(n712) );
  INV_X1 U801 ( .A(G2067), .ZN(n1003) );
  NOR2_X1 U802 ( .A1(n736), .A2(n1003), .ZN(n708) );
  XOR2_X1 U803 ( .A(n708), .B(KEYINPUT92), .Z(n710) );
  NAND2_X1 U804 ( .A1(n736), .A2(G1348), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n720) );
  NAND2_X1 U808 ( .A1(n716), .A2(G2072), .ZN(n715) );
  XNOR2_X1 U809 ( .A(n715), .B(KEYINPUT27), .ZN(n718) );
  INV_X1 U810 ( .A(G1956), .ZN(n946) );
  NOR2_X1 U811 ( .A1(n946), .A2(n716), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n928), .A2(n722), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U815 ( .A(n721), .B(KEYINPUT94), .ZN(n725) );
  OR2_X1 U816 ( .A1(n928), .A2(n722), .ZN(n723) );
  XNOR2_X1 U817 ( .A(KEYINPUT28), .B(n723), .ZN(n724) );
  NAND2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U819 ( .A(n726), .B(KEYINPUT29), .ZN(n729) );
  AND2_X1 U820 ( .A1(G171), .A2(n727), .ZN(n728) );
  NOR2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U822 ( .A(KEYINPUT95), .B(n730), .Z(n731) );
  NOR2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U824 ( .A(KEYINPUT97), .B(n733), .ZN(n748) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n748), .A2(n734), .ZN(n743) );
  INV_X1 U827 ( .A(G8), .ZN(n741) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n805), .ZN(n735) );
  XNOR2_X1 U829 ( .A(n735), .B(KEYINPUT98), .ZN(n738) );
  NOR2_X1 U830 ( .A1(n736), .A2(G2090), .ZN(n737) );
  NOR2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n739), .A2(G303), .ZN(n740) );
  OR2_X1 U833 ( .A1(n741), .A2(n740), .ZN(n742) );
  AND2_X1 U834 ( .A1(n743), .A2(n742), .ZN(n745) );
  XOR2_X1 U835 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n744) );
  XNOR2_X1 U836 ( .A(n745), .B(n744), .ZN(n754) );
  NAND2_X1 U837 ( .A1(G8), .A2(n746), .ZN(n747) );
  XOR2_X1 U838 ( .A(KEYINPUT91), .B(n747), .Z(n752) );
  INV_X1 U839 ( .A(n748), .ZN(n749) );
  NOR2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n799) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n790) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n790), .A2(n755), .ZN(n932) );
  NAND2_X1 U846 ( .A1(n799), .A2(n932), .ZN(n756) );
  XNOR2_X1 U847 ( .A(n756), .B(KEYINPUT100), .ZN(n796) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n927) );
  INV_X1 U849 ( .A(n927), .ZN(n757) );
  NOR2_X1 U850 ( .A1(n805), .A2(n757), .ZN(n794) );
  XOR2_X1 U851 ( .A(G1981), .B(G305), .Z(n919) );
  NOR2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n819) );
  NAND2_X1 U853 ( .A1(G107), .A2(n884), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G95), .A2(n888), .ZN(n761) );
  NAND2_X1 U855 ( .A1(G119), .A2(n883), .ZN(n760) );
  NAND2_X1 U856 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U857 ( .A1(G131), .A2(n891), .ZN(n762) );
  XNOR2_X1 U858 ( .A(KEYINPUT87), .B(n762), .ZN(n763) );
  NOR2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U860 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U861 ( .A(n767), .B(KEYINPUT88), .ZN(n879) );
  NAND2_X1 U862 ( .A1(G1991), .A2(n879), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G105), .A2(n888), .ZN(n768) );
  XNOR2_X1 U864 ( .A(n768), .B(KEYINPUT38), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n884), .A2(G117), .ZN(n770) );
  NAND2_X1 U866 ( .A1(G141), .A2(n891), .ZN(n769) );
  NAND2_X1 U867 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U868 ( .A1(G129), .A2(n883), .ZN(n771) );
  XNOR2_X1 U869 ( .A(KEYINPUT89), .B(n771), .ZN(n772) );
  NOR2_X1 U870 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U871 ( .A1(n775), .A2(n774), .ZN(n901) );
  NAND2_X1 U872 ( .A1(G1996), .A2(n901), .ZN(n776) );
  NAND2_X1 U873 ( .A1(n777), .A2(n776), .ZN(n978) );
  NAND2_X1 U874 ( .A1(n819), .A2(n978), .ZN(n811) );
  XNOR2_X1 U875 ( .A(n811), .B(KEYINPUT90), .ZN(n779) );
  XNOR2_X1 U876 ( .A(G1986), .B(G290), .ZN(n934) );
  NAND2_X1 U877 ( .A1(n934), .A2(n819), .ZN(n778) );
  AND2_X1 U878 ( .A1(n779), .A2(n778), .ZN(n807) );
  AND2_X1 U879 ( .A1(n919), .A2(n807), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n888), .A2(G104), .ZN(n781) );
  NAND2_X1 U881 ( .A1(G140), .A2(n891), .ZN(n780) );
  NAND2_X1 U882 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U883 ( .A(KEYINPUT34), .B(n782), .ZN(n787) );
  NAND2_X1 U884 ( .A1(G128), .A2(n883), .ZN(n784) );
  NAND2_X1 U885 ( .A1(G116), .A2(n884), .ZN(n783) );
  NAND2_X1 U886 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U887 ( .A(KEYINPUT35), .B(n785), .Z(n786) );
  NOR2_X1 U888 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U889 ( .A(KEYINPUT36), .B(n788), .ZN(n907) );
  XNOR2_X1 U890 ( .A(KEYINPUT37), .B(G2067), .ZN(n817) );
  NOR2_X1 U891 ( .A1(n907), .A2(n817), .ZN(n990) );
  NAND2_X1 U892 ( .A1(n819), .A2(n990), .ZN(n816) );
  NAND2_X1 U893 ( .A1(n789), .A2(n816), .ZN(n793) );
  NAND2_X1 U894 ( .A1(n790), .A2(KEYINPUT33), .ZN(n791) );
  NOR2_X1 U895 ( .A1(n791), .A2(n805), .ZN(n792) );
  NOR2_X1 U896 ( .A1(n793), .A2(n792), .ZN(n821) );
  AND2_X1 U897 ( .A1(n794), .A2(n821), .ZN(n795) );
  NAND2_X1 U898 ( .A1(n796), .A2(n795), .ZN(n829) );
  NOR2_X1 U899 ( .A1(G2090), .A2(G303), .ZN(n797) );
  NAND2_X1 U900 ( .A1(G8), .A2(n797), .ZN(n798) );
  NAND2_X1 U901 ( .A1(n799), .A2(n798), .ZN(n802) );
  AND2_X1 U902 ( .A1(n805), .A2(n807), .ZN(n800) );
  AND2_X1 U903 ( .A1(n800), .A2(n816), .ZN(n801) );
  AND2_X1 U904 ( .A1(n802), .A2(n801), .ZN(n827) );
  NOR2_X1 U905 ( .A1(G1981), .A2(G305), .ZN(n803) );
  XOR2_X1 U906 ( .A(n803), .B(KEYINPUT24), .Z(n804) );
  NOR2_X1 U907 ( .A1(n805), .A2(n804), .ZN(n806) );
  AND2_X1 U908 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U909 ( .A1(n816), .A2(n808), .ZN(n825) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U911 ( .A1(n879), .A2(G1991), .ZN(n979) );
  NOR2_X1 U912 ( .A1(n809), .A2(n979), .ZN(n810) );
  XNOR2_X1 U913 ( .A(n810), .B(KEYINPUT101), .ZN(n812) );
  NAND2_X1 U914 ( .A1(n812), .A2(n811), .ZN(n813) );
  OR2_X1 U915 ( .A1(n901), .A2(G1996), .ZN(n982) );
  NAND2_X1 U916 ( .A1(n813), .A2(n982), .ZN(n814) );
  XOR2_X1 U917 ( .A(KEYINPUT39), .B(n814), .Z(n815) );
  NAND2_X1 U918 ( .A1(n816), .A2(n815), .ZN(n818) );
  NAND2_X1 U919 ( .A1(n907), .A2(n817), .ZN(n987) );
  NAND2_X1 U920 ( .A1(n818), .A2(n987), .ZN(n820) );
  NAND2_X1 U921 ( .A1(n820), .A2(n819), .ZN(n823) );
  NAND2_X1 U922 ( .A1(n821), .A2(KEYINPUT33), .ZN(n822) );
  AND2_X1 U923 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U924 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U925 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U930 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U932 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(KEYINPUT105), .B(n835), .Z(G188) );
  XOR2_X1 U934 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  XOR2_X1 U935 ( .A(n836), .B(G286), .Z(n838) );
  XNOR2_X1 U936 ( .A(G171), .B(n922), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n839), .B(n938), .ZN(n840) );
  NOR2_X1 U939 ( .A1(G37), .A2(n840), .ZN(G397) );
  XOR2_X1 U940 ( .A(KEYINPUT41), .B(G1961), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n843), .B(KEYINPUT109), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1981), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1956), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U950 ( .A(KEYINPUT108), .B(G2474), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U952 ( .A(KEYINPUT107), .B(G2072), .Z(n853) );
  XNOR2_X1 U953 ( .A(G2084), .B(G2078), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n854), .B(G2100), .Z(n856) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2090), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(G2096), .B(G2678), .Z(n858) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U961 ( .A(n860), .B(n859), .Z(G227) );
  NAND2_X1 U962 ( .A1(G100), .A2(n888), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G112), .A2(n884), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G124), .A2(n883), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n863), .B(KEYINPUT44), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n864), .B(KEYINPUT110), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G136), .A2(n891), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U970 ( .A(KEYINPUT111), .B(n867), .Z(n868) );
  NOR2_X1 U971 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U972 ( .A1(n888), .A2(G106), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G142), .A2(n891), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n872), .B(KEYINPUT45), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G130), .A2(n883), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n884), .A2(G118), .ZN(n875) );
  XOR2_X1 U979 ( .A(KEYINPUT112), .B(n875), .Z(n876) );
  NOR2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n905) );
  XNOR2_X1 U982 ( .A(G160), .B(n977), .ZN(n899) );
  XOR2_X1 U983 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n881) );
  XNOR2_X1 U984 ( .A(KEYINPUT118), .B(KEYINPUT117), .ZN(n880) );
  XNOR2_X1 U985 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U986 ( .A(n882), .B(KEYINPUT48), .Z(n897) );
  NAND2_X1 U987 ( .A1(G127), .A2(n883), .ZN(n886) );
  NAND2_X1 U988 ( .A1(G115), .A2(n884), .ZN(n885) );
  NAND2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n887), .B(KEYINPUT47), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G103), .A2(n888), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n894) );
  NAND2_X1 U993 ( .A1(G139), .A2(n891), .ZN(n892) );
  XNOR2_X1 U994 ( .A(KEYINPUT115), .B(n892), .ZN(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U996 ( .A(KEYINPUT116), .B(n895), .Z(n972) );
  XNOR2_X1 U997 ( .A(n972), .B(KEYINPUT46), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U1000 ( .A(n900), .B(G162), .Z(n903) );
  XOR2_X1 U1001 ( .A(G164), .B(n901), .Z(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n907), .B(n906), .Z(n908) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n908), .ZN(n909) );
  XOR2_X1 U1006 ( .A(KEYINPUT119), .B(n909), .Z(G395) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(G397), .A2(n911), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(n918), .A2(G401), .ZN(n912) );
  XOR2_X1 U1011 ( .A(KEYINPUT120), .B(n912), .Z(n913) );
  NOR2_X1 U1012 ( .A1(G395), .A2(n913), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(G225) );
  XNOR2_X1 U1014 ( .A(KEYINPUT121), .B(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(G325) );
  INV_X1 U1019 ( .A(G325), .ZN(G261) );
  INV_X1 U1020 ( .A(n918), .ZN(G319) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1022 ( .A(G16), .B(KEYINPUT56), .ZN(n944) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G168), .ZN(n920) );
  NAND2_X1 U1024 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1025 ( .A(n921), .B(KEYINPUT57), .ZN(n942) );
  XNOR2_X1 U1026 ( .A(G1348), .B(n922), .ZN(n923) );
  XNOR2_X1 U1027 ( .A(n923), .B(KEYINPUT125), .ZN(n925) );
  XNOR2_X1 U1028 ( .A(G171), .B(n945), .ZN(n924) );
  NOR2_X1 U1029 ( .A1(n925), .A2(n924), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(G1971), .A2(G303), .ZN(n926) );
  NAND2_X1 U1031 ( .A1(n927), .A2(n926), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(n946), .B(n928), .ZN(n929) );
  NOR2_X1 U1033 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(n935), .B(KEYINPUT126), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n940) );
  XNOR2_X1 U1038 ( .A(G1341), .B(n938), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n971) );
  INV_X1 U1042 ( .A(G16), .ZN(n969) );
  XNOR2_X1 U1043 ( .A(G5), .B(n945), .ZN(n958) );
  XNOR2_X1 U1044 ( .A(G20), .B(n946), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G1341), .B(G19), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G6), .B(G1981), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1049 ( .A(KEYINPUT59), .B(G1348), .Z(n951) );
  XNOR2_X1 U1050 ( .A(G4), .B(n951), .ZN(n952) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1052 ( .A(KEYINPUT60), .B(n954), .Z(n956) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G21), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(G1986), .B(KEYINPUT127), .ZN(n961) );
  XNOR2_X1 U1060 ( .A(n961), .B(G24), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(KEYINPUT58), .B(n964), .ZN(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(KEYINPUT61), .B(n967), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n1023) );
  XOR2_X1 U1067 ( .A(G164), .B(G2078), .Z(n974) );
  XNOR2_X1 U1068 ( .A(G2072), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1070 ( .A(KEYINPUT50), .B(n975), .Z(n993) );
  XOR2_X1 U1071 ( .A(G2084), .B(G160), .Z(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G162), .B(G2090), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT51), .B(n984), .Z(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1081 ( .A(KEYINPUT122), .B(n991), .Z(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1083 ( .A(KEYINPUT52), .B(n994), .Z(n995) );
  NOR2_X1 U1084 ( .A1(KEYINPUT55), .A2(n995), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(n996), .B(KEYINPUT123), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n997), .A2(G29), .ZN(n1021) );
  XOR2_X1 U1087 ( .A(G2090), .B(G35), .Z(n1000) );
  XOR2_X1 U1088 ( .A(G34), .B(KEYINPUT54), .Z(n998) );
  XNOR2_X1 U1089 ( .A(G2084), .B(n998), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1014) );
  XNOR2_X1 U1091 ( .A(G1996), .B(G32), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G33), .B(G2072), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(G26), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(G28), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(G25), .B(G1991), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(G27), .B(n1009), .Z(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1012), .B(KEYINPUT53), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(KEYINPUT55), .B(n1015), .ZN(n1017) );
  INV_X1 U1104 ( .A(G29), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(G11), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT124), .B(n1019), .Z(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(n1024), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

