//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(KEYINPUT67), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n467), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n471), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n469), .A2(G2105), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n479), .A2(KEYINPUT68), .A3(G101), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT68), .B1(new_n479), .B2(G101), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n477), .A2(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n475), .A2(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n476), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n465), .A2(new_n466), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n463), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OAI22_X1  g071(.A1(new_n484), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n467), .A2(new_n472), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n463), .C1(new_n465), .C2(new_n466), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n500), .A2(new_n501), .B1(KEYINPUT4), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n467), .A2(new_n472), .A3(KEYINPUT69), .A4(new_n499), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n497), .B1(new_n503), .B2(new_n504), .ZN(G164));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT70), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(new_n506), .ZN(new_n514));
  AOI22_X1  g089(.A1(G50), .A2(new_n513), .B1(new_n514), .B2(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n509), .A2(KEYINPUT70), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n511), .A2(new_n506), .ZN(new_n523));
  OAI221_X1 g098(.A(new_n520), .B1(new_n512), .B2(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT71), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(G168));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n523), .A2(new_n528), .B1(new_n512), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n508), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(new_n532), .ZN(G171));
  INV_X1    g108(.A(G81), .ZN(new_n534));
  INV_X1    g109(.A(G43), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n523), .A2(new_n534), .B1(new_n512), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n508), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  NAND4_X1  g115(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(G188));
  NAND3_X1  g119(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT9), .B1(new_n545), .B2(KEYINPUT72), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(KEYINPUT72), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(KEYINPUT73), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n508), .B1(new_n549), .B2(KEYINPUT73), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n550), .A2(new_n551), .B1(G91), .B2(new_n514), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G299));
  OR2_X1    g128(.A1(new_n530), .A2(new_n532), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT74), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n556));
  NAND2_X1  g131(.A1(G171), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(G301));
  INV_X1    g134(.A(G168), .ZN(G286));
  INV_X1    g135(.A(G166), .ZN(G303));
  NAND2_X1  g136(.A1(new_n514), .A2(G87), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n506), .A2(G74), .ZN(new_n564));
  AOI22_X1  g139(.A1(G49), .A2(new_n513), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(G288));
  INV_X1    g141(.A(G86), .ZN(new_n567));
  INV_X1    g142(.A(G48), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n523), .A2(new_n567), .B1(new_n512), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n508), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G305));
  INV_X1    g148(.A(G85), .ZN(new_n574));
  INV_X1    g149(.A(G47), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n523), .A2(new_n574), .B1(new_n512), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n508), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G290));
  AND3_X1   g157(.A1(G301), .A2(KEYINPUT77), .A3(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n514), .A2(G92), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT10), .Z(new_n585));
  NAND2_X1  g160(.A1(new_n506), .A2(G66), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n508), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G54), .B2(new_n513), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT78), .ZN(new_n591));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT77), .B1(G301), .B2(G868), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n583), .B1(new_n593), .B2(new_n594), .ZN(G284));
  AOI21_X1  g170(.A(new_n583), .B1(new_n593), .B2(new_n594), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(G299), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G297));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G280));
  AND2_X1   g175(.A1(new_n585), .A2(new_n589), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT78), .ZN(new_n602));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G860), .ZN(G148));
  INV_X1    g179(.A(new_n539), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(new_n592), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n591), .A2(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n592), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n488), .A2(G135), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT79), .Z(new_n611));
  INV_X1    g186(.A(G111), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n612), .A2(KEYINPUT80), .A3(G2105), .ZN(new_n613));
  AOI21_X1  g188(.A(KEYINPUT80), .B1(new_n612), .B2(G2105), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n485), .A2(G123), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT81), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2096), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n467), .A2(new_n472), .A3(new_n479), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT82), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2430), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(KEYINPUT14), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n632), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  OAI21_X1  g213(.A(G14), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT84), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n644), .B(KEYINPUT17), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n646), .B1(new_n641), .B2(new_n647), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n648), .B(new_n651), .C1(new_n652), .C2(new_n643), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT85), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n658), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n658), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1981), .B(G1986), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  NAND2_X1  g249(.A1(new_n619), .A2(G29), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT31), .B(G11), .ZN(new_n676));
  INV_X1    g251(.A(G28), .ZN(new_n677));
  OAI21_X1  g252(.A(KEYINPUT96), .B1(new_n677), .B2(KEYINPUT30), .ZN(new_n678));
  AOI21_X1  g253(.A(G29), .B1(new_n677), .B2(KEYINPUT30), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n677), .A2(KEYINPUT96), .A3(KEYINPUT30), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n676), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NOR2_X1   g258(.A1(G171), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G5), .B2(new_n683), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n682), .B1(new_n686), .B2(G1961), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(G21), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G168), .B2(new_n683), .ZN(new_n689));
  INV_X1    g264(.A(G1966), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n675), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT97), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n683), .A2(G4), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n602), .B2(new_n683), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1348), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G26), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  OR2_X1    g274(.A1(G104), .A2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n700), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT93), .ZN(new_n702));
  INV_X1    g277(.A(G128), .ZN(new_n703));
  INV_X1    g278(.A(G140), .ZN(new_n704));
  OAI22_X1  g279(.A1(new_n703), .A2(new_n484), .B1(new_n477), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n699), .B1(new_n706), .B2(new_n697), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2067), .ZN(new_n708));
  INV_X1    g283(.A(G1961), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n685), .ZN(new_n710));
  INV_X1    g285(.A(G34), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(KEYINPUT24), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(KEYINPUT24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n697), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G160), .B2(new_n697), .ZN(new_n715));
  INV_X1    g290(.A(G2084), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n683), .A2(G19), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT92), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n539), .B2(new_n683), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1341), .Z(new_n721));
  NOR2_X1   g296(.A1(G29), .A2(G35), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G162), .B2(G29), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT29), .B(G2090), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n710), .A2(new_n717), .A3(new_n721), .A4(new_n725), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n693), .A2(new_n696), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n697), .A2(G27), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G164), .B2(new_n697), .ZN(new_n729));
  INV_X1    g304(.A(G2078), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT26), .Z(new_n733));
  INV_X1    g308(.A(G129), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n484), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n488), .A2(G141), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n479), .A2(G105), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G29), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT95), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G29), .B2(G32), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(KEYINPUT95), .B2(new_n740), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n683), .A2(G20), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G299), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(G1956), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n753));
  OR3_X1    g328(.A1(new_n753), .A2(G29), .A3(G33), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(G29), .B2(G33), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n467), .A2(new_n472), .A3(G127), .ZN(new_n756));
  INV_X1    g331(.A(G115), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n469), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G2105), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n488), .A2(G139), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n754), .B(new_n755), .C1(new_n765), .C2(new_n697), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G2072), .Z(new_n767));
  NOR3_X1   g342(.A1(new_n746), .A2(new_n752), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n727), .A2(new_n731), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n683), .A2(G24), .ZN(new_n770));
  INV_X1    g345(.A(G290), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n683), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1986), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n697), .A2(G25), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT87), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n485), .A2(G119), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n488), .A2(G131), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n463), .A2(G107), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(KEYINPUT88), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT88), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n775), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT35), .B(G1991), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT89), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n784), .B(new_n786), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n683), .A2(G23), .ZN(new_n788));
  INV_X1    g363(.A(G288), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n683), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT33), .B(G1976), .Z(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n683), .A2(G6), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n572), .B2(new_n683), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT32), .B(G1981), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT90), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n790), .A2(new_n791), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n792), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n683), .A2(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n683), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G1971), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(G1971), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n802), .A2(KEYINPUT91), .A3(new_n803), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n799), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n773), .B(new_n787), .C1(new_n808), .C2(KEYINPUT34), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n810));
  OR3_X1    g385(.A1(new_n809), .A2(new_n810), .A3(KEYINPUT36), .ZN(new_n811));
  OAI21_X1  g386(.A(KEYINPUT36), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n769), .B1(new_n811), .B2(new_n812), .ZN(G311));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n814));
  XNOR2_X1  g389(.A(G311), .B(new_n814), .ZN(G150));
  NOR2_X1   g390(.A1(new_n591), .A2(new_n603), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT38), .ZN(new_n817));
  INV_X1    g392(.A(G93), .ZN(new_n818));
  INV_X1    g393(.A(G55), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n523), .A2(new_n818), .B1(new_n512), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n508), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n539), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n817), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n827));
  AOI21_X1  g402(.A(G860), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  OAI21_X1  g404(.A(G860), .B1(new_n820), .B2(new_n822), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(G145));
  INV_X1    g407(.A(new_n765), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n500), .A2(new_n501), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n504), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n497), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n706), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n834), .B1(new_n840), .B2(new_n739), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n739), .B2(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n833), .A2(KEYINPUT100), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n485), .A2(G130), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n463), .A2(G118), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n488), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(new_n622), .Z(new_n850));
  INV_X1    g425(.A(new_n783), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n844), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n844), .A2(new_n852), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n619), .B(G162), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G160), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n853), .B2(new_n854), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g436(.A(new_n607), .B(new_n824), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n601), .B2(G299), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n598), .A2(KEYINPUT102), .A3(new_n590), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n601), .A2(G299), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT101), .B1(new_n601), .B2(G299), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n598), .A2(new_n590), .A3(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n865), .B(new_n864), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n873), .B2(new_n868), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n862), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n862), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT42), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n875), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n771), .A2(new_n789), .ZN(new_n882));
  NAND2_X1  g457(.A1(G290), .A2(G288), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(KEYINPUT103), .A3(new_n883), .ZN(new_n887));
  XNOR2_X1  g462(.A(G166), .B(new_n572), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G166), .B(G305), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n884), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n878), .B2(new_n879), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n880), .B1(new_n875), .B2(new_n877), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n881), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n881), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(G868), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(G868), .B2(new_n823), .ZN(G295));
  OAI21_X1  g474(.A(new_n898), .B1(G868), .B2(new_n823), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n901));
  OR3_X1    g476(.A1(G168), .A2(KEYINPUT105), .A3(new_n554), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT105), .B1(G168), .B2(new_n554), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n555), .A2(G168), .A3(new_n557), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n825), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n902), .A2(new_n824), .A3(new_n903), .A4(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n873), .A2(new_n906), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n910), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n874), .A2(new_n908), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n914), .B2(new_n892), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n906), .A3(new_n912), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n867), .A2(KEYINPUT41), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n917), .B(new_n918), .C1(KEYINPUT41), .C2(new_n873), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n909), .A2(new_n907), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n915), .B(new_n916), .C1(new_n892), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n874), .A2(new_n908), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n909), .A2(new_n913), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n893), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n916), .B1(new_n915), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI211_X1 g504(.A(KEYINPUT107), .B(new_n916), .C1(new_n915), .C2(new_n926), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n901), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n892), .A2(new_n923), .A3(new_n924), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n858), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n892), .B1(new_n919), .B2(new_n920), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n915), .A2(new_n916), .A3(new_n926), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT44), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n931), .B1(new_n939), .B2(new_n940), .ZN(G397));
  INV_X1    g516(.A(KEYINPUT119), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT115), .ZN(new_n943));
  INV_X1    g518(.A(G40), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n475), .A2(new_n482), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n837), .B2(new_n838), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT50), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n943), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n839), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n943), .B1(new_n952), .B2(new_n945), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n751), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(G299), .B(KEYINPUT57), .Z(new_n955));
  NAND2_X1  g530(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n945), .B1(new_n946), .B2(KEYINPUT45), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT56), .B(G2072), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n954), .A2(new_n955), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT118), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n955), .B1(new_n954), .B2(new_n961), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n954), .A2(new_n961), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT118), .ZN(new_n967));
  INV_X1    g542(.A(new_n955), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n942), .B1(new_n965), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT120), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n962), .A2(KEYINPUT61), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n964), .ZN(new_n975));
  INV_X1    g550(.A(new_n964), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n976), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n962), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT59), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n839), .A2(new_n949), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n983), .A3(new_n945), .A4(new_n956), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n946), .A2(new_n945), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT58), .B(G1341), .Z(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n979), .B1(new_n988), .B2(new_n539), .ZN(new_n989));
  AOI211_X1 g564(.A(KEYINPUT59), .B(new_n605), .C1(new_n984), .C2(new_n987), .ZN(new_n990));
  INV_X1    g565(.A(G2067), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n946), .A2(new_n991), .A3(new_n945), .ZN(new_n992));
  INV_X1    g567(.A(new_n945), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n952), .A2(new_n950), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n980), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n992), .B1(new_n997), .B2(G1348), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n590), .A2(KEYINPUT60), .ZN(new_n999));
  OAI22_X1  g574(.A1(new_n989), .A2(new_n990), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n601), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n590), .B(new_n992), .C1(new_n997), .C2(G1348), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(KEYINPUT60), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT61), .B1(new_n964), .B2(new_n967), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1005), .B(KEYINPUT119), .C1(new_n964), .C2(new_n963), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n972), .A2(new_n978), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n964), .B1(new_n1001), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1008), .B2(new_n1001), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n962), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n995), .A2(new_n996), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n945), .A2(new_n716), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n690), .B1(new_n957), .B2(new_n958), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(G168), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1014), .B1(new_n995), .B2(new_n996), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n993), .B1(new_n980), .B2(new_n981), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1966), .B1(new_n1020), .B2(new_n956), .ZN(new_n1021));
  OAI21_X1  g596(.A(G286), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1022), .A3(G8), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT51), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1018), .A2(new_n1025), .A3(G8), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1020), .A2(new_n730), .A3(new_n956), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n959), .A2(KEYINPUT53), .A3(new_n730), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n997), .A2(G1961), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(G301), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(G171), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(KEYINPUT54), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1027), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1040));
  AOI21_X1  g615(.A(G301), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1032), .A2(new_n1034), .A3(new_n558), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT122), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT122), .B(new_n1040), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1039), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n945), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n995), .B2(new_n996), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1050), .A2(KEYINPUT111), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n1052), .B(new_n1049), .C1(new_n995), .C2(new_n996), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1971), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n957), .B2(new_n958), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G166), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT55), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1057), .A2(new_n1058), .A3(G8), .A4(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1056), .B1(new_n1050), .B2(KEYINPUT111), .ZN(new_n1063));
  OAI211_X1 g638(.A(G8), .B(new_n1061), .C1(new_n1063), .C2(new_n1053), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT112), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n571), .B1(new_n569), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1067), .B2(new_n569), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(G1981), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT114), .ZN(new_n1071));
  OR2_X1    g646(.A1(G305), .A2(G1981), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1073), .A3(G1981), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1071), .A2(KEYINPUT49), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n985), .A2(G8), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G288), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT52), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1080), .B(new_n1085), .C1(new_n1082), .C2(G288), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1081), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1061), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n951), .A2(new_n953), .A3(G2090), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1056), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT116), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n953), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1092), .A2(new_n1048), .A3(new_n950), .A4(new_n948), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n1056), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(G8), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1087), .B1(new_n1088), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1066), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1012), .A2(new_n1047), .A3(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1081), .A2(new_n1082), .A3(new_n789), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1072), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1080), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1066), .B2(new_n1087), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT123), .B1(new_n1027), .B2(KEYINPUT62), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1106), .B(new_n1107), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1024), .A2(new_n1107), .A3(new_n1026), .ZN(new_n1110));
  AND4_X1   g685(.A1(new_n1066), .A2(new_n1097), .A3(new_n1110), .A4(new_n1041), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1104), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1059), .B(G286), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1098), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1061), .B1(new_n1057), .B2(G8), .ZN(new_n1117));
  NOR4_X1   g692(.A1(new_n1117), .A2(new_n1087), .A3(new_n1115), .A4(new_n1113), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n1066), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1100), .A2(new_n1112), .A3(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n706), .B(new_n991), .ZN(new_n1122));
  INV_X1    g697(.A(new_n739), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(G1996), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n980), .A2(new_n981), .A3(new_n945), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(G1996), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT109), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1129), .B2(new_n739), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n783), .B(new_n786), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1125), .ZN(new_n1133));
  XNOR2_X1  g708(.A(G290), .B(G1986), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1121), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1123), .B2(new_n1122), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1128), .A2(KEYINPUT46), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1128), .A2(KEYINPUT46), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1144), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n851), .A2(new_n786), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT124), .Z(new_n1149));
  AOI22_X1  g724(.A1(new_n1130), .A2(new_n1149), .B1(new_n991), .B2(new_n706), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1125), .A2(G290), .A3(G1986), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT127), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT48), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1150), .A2(new_n1125), .B1(new_n1132), .B2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1146), .A2(new_n1147), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1136), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g731(.A1(G229), .A2(new_n461), .A3(G227), .A4(G401), .ZN(new_n1158));
  OAI211_X1 g732(.A(new_n860), .B(new_n1158), .C1(new_n929), .C2(new_n930), .ZN(G225));
  INV_X1    g733(.A(G225), .ZN(G308));
endmodule


