//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G250), .B(G257), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  INV_X1    g0041(.A(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n218), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT68), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT68), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AND3_X1   g0053(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n205), .B(G274), .C1(new_n255), .C2(new_n214), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT69), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  INV_X1    g0058(.A(new_n214), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT69), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .A4(new_n205), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G226), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n265), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT70), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1698), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G222), .ZN(new_n278));
  INV_X1    g0078(.A(G77), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n276), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(G1698), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n278), .B1(new_n279), .B2(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n267), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n272), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n270), .A2(new_n271), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G190), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n214), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n242), .B1(new_n205), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(new_n297), .B1(new_n242), .B2(new_n293), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT8), .B(G58), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n206), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G150), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n299), .A2(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n206), .B1(new_n201), .B2(new_n242), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n298), .B(new_n306), .C1(KEYINPUT72), .C2(KEYINPUT9), .ZN(new_n307));
  NAND2_X1  g0107(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n308));
  XOR2_X1   g0108(.A(new_n307), .B(new_n308), .Z(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n289), .B(new_n309), .C1(new_n310), .C2(new_n288), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n288), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n298), .A2(new_n306), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n314), .B(new_n315), .C1(G169), .C2(new_n288), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G58), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n218), .ZN(new_n319));
  OAI21_X1  g0119(.A(G20), .B1(new_n319), .B2(new_n201), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n302), .A2(G159), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n275), .A2(new_n206), .A3(new_n276), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n276), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n326), .A2(KEYINPUT75), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(G68), .B1(new_n326), .B2(KEYINPUT75), .ZN(new_n329));
  OAI211_X1 g0129(.A(KEYINPUT16), .B(new_n323), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n218), .B1(new_n326), .B2(new_n327), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n322), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n295), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n299), .B1(new_n205), .B2(G20), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n296), .A2(new_n335), .B1(new_n293), .B2(new_n299), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n267), .A2(G232), .A3(new_n268), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G87), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n266), .A2(G1698), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G223), .B2(G1698), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n339), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n345), .B2(new_n284), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n265), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G169), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n265), .A2(new_n346), .A3(G179), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n337), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT18), .ZN(new_n352));
  INV_X1    g0152(.A(new_n336), .ZN(new_n353));
  INV_X1    g0153(.A(new_n295), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT7), .B1(new_n344), .B2(new_n206), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT75), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n218), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n326), .A2(KEYINPUT75), .A3(new_n327), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n322), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n354), .B1(new_n359), .B2(KEYINPUT16), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n353), .B1(new_n360), .B2(new_n333), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n347), .A2(new_n310), .ZN(new_n362));
  INV_X1    g0162(.A(G190), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n265), .A2(new_n346), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n361), .A2(KEYINPUT76), .A3(KEYINPUT17), .A4(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n365), .A2(new_n334), .A3(KEYINPUT76), .A4(new_n336), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT17), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n337), .A2(new_n370), .A3(new_n350), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n352), .A2(new_n366), .A3(new_n369), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G1698), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n280), .A2(G232), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n375), .B1(new_n376), .B2(new_n280), .C1(new_n282), .C2(new_n217), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n284), .ZN(new_n378));
  INV_X1    g0178(.A(G244), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n378), .B(new_n265), .C1(new_n379), .C2(new_n269), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(G179), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n299), .A2(new_n303), .B1(new_n206), .B2(new_n279), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n300), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n295), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT71), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n205), .A2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G77), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n296), .A2(new_n389), .B1(new_n279), .B2(new_n293), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G169), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n380), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n381), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n380), .A2(G200), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n395), .B(new_n396), .C1(new_n363), .C2(new_n380), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  OR3_X1    g0198(.A1(new_n292), .A2(KEYINPUT73), .A3(G68), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT73), .B1(new_n292), .B2(G68), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(KEYINPUT12), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n296), .A2(G68), .A3(new_n387), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n400), .A2(KEYINPUT12), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n303), .A2(new_n242), .B1(new_n206), .B2(G68), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n300), .A2(new_n279), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n295), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT11), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT14), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n267), .A2(G238), .A3(new_n268), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n265), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G97), .ZN(new_n417));
  INV_X1    g0217(.A(new_n277), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n416), .B(new_n417), .C1(new_n418), .C2(new_n266), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n284), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n414), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n415), .B1(new_n414), .B2(new_n420), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n412), .B(G169), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n423), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n421), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n424), .B1(new_n313), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n412), .B1(new_n426), .B2(G169), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n411), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n411), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(G200), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n430), .B(new_n431), .C1(new_n363), .C2(new_n426), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AND4_X1   g0234(.A1(new_n317), .A2(new_n373), .A3(new_n398), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT23), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n206), .B2(G107), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n376), .A2(KEYINPUT23), .A3(G20), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(KEYINPUT78), .A2(G116), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(KEYINPUT78), .A2(G116), .ZN(new_n442));
  OAI21_X1  g0242(.A(G33), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n439), .B1(new_n443), .B2(G20), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n206), .B(G87), .C1(new_n342), .C2(new_n343), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT22), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(new_n206), .A3(G87), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT84), .B1(new_n344), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT84), .ZN(new_n450));
  INV_X1    g0250(.A(G87), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n451), .A2(KEYINPUT22), .A3(G20), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n280), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  AOI221_X4 g0253(.A(KEYINPUT85), .B1(new_n446), .B2(KEYINPUT22), .C1(new_n449), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT85), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n449), .A2(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n446), .A2(KEYINPUT22), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n445), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT24), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(KEYINPUT24), .B(new_n445), .C1(new_n454), .C2(new_n458), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(new_n295), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n293), .A2(new_n376), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n464), .B2(new_n465), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n274), .A2(G1), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n293), .A2(new_n295), .A3(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n466), .A2(new_n468), .B1(G107), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT5), .B1(new_n250), .B2(new_n252), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n253), .A2(G1), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G264), .B(new_n267), .C1(new_n472), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT88), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT68), .B(G41), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n474), .B(new_n473), .C1(new_n479), .C2(KEYINPUT5), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(KEYINPUT88), .A3(G264), .A4(new_n267), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n280), .A2(G257), .A3(G1698), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G294), .ZN(new_n483));
  INV_X1    g0283(.A(G250), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n482), .B(new_n483), .C1(new_n418), .C2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n478), .A2(new_n481), .B1(new_n485), .B2(new_n284), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n473), .A2(new_n474), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n487), .B(new_n261), .C1(KEYINPUT5), .C2(new_n479), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(G190), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n488), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G200), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n463), .A2(new_n471), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n471), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n354), .B1(new_n459), .B2(new_n460), .ZN(new_n495));
  AOI211_X1 g0295(.A(KEYINPUT87), .B(new_n494), .C1(new_n495), .C2(new_n462), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT87), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n463), .B2(new_n471), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n490), .A2(G169), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n313), .B2(new_n490), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n493), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT21), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n354), .B(new_n292), .C1(G1), .C2(new_n274), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n441), .A2(new_n442), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n504), .A2(new_n505), .B1(new_n507), .B2(new_n292), .ZN(new_n508));
  AOI21_X1  g0308(.A(G20), .B1(G33), .B2(G283), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n274), .A2(G97), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n509), .A2(new_n510), .B1(new_n294), .B2(new_n214), .ZN(new_n511));
  INV_X1    g0311(.A(new_n442), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(G20), .A3(new_n440), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT20), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT20), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT83), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n508), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G264), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n521));
  OAI211_X1 g0321(.A(G257), .B(new_n374), .C1(new_n342), .C2(new_n343), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n275), .A2(G303), .A3(new_n276), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n284), .ZN(new_n525));
  OAI211_X1 g0325(.A(G270), .B(new_n267), .C1(new_n472), .C2(new_n475), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n488), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G169), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n503), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n511), .A2(new_n513), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n511), .A2(new_n513), .A3(new_n516), .A4(KEYINPUT20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n519), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n470), .A2(G116), .B1(new_n506), .B2(new_n293), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(KEYINPUT21), .A3(G169), .A4(new_n527), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n527), .A2(G200), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n525), .A2(G190), .A3(new_n488), .A4(new_n526), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n520), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n525), .A2(G179), .A3(new_n488), .A4(new_n526), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  AND4_X1   g0343(.A1(new_n529), .A2(new_n537), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  AND2_X1   g0345(.A1(G97), .A2(G107), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n376), .A2(KEYINPUT77), .A3(KEYINPUT6), .A4(G97), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT77), .ZN(new_n550));
  NAND2_X1  g0350(.A1(KEYINPUT6), .A2(G97), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n548), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G20), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n302), .A2(G77), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n376), .B1(new_n326), .B2(new_n327), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n295), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n292), .A2(G97), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G97), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(new_n504), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(G257), .B(new_n267), .C1(new_n472), .C2(new_n475), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n488), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G283), .ZN(new_n567));
  OAI211_X1 g0367(.A(G250), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n568));
  OAI211_X1 g0368(.A(G244), .B(new_n374), .C1(new_n342), .C2(new_n343), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT4), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT4), .B1(new_n277), .B2(G244), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n284), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n392), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n566), .A2(new_n573), .A3(new_n313), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n564), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(G200), .ZN(new_n578));
  INV_X1    g0378(.A(new_n327), .ZN(new_n579));
  OAI21_X1  g0379(.A(G107), .B1(new_n355), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n554), .A3(new_n555), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n562), .B1(new_n581), .B2(new_n295), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n566), .A2(new_n573), .A3(G190), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g0385(.A1(G238), .A2(G1698), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n379), .A2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n586), .B(new_n587), .C1(new_n342), .C2(new_n343), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n443), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT79), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT79), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(new_n443), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n284), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT80), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n473), .A2(new_n258), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n484), .B1(new_n253), .B2(G1), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n267), .A3(new_n596), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n594), .B1(new_n593), .B2(new_n597), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n392), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n280), .A2(new_n206), .A3(G68), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n206), .B1(new_n417), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n547), .A2(new_n451), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n206), .A2(G33), .A3(G97), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n606), .A2(KEYINPUT81), .A3(new_n602), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT81), .B1(new_n606), .B2(new_n602), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n601), .B(new_n605), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n295), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n293), .A2(new_n383), .ZN(new_n611));
  INV_X1    g0411(.A(new_n383), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n470), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT82), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT82), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n610), .A2(new_n616), .A3(new_n611), .A4(new_n613), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n588), .A2(new_n591), .A3(new_n443), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n591), .B1(new_n588), .B2(new_n443), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n619), .A2(new_n620), .A3(new_n267), .ZN(new_n621));
  INV_X1    g0421(.A(new_n597), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT80), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n313), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n600), .A2(new_n618), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(G200), .B1(new_n598), .B2(new_n599), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n623), .A2(G190), .A3(new_n624), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n610), .A2(new_n611), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(G87), .B2(new_n470), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n544), .A2(new_n585), .A3(new_n626), .A4(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n435), .A2(new_n502), .A3(new_n632), .ZN(G372));
  INV_X1    g0433(.A(new_n394), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n432), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n429), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n369), .A3(new_n366), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n352), .A3(new_n371), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n312), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n316), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n558), .A2(new_n563), .B1(new_n574), .B2(new_n392), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT90), .B1(new_n642), .B2(new_n576), .ZN(new_n643));
  AND4_X1   g0443(.A1(KEYINPUT90), .A2(new_n564), .A3(new_n575), .A4(new_n576), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n392), .B1(new_n621), .B2(new_n622), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n618), .A2(new_n625), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n310), .B1(new_n593), .B2(new_n597), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT89), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT89), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n628), .A3(new_n630), .A4(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n645), .A2(new_n646), .A3(new_n648), .A4(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n577), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n626), .A2(new_n631), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT26), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(new_n648), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n492), .A2(new_n585), .A3(new_n648), .A4(new_n652), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n529), .A2(new_n537), .A3(new_n543), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n344), .A2(KEYINPUT84), .A3(new_n448), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n450), .B1(new_n280), .B2(new_n452), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n457), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT85), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n456), .A2(new_n455), .A3(new_n457), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n444), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n295), .B1(new_n665), .B2(KEYINPUT24), .ZN(new_n666));
  INV_X1    g0466(.A(new_n462), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n471), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n659), .B1(new_n668), .B2(new_n501), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n658), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n657), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n435), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n641), .A2(new_n672), .ZN(G369));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n291), .A2(new_n206), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(G213), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n544), .B1(new_n520), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n659), .A2(new_n536), .A3(new_n680), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(KEYINPUT91), .A3(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n683), .A2(KEYINPUT91), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n674), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n499), .A2(new_n680), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n502), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n499), .A2(new_n501), .A3(new_n680), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n668), .A2(new_n501), .A3(new_n681), .ZN(new_n695));
  INV_X1    g0495(.A(new_n659), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n680), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n502), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n694), .A2(new_n695), .A3(new_n698), .ZN(G399));
  NAND2_X1  g0499(.A1(new_n209), .A2(new_n479), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n604), .A2(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n212), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT29), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n671), .A2(new_n705), .A3(new_n681), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n652), .A2(new_n648), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT90), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n577), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n642), .A2(KEYINPUT90), .A3(new_n576), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT26), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n626), .A2(new_n631), .A3(new_n646), .A4(new_n654), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n648), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n668), .A2(KEYINPUT87), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n463), .A2(new_n497), .A3(new_n471), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n716), .A3(new_n501), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n696), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n492), .A2(new_n648), .A3(new_n652), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n577), .A2(new_n584), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT97), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n577), .A2(new_n584), .A3(KEYINPUT97), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT98), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n714), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n718), .A2(new_n725), .A3(KEYINPUT98), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n680), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n706), .B1(new_n730), .B2(new_n705), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n502), .A2(KEYINPUT96), .A3(new_n632), .A4(new_n681), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n632), .A2(new_n717), .A3(new_n492), .A4(new_n681), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT96), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT95), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n485), .A2(new_n284), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n478), .A2(new_n481), .ZN(new_n740));
  AND4_X1   g0540(.A1(new_n739), .A2(new_n740), .A3(new_n573), .A4(new_n566), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(new_n623), .A3(new_n624), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n541), .B(KEYINPUT94), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n541), .B(KEYINPUT94), .Z(new_n745));
  NOR2_X1   g0545(.A1(new_n598), .A2(new_n599), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT30), .A4(new_n741), .ZN(new_n747));
  AOI21_X1  g0547(.A(G179), .B1(new_n593), .B2(new_n597), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n490), .A2(new_n527), .A3(new_n574), .A4(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n744), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n737), .B(KEYINPUT31), .C1(new_n750), .C2(new_n680), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n680), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n755));
  NAND3_X1  g0555(.A1(new_n750), .A2(new_n680), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT95), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n751), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n674), .B1(new_n736), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n731), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n704), .B1(new_n760), .B2(G1), .ZN(G364));
  INV_X1    g0561(.A(new_n700), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n290), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n205), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n209), .A2(new_n280), .ZN(new_n767));
  INV_X1    g0567(.A(G355), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n767), .A2(new_n768), .B1(G116), .B2(new_n209), .ZN(new_n769));
  INV_X1    g0569(.A(new_n209), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n280), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n253), .B2(new_n213), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n247), .A2(new_n253), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n769), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n214), .B1(G20), .B2(new_n392), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n766), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n313), .A2(new_n310), .A3(KEYINPUT101), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(KEYINPUT101), .B1(new_n313), .B2(new_n310), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(new_n206), .A3(G190), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G329), .ZN(new_n788));
  INV_X1    g0588(.A(G283), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n206), .A2(G179), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(new_n363), .A3(G200), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n788), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n786), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n206), .B1(new_n793), .B2(G190), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n792), .B1(G294), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(G20), .A2(G179), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT99), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G200), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n280), .B1(new_n802), .B2(G303), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT103), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n800), .A2(G322), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n798), .A2(new_n363), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n799), .A2(new_n310), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G311), .A2(new_n807), .B1(new_n808), .B2(G326), .ZN(new_n809));
  INV_X1    g0609(.A(new_n803), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n806), .A2(new_n310), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT33), .B(G317), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n810), .A2(KEYINPUT103), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n796), .A2(new_n805), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n787), .A2(G159), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT32), .Z(new_n816));
  INV_X1    g0616(.A(new_n791), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G107), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n802), .A2(G87), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(new_n819), .A3(new_n280), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G68), .B2(new_n811), .ZN(new_n821));
  INV_X1    g0621(.A(new_n808), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n816), .B(new_n821), .C1(new_n242), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n800), .ZN(new_n824));
  INV_X1    g0624(.A(new_n807), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n318), .A2(new_n824), .B1(new_n825), .B2(new_n279), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n826), .A2(KEYINPUT100), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n794), .B(KEYINPUT102), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G97), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n826), .A2(KEYINPUT100), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n814), .B1(new_n823), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n782), .B1(new_n832), .B2(new_n779), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n687), .A2(new_n688), .ZN(new_n834));
  INV_X1    g0634(.A(new_n778), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n689), .ZN(new_n837));
  INV_X1    g0637(.A(new_n766), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n834), .A2(G330), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(G396));
  NAND2_X1  g0641(.A1(new_n671), .A2(new_n681), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n394), .A2(new_n680), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n397), .B1(new_n395), .B2(new_n681), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(new_n394), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n681), .B(new_n845), .C1(new_n657), .C2(new_n670), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n759), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n766), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n759), .A2(new_n847), .A3(new_n848), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n779), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n777), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n766), .B1(G77), .B2(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G143), .A2(new_n800), .B1(new_n807), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  INV_X1    g0657(.A(new_n811), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n856), .B1(new_n857), .B2(new_n822), .C1(new_n301), .C2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT34), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n280), .B1(new_n801), .B2(new_n242), .C1(new_n218), .C2(new_n791), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G132), .B2(new_n787), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(new_n318), .C2(new_n794), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n859), .A2(new_n860), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G283), .A2(new_n811), .B1(new_n808), .B2(G303), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n506), .B2(new_n825), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT104), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n787), .A2(G311), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n817), .A2(G87), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n280), .B1(new_n802), .B2(G107), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(G294), .B2(new_n800), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n870), .A2(new_n829), .A3(new_n875), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n864), .A2(new_n865), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n855), .B1(new_n877), .B2(new_n779), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n845), .B2(new_n777), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n852), .A2(new_n879), .ZN(G384));
  NOR2_X1   g0680(.A1(new_n763), .A2(new_n205), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n750), .A2(new_n680), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(new_n755), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n733), .A2(new_n734), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n733), .A2(new_n734), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n435), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT106), .Z(new_n890));
  NOR2_X1   g0690(.A1(new_n430), .A2(new_n681), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n429), .B2(new_n432), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n429), .A2(new_n432), .A3(new_n892), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n846), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n323), .B1(new_n328), .B2(new_n329), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n331), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n353), .B1(new_n360), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(new_n678), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n372), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n365), .A2(new_n334), .A3(new_n336), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n899), .B2(new_n678), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n348), .A2(new_n349), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n678), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n337), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n351), .A2(new_n908), .A3(new_n909), .A4(new_n902), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n901), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n901), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT40), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n888), .A2(new_n896), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n884), .B1(new_n732), .B2(new_n735), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n901), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n919));
  XOR2_X1   g0719(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n908), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n372), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n351), .A2(new_n908), .A3(new_n902), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n910), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n921), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n429), .A2(new_n432), .A3(new_n892), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n845), .B1(new_n929), .B2(new_n893), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n918), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n917), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n674), .B1(new_n890), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n890), .B2(new_n933), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n640), .B1(new_n731), .B2(new_n435), .ZN(new_n936));
  INV_X1    g0736(.A(new_n843), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n848), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n914), .A2(new_n915), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n894), .A2(new_n895), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n919), .B2(new_n927), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n429), .A2(new_n680), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n352), .ZN(new_n948));
  INV_X1    g0748(.A(new_n371), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n678), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n941), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n936), .B(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n881), .B1(new_n935), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n952), .B2(new_n935), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n553), .A2(KEYINPUT35), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n553), .A2(KEYINPUT35), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n955), .A2(G116), .A3(new_n215), .A4(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT36), .ZN(new_n958));
  OAI21_X1  g0758(.A(G77), .B1(new_n318), .B2(new_n218), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n243), .B1(new_n212), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(G1), .A3(new_n290), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n958), .A3(new_n961), .ZN(G367));
  NAND2_X1  g0762(.A1(new_n231), .A2(new_n771), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(new_n780), .C1(new_n209), .C2(new_n383), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n964), .A2(KEYINPUT108), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(KEYINPUT108), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n965), .A2(new_n966), .A3(new_n838), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n630), .A2(new_n681), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n707), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n968), .A2(new_n625), .A3(new_n618), .A4(new_n647), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G294), .A2(new_n811), .B1(new_n808), .B2(G311), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n789), .B2(new_n825), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n802), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n974), .B(new_n344), .C1(new_n561), .C2(new_n791), .ZN(new_n975));
  INV_X1    g0775(.A(new_n787), .ZN(new_n976));
  INV_X1    g0776(.A(G317), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n801), .A2(new_n506), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n976), .A2(new_n977), .B1(KEYINPUT46), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(G303), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n824), .A2(new_n980), .B1(new_n794), .B2(new_n376), .ZN(new_n981));
  NOR4_X1   g0781(.A1(new_n973), .A2(new_n975), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT109), .Z(new_n983));
  NOR2_X1   g0783(.A1(new_n824), .A2(new_n301), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n344), .B1(new_n802), .B2(G58), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n279), .B2(new_n791), .C1(new_n976), .C2(new_n857), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n984), .B(new_n986), .C1(G143), .C2(new_n808), .ZN(new_n987));
  INV_X1    g0787(.A(G159), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n242), .A2(new_n825), .B1(new_n858), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n828), .A2(G68), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n987), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n983), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT111), .Z(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n967), .B1(new_n835), .B2(new_n971), .C1(new_n996), .C2(new_n853), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n722), .A2(new_n723), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n582), .A2(new_n681), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n577), .B2(new_n681), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n698), .A2(new_n1002), .A3(new_n695), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n698), .A2(new_n1002), .A3(KEYINPUT45), .A4(new_n695), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1002), .B1(new_n698), .B2(new_n695), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1008), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1002), .C1(new_n695), .C2(new_n698), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1007), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n694), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n694), .B(new_n1007), .C1(new_n1013), .C2(new_n1012), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n698), .B1(new_n693), .B2(new_n697), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n689), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n760), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n760), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n700), .B(KEYINPUT41), .Z(new_n1023));
  AOI21_X1  g0823(.A(new_n765), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1002), .A2(new_n502), .A3(new_n697), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT42), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n577), .B1(new_n1001), .B2(new_n717), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1025), .A2(KEYINPUT42), .B1(new_n681), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n971), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT43), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1026), .A2(new_n1028), .A3(new_n1031), .A4(new_n1030), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1015), .A2(new_n1002), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1036), .B(new_n1037), .Z(new_n1038));
  OAI21_X1  g0838(.A(new_n997), .B1(new_n1024), .B2(new_n1038), .ZN(G387));
  NAND3_X1  g0839(.A1(new_n691), .A2(new_n692), .A3(new_n778), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n767), .A2(new_n701), .B1(G107), .B2(new_n209), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n235), .A2(G45), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n701), .ZN(new_n1043));
  AOI211_X1 g0843(.A(G45), .B(new_n1043), .C1(G68), .C2(G77), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n299), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n772), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1041), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n766), .B1(new_n1048), .B2(new_n781), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n299), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G68), .A2(new_n807), .B1(new_n811), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT113), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n828), .A2(new_n612), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n824), .A2(new_n242), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n976), .A2(new_n301), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n280), .B1(new_n801), .B2(new_n279), .C1(new_n561), .C2(new_n791), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n808), .A2(G159), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT112), .Z(new_n1059));
  NAND4_X1  g0859(.A1(new_n1052), .A2(new_n1053), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(G294), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n794), .A2(new_n789), .B1(new_n1061), .B2(new_n801), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G311), .A2(new_n811), .B1(new_n808), .B2(G322), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n980), .B2(new_n825), .C1(new_n977), .C2(new_n824), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT48), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT49), .Z(new_n1068));
  NAND2_X1  g0868(.A1(new_n787), .A2(G326), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n344), .C1(new_n506), .C2(new_n791), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1060), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1049), .B1(new_n1071), .B2(new_n779), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1020), .A2(new_n765), .B1(new_n1040), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1021), .A2(new_n762), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n760), .A2(new_n1020), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(G393));
  NAND3_X1  g0876(.A1(new_n1016), .A2(new_n765), .A3(new_n1017), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n240), .A2(new_n772), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n780), .B1(new_n561), .B2(new_n209), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n766), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G50), .A2(new_n811), .B1(new_n807), .B2(new_n1050), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT114), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n828), .A2(G77), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n872), .B(new_n280), .C1(new_n218), .C2(new_n801), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G143), .B2(new_n787), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G150), .A2(new_n808), .B1(new_n800), .B2(G159), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G311), .A2(new_n800), .B1(new_n808), .B2(G317), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n795), .A2(new_n507), .B1(G294), .B2(new_n807), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n818), .B(new_n344), .C1(new_n789), .C2(new_n801), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G322), .B2(new_n787), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(new_n980), .C2(new_n858), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1086), .A2(new_n1088), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1080), .B1(new_n1095), .B2(new_n779), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT115), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n835), .B2(new_n1002), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1077), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n762), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(G390));
  NOR2_X1   g0903(.A1(new_n929), .A2(new_n893), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n937), .B2(new_n848), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n943), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n944), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1105), .A2(new_n946), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n726), .A2(new_n727), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n714), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n729), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n844), .A2(new_n394), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n681), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1104), .B1(new_n1113), .B2(new_n937), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n928), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n945), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1108), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n918), .A2(new_n930), .A3(KEYINPUT116), .A4(new_n674), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n888), .A2(KEYINPUT116), .A3(G330), .A4(new_n896), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1120), .A2(new_n759), .A3(new_n845), .A4(new_n940), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n1108), .C1(new_n1114), .C2(new_n1116), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1119), .A2(new_n765), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n776), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n766), .B1(new_n1050), .B2(new_n854), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT117), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n280), .B1(new_n791), .B2(new_n242), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n801), .A2(new_n301), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1127), .B(new_n1130), .C1(G125), .C2(new_n787), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n828), .A2(G159), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT54), .B(G143), .Z(new_n1133));
  AOI22_X1  g0933(.A1(G137), .A2(new_n811), .B1(new_n807), .B2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G128), .A2(new_n808), .B1(new_n800), .B2(G132), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT119), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n376), .A2(new_n858), .B1(new_n824), .B2(new_n505), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G283), .B2(new_n808), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n976), .A2(new_n1061), .B1(new_n218), .B2(new_n791), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT120), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n344), .B(new_n819), .C1(new_n825), .C2(new_n561), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1143), .B2(new_n1142), .ZN(new_n1146));
  AND4_X1   g0946(.A1(new_n1083), .A2(new_n1141), .A3(new_n1144), .A4(new_n1146), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1138), .A2(new_n1139), .A3(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1124), .B(new_n1126), .C1(new_n853), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1123), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n940), .B1(new_n759), .B2(new_n845), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n918), .A2(new_n674), .A3(new_n930), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n938), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n843), .B1(new_n730), .B2(new_n1112), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n736), .A2(new_n758), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1156), .A2(G330), .A3(new_n845), .A4(new_n940), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n918), .A2(new_n674), .A3(new_n846), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1155), .B(new_n1157), .C1(new_n1158), .C2(new_n940), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n705), .B1(new_n1111), .B2(new_n681), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n706), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n435), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n435), .A2(G330), .A3(new_n888), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n641), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n700), .B1(new_n1151), .B2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1119), .A2(new_n1122), .A3(new_n1160), .A4(new_n1166), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1150), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(G378));
  NAND2_X1  g0971(.A1(new_n312), .A2(new_n316), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n315), .A2(new_n907), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT121), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n317), .A2(new_n1173), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT121), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n1180), .A3(new_n1175), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1178), .A2(new_n1183), .A3(new_n1181), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n888), .A2(new_n1115), .A3(new_n896), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n930), .B1(new_n736), .B2(new_n885), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1188), .A2(KEYINPUT40), .B1(new_n1189), .B2(new_n916), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1190), .A2(new_n951), .A3(new_n674), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n941), .A2(new_n947), .A3(new_n950), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n933), .B2(G330), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1187), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n951), .B1(new_n1190), .B2(new_n674), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n933), .A2(G330), .A3(new_n1192), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n1186), .A4(new_n1185), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n765), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n766), .B1(G50), .B2(new_n854), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n344), .A2(new_n479), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G77), .B2(new_n802), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n318), .B2(new_n791), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G283), .B2(new_n787), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G107), .A2(new_n800), .B1(new_n807), .B2(new_n612), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G97), .A2(new_n811), .B1(new_n808), .B2(G116), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n991), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT58), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G50), .B1(new_n274), .B2(new_n249), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1207), .A2(new_n1208), .B1(new_n1201), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n828), .A2(G150), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n800), .A2(G128), .B1(new_n802), .B2(new_n1133), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n807), .A2(G137), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G125), .A2(new_n808), .B1(new_n811), .B2(G132), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n274), .B(new_n249), .C1(new_n791), .C2(new_n988), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n787), .B2(G124), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1210), .B1(new_n1208), .B2(new_n1207), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1200), .B1(new_n1221), .B2(new_n779), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1187), .B2(new_n777), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1199), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT122), .B1(new_n936), .B2(new_n1164), .ZN(new_n1225));
  AND4_X1   g1025(.A1(KEYINPUT122), .A2(new_n1163), .A3(new_n641), .A4(new_n1164), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1169), .A2(new_n1227), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n762), .B1(new_n1228), .B2(KEYINPUT57), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1169), .A2(new_n1227), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1230), .A2(KEYINPUT57), .A3(new_n1198), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1224), .B1(new_n1229), .B2(new_n1231), .ZN(G375));
  NAND3_X1  g1032(.A1(new_n1165), .A2(new_n1154), .A3(new_n1159), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT123), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT123), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1165), .A2(new_n1154), .A3(new_n1159), .A4(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1234), .A2(new_n1023), .A3(new_n1167), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1104), .A2(new_n776), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n766), .B1(G68), .B2(new_n854), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n828), .A2(G50), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n280), .B1(new_n801), .B2(new_n988), .C1(new_n318), .C2(new_n791), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G128), .B2(new_n787), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G137), .A2(new_n800), .B1(new_n811), .B2(new_n1133), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G132), .A2(new_n808), .B1(new_n807), .B2(G150), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1240), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1053), .B1(new_n789), .B2(new_n824), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT125), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G294), .A2(new_n808), .B1(new_n811), .B2(new_n507), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n807), .A2(G107), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n787), .A2(G303), .B1(G97), .B2(new_n802), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n344), .B1(new_n791), .B2(new_n279), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT124), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1245), .B1(new_n1247), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1239), .B1(new_n1254), .B2(new_n779), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1160), .A2(new_n765), .B1(new_n1238), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1237), .A2(new_n1256), .ZN(G381));
  OR4_X1    g1057(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1258), .A2(G387), .A3(G378), .A4(G381), .ZN(new_n1259));
  INV_X1    g1059(.A(G375), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(G407));
  NAND2_X1  g1061(.A1(new_n679), .A2(G213), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1170), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(G213), .A3(new_n1264), .ZN(G409));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  INV_X1    g1066(.A(G390), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G390), .B(new_n997), .C1(new_n1024), .C2(new_n1038), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(G393), .B(G396), .ZN(new_n1270));
  AND4_X1   g1070(.A1(new_n1266), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(KEYINPUT126), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1272), .A2(new_n1270), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1224), .C1(new_n1229), .C2(new_n1231), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1228), .A2(new_n1023), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1199), .A2(new_n1223), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1170), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1165), .A2(new_n1154), .A3(new_n1159), .A4(KEYINPUT60), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1280), .A2(new_n762), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT60), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1281), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1285), .A2(G384), .A3(new_n1256), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G384), .B1(new_n1285), .B2(new_n1256), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1279), .A2(new_n1288), .A3(new_n1262), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1274), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1263), .A2(G2897), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1285), .A2(new_n1256), .ZN(new_n1295));
  INV_X1    g1095(.A(G384), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1285), .A2(G384), .A3(new_n1256), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1292), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1279), .A2(new_n1262), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT61), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1263), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1288), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1291), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1306), .B1(new_n1307), .B2(new_n1303), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1289), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1303), .A2(KEYINPUT62), .A3(new_n1288), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1274), .B(KEYINPUT127), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1305), .B1(new_n1312), .B2(new_n1313), .ZN(G405));
  NAND2_X1  g1114(.A1(G375), .A2(new_n1170), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1275), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1288), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1315), .B(new_n1275), .C1(new_n1287), .C2(new_n1286), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(new_n1274), .ZN(G402));
endmodule


