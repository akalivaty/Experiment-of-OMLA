//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n459), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n459), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OR3_X1    g044(.A1(new_n463), .A2(KEYINPUT67), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT67), .B1(new_n463), .B2(new_n469), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n464), .A2(new_n465), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT68), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n478), .B1(new_n474), .B2(new_n459), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n460), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n477), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(KEYINPUT70), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n459), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(new_n487), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n460), .A2(G126), .A3(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT71), .A2(G138), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n459), .B(new_n497), .C1(new_n464), .C2(new_n465), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n459), .A4(new_n497), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n495), .A2(new_n496), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT72), .A3(G651), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n506), .A2(new_n508), .B1(KEYINPUT6), .B2(new_n505), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT73), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(G651), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n509), .A2(G88), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n510), .A2(new_n519), .A3(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  AND2_X1   g098(.A1(new_n509), .A2(new_n520), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT74), .B(G89), .Z(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n506), .A2(new_n508), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n527), .A2(G543), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n520), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n526), .A2(new_n530), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n524), .A2(G90), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n505), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n529), .A2(G52), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND4_X1  g118(.A1(new_n527), .A2(G43), .A3(G543), .A4(new_n528), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n527), .A2(G81), .A3(new_n528), .A4(new_n520), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AND2_X1   g122(.A1(KEYINPUT5), .A2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(KEYINPUT5), .A2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n505), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g129(.A(KEYINPUT75), .B(new_n547), .C1(new_n550), .C2(new_n551), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n546), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n527), .A2(G543), .A3(new_n528), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n509), .A2(new_n565), .A3(G53), .A4(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n509), .A2(G91), .A3(new_n520), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n516), .B2(new_n517), .ZN(new_n570));
  AND2_X1   g145(.A1(G78), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n567), .A2(new_n573), .ZN(G299));
  NAND3_X1  g149(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n509), .A2(G87), .A3(new_n520), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n516), .B2(new_n517), .ZN(new_n580));
  AND2_X1   g155(.A1(G73), .A2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n527), .A2(G48), .A3(G543), .A4(new_n528), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n527), .A2(G86), .A3(new_n528), .A4(new_n520), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G305));
  NAND3_X1  g160(.A1(new_n509), .A2(G85), .A3(new_n520), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n527), .A2(G47), .A3(G543), .A4(new_n528), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n516), .B2(new_n517), .ZN(new_n589));
  AND2_X1   g164(.A1(G72), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n586), .A2(new_n591), .A3(KEYINPUT76), .A4(new_n587), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n527), .A2(G92), .A3(new_n528), .A4(new_n520), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n509), .A2(KEYINPUT10), .A3(G92), .A4(new_n520), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(G66), .B1(new_n548), .B2(new_n549), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n505), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n529), .B2(G54), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(new_n611), .B2(G168), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n554), .A2(new_n555), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n617), .A2(new_n544), .A3(new_n545), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n611), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n607), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n611), .ZN(G323));
  XOR2_X1   g196(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n622));
  XNOR2_X1  g197(.A(G323), .B(new_n622), .ZN(G282));
  NOR2_X1   g198(.A1(new_n474), .A2(new_n468), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT13), .Z(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT78), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n475), .A2(G135), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  AOI211_X1 g210(.A(new_n632), .B(new_n635), .C1(new_n481), .C2(G123), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n627), .A2(G2100), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n629), .B(new_n637), .C1(new_n630), .C2(new_n636), .ZN(G156));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT79), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n644), .B2(new_n645), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  AND2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n652), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n648), .A2(new_n649), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n648), .A2(new_n649), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n641), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n652), .B1(new_n650), .B2(new_n651), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n654), .A3(new_n656), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n660), .A3(new_n640), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(G14), .A3(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n668));
  AOI21_X1  g243(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT81), .ZN(new_n670));
  INV_X1    g245(.A(new_n668), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n665), .A2(new_n666), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n681), .A2(new_n688), .A3(new_n684), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n681), .A2(new_n688), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT20), .Z(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n694), .B1(new_n690), .B2(new_n692), .ZN(new_n698));
  AND3_X1   g273(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n697), .B1(new_n695), .B2(new_n698), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n679), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(new_n698), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(new_n696), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n703), .A2(new_n678), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G26), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n481), .A2(G128), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n712));
  INV_X1    g287(.A(G116), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(G2105), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n475), .B2(G140), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n710), .B1(new_n716), .B2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G2067), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G5), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G171), .B2(new_n720), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n719), .B1(G1961), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G34), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(new_n708), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n472), .B2(new_n708), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2084), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT84), .B(G16), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G19), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n556), .B2(new_n729), .ZN(new_n731));
  INV_X1    g306(.A(G1341), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n722), .A2(G1961), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n708), .A2(G27), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G164), .B2(new_n708), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2078), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n723), .A2(new_n728), .A3(new_n733), .A4(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n708), .A2(G32), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT26), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n741), .B(new_n743), .C1(G141), .C2(new_n475), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n481), .A2(G129), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(G29), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT27), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G1996), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n747), .A2(new_n748), .ZN(new_n752));
  OR3_X1    g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n608), .A2(new_n720), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G4), .B2(new_n720), .ZN(new_n755));
  INV_X1    g330(.A(G1348), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n755), .A2(new_n756), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n753), .A2(new_n757), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n720), .A2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G168), .B2(new_n720), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT95), .B(KEYINPUT23), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT96), .ZN(new_n766));
  INV_X1    g341(.A(new_n729), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G20), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G16), .B2(G299), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n636), .A2(G29), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT30), .B(G28), .ZN(new_n774));
  OR2_X1    g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n774), .A2(new_n708), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND3_X1   g352(.A1(new_n772), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n773), .B1(new_n772), .B2(new_n777), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n764), .B(new_n771), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n739), .A2(new_n760), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n460), .A2(G127), .ZN(new_n782));
  AND2_X1   g357(.A1(G115), .A2(G2104), .ZN(new_n783));
  OAI21_X1  g358(.A(G2105), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT25), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n475), .A2(G139), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT89), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT89), .B1(new_n786), .B2(new_n787), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT90), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT90), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(new_n784), .C1(new_n788), .C2(new_n789), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n791), .A2(G29), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G29), .A2(G33), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT88), .Z(new_n796));
  AND2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(G2072), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n485), .A2(G29), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT29), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n708), .A2(G35), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT93), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n800), .B1(new_n799), .B2(new_n802), .ZN(new_n804));
  OAI21_X1  g379(.A(G2090), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n797), .A2(G2072), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n798), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n803), .A2(new_n804), .ZN(new_n808));
  INV_X1    g383(.A(G2090), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT94), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(KEYINPUT94), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n767), .B1(G290), .B2(KEYINPUT85), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(KEYINPUT85), .B2(G290), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n767), .A2(G24), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(G1986), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n708), .A2(G25), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n481), .A2(G119), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n821));
  INV_X1    g396(.A(G107), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(G2105), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n475), .B2(G131), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n819), .B1(new_n825), .B2(G29), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT35), .B(G1991), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT83), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n826), .A2(new_n829), .ZN(new_n831));
  AOI211_X1 g406(.A(new_n830), .B(new_n831), .C1(KEYINPUT87), .C2(KEYINPUT36), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n817), .A2(G1986), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n818), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(G16), .A2(G23), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT86), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G288), .B2(new_n720), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT33), .ZN(new_n838));
  INV_X1    g413(.A(G1976), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n729), .A2(G22), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G166), .B2(new_n729), .ZN(new_n842));
  INV_X1    g417(.A(G1971), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(G6), .A2(G16), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(G16), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT32), .B(G1981), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n840), .A2(KEYINPUT34), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT34), .B1(new_n840), .B2(new_n851), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n834), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n781), .B(new_n813), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT97), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n813), .A2(new_n781), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n854), .A2(new_n855), .ZN(new_n861));
  OAI221_X1 g436(.A(new_n834), .B1(KEYINPUT87), .B2(KEYINPUT36), .C1(new_n852), .C2(new_n853), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n858), .A2(new_n863), .ZN(G311));
  NAND3_X1  g439(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(G150));
  NAND4_X1  g440(.A1(new_n527), .A2(G55), .A3(G543), .A4(new_n528), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n527), .A2(G93), .A3(new_n528), .A4(new_n520), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n869));
  INV_X1    g444(.A(G67), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n516), .B2(new_n517), .ZN(new_n871));
  NAND2_X1  g446(.A1(G80), .A2(G543), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g449(.A(KEYINPUT99), .B(new_n872), .C1(new_n550), .C2(new_n870), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(G651), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n868), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT100), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n868), .A2(new_n880), .A3(new_n876), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n878), .A2(new_n618), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n868), .A2(new_n880), .A3(new_n876), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n880), .B1(new_n868), .B2(new_n876), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n883), .A2(new_n884), .A3(new_n556), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n556), .A2(new_n877), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT101), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n882), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n607), .A2(new_n615), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n891));
  XOR2_X1   g466(.A(new_n890), .B(new_n891), .Z(new_n892));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n893));
  AOI21_X1  g468(.A(G860), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n878), .A2(new_n881), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(G860), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT102), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n899), .ZN(G145));
  NAND2_X1  g475(.A1(new_n481), .A2(G130), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n475), .A2(G142), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n459), .A2(G118), .ZN(new_n903));
  OAI21_X1  g478(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n625), .ZN(new_n906));
  INV_X1    g481(.A(new_n825), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n711), .A2(new_n715), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n746), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n716), .A2(new_n745), .A3(new_n744), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n502), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n502), .B1(new_n911), .B2(new_n912), .ZN(new_n915));
  OAI211_X1 g490(.A(KEYINPUT103), .B(new_n790), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n915), .ZN(new_n917));
  INV_X1    g492(.A(new_n793), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n790), .A2(KEYINPUT90), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(KEYINPUT103), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n920), .A3(new_n913), .ZN(new_n921));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n916), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n916), .B2(new_n921), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n909), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n917), .A2(new_n920), .A3(new_n913), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n790), .A2(KEYINPUT103), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n917), .B2(new_n913), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n916), .A2(new_n921), .A3(new_n923), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n908), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G160), .B(new_n485), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(new_n636), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n926), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G37), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n926), .B2(new_n932), .ZN(new_n938));
  XOR2_X1   g513(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n939));
  OR3_X1    g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(new_n937), .B2(new_n938), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(G395));
  OR2_X1    g517(.A1(new_n888), .A2(new_n620), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n888), .A2(new_n620), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n567), .A2(new_n602), .A3(new_n573), .A4(new_n606), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n567), .A2(new_n573), .B1(new_n602), .B2(new_n606), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(G299), .A2(new_n607), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n948), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n951), .B1(new_n953), .B2(KEYINPUT41), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n945), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n953), .B(KEYINPUT107), .Z(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n943), .A3(new_n944), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n594), .B2(new_n595), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n594), .A2(new_n960), .A3(new_n595), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g539(.A1(G303), .A2(KEYINPUT109), .ZN(new_n965));
  NAND2_X1  g540(.A1(G303), .A2(KEYINPUT109), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n846), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n966), .A3(G305), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n964), .A2(KEYINPUT110), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n962), .A2(KEYINPUT110), .A3(new_n963), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  INV_X1    g548(.A(new_n963), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n961), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n970), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n955), .A2(new_n978), .A3(new_n957), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n959), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n959), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g556(.A(G868), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n896), .A2(new_n611), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(G295));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n983), .ZN(G331));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n986));
  XNOR2_X1  g561(.A(G286), .B(G301), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n888), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n879), .B1(new_n556), .B2(new_n877), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n896), .B2(new_n556), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n987), .A3(new_n882), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n954), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n989), .A2(new_n992), .A3(new_n954), .A4(KEYINPUT112), .ZN(new_n996));
  INV_X1    g571(.A(new_n953), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n888), .A2(new_n988), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n987), .B1(new_n991), .B2(new_n882), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n995), .A2(new_n977), .A3(new_n996), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n936), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n989), .A2(new_n992), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n993), .A2(new_n994), .B1(new_n1003), .B2(new_n997), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n977), .B1(new_n1004), .B2(new_n996), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n986), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n952), .A2(new_n948), .A3(new_n946), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1009), .A2(KEYINPUT113), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT41), .B1(new_n949), .B2(new_n950), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(KEYINPUT113), .A3(new_n1009), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n989), .A2(new_n992), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1013), .A2(KEYINPUT114), .B1(new_n1003), .B2(new_n956), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1012), .A2(new_n1010), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n989), .A4(new_n992), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n977), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT43), .B1(new_n1002), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT115), .B(KEYINPUT43), .C1(new_n1002), .C2(new_n1018), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1008), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1024));
  INV_X1    g599(.A(new_n977), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1026), .A2(new_n1007), .A3(new_n936), .A4(new_n1001), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT43), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1023), .A2(new_n1031), .ZN(G397));
  INV_X1    g607(.A(KEYINPUT127), .ZN(new_n1033));
  INV_X1    g608(.A(G1384), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n502), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n461), .A2(new_n462), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G2105), .ZN(new_n1039));
  INV_X1    g614(.A(new_n469), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1039), .A2(G40), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n1034), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n763), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1040), .A3(G40), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n1035), .B2(KEYINPUT50), .ZN(new_n1046));
  INV_X1    g621(.A(G2084), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n502), .A2(new_n1048), .A3(new_n1034), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1044), .A2(G168), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(G168), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT51), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1056), .A3(G8), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT117), .B(G1981), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n846), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G305), .A2(G1981), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n502), .A2(new_n1034), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n1041), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1060), .A2(new_n1061), .A3(KEYINPUT49), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n960), .A2(new_n1070), .A3(G1976), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT116), .B1(G288), .B2(new_n839), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n463), .A2(new_n469), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1073), .A2(new_n502), .A3(G40), .A4(new_n1034), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .A4(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT52), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n839), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1067), .A2(new_n1072), .A3(new_n1071), .A4(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1069), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G303), .A2(G8), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(KEYINPUT55), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1043), .A2(new_n843), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1046), .A2(new_n809), .A3(new_n1049), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1065), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1079), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1045), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1090));
  INV_X1    g665(.A(G2078), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(KEYINPUT53), .A3(new_n1091), .A4(new_n1042), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1043), .B2(G2078), .ZN(new_n1095));
  AOI21_X1  g670(.A(G301), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G8), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(KEYINPUT120), .A3(new_n1081), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1085), .B2(new_n1082), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1086), .A2(new_n1096), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1033), .B1(new_n1058), .B2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1086), .A2(new_n1101), .A3(new_n1099), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(KEYINPUT127), .A4(new_n1096), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1057), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1053), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(G8), .A3(new_n1051), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1109), .B2(KEYINPUT51), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(new_n1055), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1103), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(new_n732), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1074), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1074), .A2(KEYINPUT124), .A3(new_n1114), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1043), .A2(G1996), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n556), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT59), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1123), .B(new_n556), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1090), .A2(new_n1042), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1035), .A2(KEYINPUT50), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1128), .A2(new_n1041), .A3(new_n1049), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1127), .B1(new_n1129), .B2(G1956), .ZN(new_n1130));
  XNOR2_X1  g705(.A(G299), .B(KEYINPUT57), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1125), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(G1956), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n1135));
  XNOR2_X1  g710(.A(G299), .B(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1136), .A3(new_n1127), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1122), .A2(new_n1124), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1134), .B2(new_n1127), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT61), .B1(new_n1139), .B2(KEYINPUT125), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(new_n1137), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT122), .B1(new_n1074), .B2(G2067), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1066), .A2(new_n1041), .A3(new_n1146), .A4(new_n718), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(G1348), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n1150));
  NOR4_X1   g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n608), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n607), .B1(new_n1152), .B2(KEYINPUT60), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1150), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1151), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1138), .A2(new_n1144), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1152), .A2(new_n607), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1139), .B1(new_n1157), .B2(new_n1137), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1086), .A2(new_n1101), .A3(new_n1099), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1095), .A2(new_n1089), .A3(G301), .A4(new_n1092), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT54), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1096), .A2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1110), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1166), .B(new_n1167), .C1(new_n1096), .C2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1159), .A2(new_n1164), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1172));
  NOR2_X1   g747(.A1(G286), .A2(new_n1065), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1172), .A2(KEYINPUT121), .A3(new_n1173), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1171), .B1(new_n1160), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1171), .B1(new_n1098), .B2(new_n1081), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1178), .A2(new_n1086), .A3(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(G288), .A2(G1976), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT118), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1060), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1067), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1085), .A2(new_n1082), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1187), .B1(new_n1188), .B2(new_n1079), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT119), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1187), .B(KEYINPUT119), .C1(new_n1188), .C2(new_n1079), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1180), .A2(new_n1182), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1112), .A2(new_n1170), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1037), .A2(new_n1045), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n910), .A2(new_n718), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n716), .A2(G2067), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n746), .B(new_n751), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n825), .A2(new_n828), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n907), .A2(new_n829), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(G290), .B(G1986), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1195), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1194), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(G290), .A2(G1986), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1195), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1208), .A2(KEYINPUT48), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1208), .A2(KEYINPUT48), .ZN(new_n1210));
  AOI211_X1 g785(.A(new_n1209), .B(new_n1210), .C1(new_n1195), .C2(new_n1202), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1198), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1195), .B1(new_n1212), .B2(new_n746), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1195), .A2(new_n751), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1214), .B(KEYINPUT46), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n1216), .B(KEYINPUT47), .Z(new_n1217));
  NAND2_X1  g792(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1196), .B1(new_n1218), .B2(new_n1201), .ZN(new_n1219));
  AOI211_X1 g794(.A(new_n1211), .B(new_n1217), .C1(new_n1195), .C2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1205), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g796(.A(G319), .ZN(new_n1223));
  NOR2_X1   g797(.A1(G227), .A2(new_n1223), .ZN(new_n1224));
  AND3_X1   g798(.A1(new_n706), .A2(new_n662), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g799(.A(new_n1225), .B1(new_n937), .B2(new_n938), .ZN(new_n1226));
  AOI21_X1  g800(.A(new_n1226), .B1(new_n1028), .B2(new_n1027), .ZN(G308));
  OAI211_X1 g801(.A(new_n1029), .B(new_n1225), .C1(new_n938), .C2(new_n937), .ZN(G225));
endmodule


