//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT66), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G116), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G119), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n194), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(new_n196), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n200), .A2(new_n194), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G104), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G101), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n204), .A2(new_n207), .A3(new_n211), .A4(new_n208), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n214), .A3(G101), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n202), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n203), .A2(G107), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n206), .A2(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(G101), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT5), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(new_n193), .B2(new_n198), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT83), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n195), .B2(KEYINPUT5), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n221), .A2(new_n191), .A3(KEYINPUT83), .A4(G116), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(G113), .A3(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n220), .B(new_n201), .C1(new_n222), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n216), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G110), .B(G122), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n216), .A2(new_n227), .A3(new_n229), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(KEYINPUT6), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G146), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n235), .A2(G146), .ZN(new_n238));
  INV_X1    g052(.A(G146), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G143), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n237), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n235), .A2(G146), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(G128), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n236), .B(new_n241), .C1(new_n234), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G125), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n248), .B(new_n249), .C1(new_n238), .C2(new_n240), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n242), .A2(new_n243), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(G125), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G224), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n256), .B(KEYINPUT84), .Z(new_n257));
  XNOR2_X1  g071(.A(new_n254), .B(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n228), .A2(new_n259), .A3(new_n230), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n233), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n233), .A2(new_n258), .A3(KEYINPUT85), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G902), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n200), .A2(new_n194), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n197), .B1(new_n195), .B2(new_n196), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT5), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n224), .A2(G113), .A3(new_n225), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n220), .A2(new_n201), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n200), .A2(new_n221), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n226), .A2(new_n274), .ZN(new_n275));
  OAI22_X1  g089(.A1(new_n272), .A2(new_n220), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n229), .B(KEYINPUT8), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n256), .A2(KEYINPUT7), .ZN(new_n279));
  AOI21_X1  g093(.A(G128), .B1(new_n242), .B2(new_n243), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n242), .A2(new_n243), .A3(G128), .ZN(new_n281));
  INV_X1    g095(.A(new_n234), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(G125), .B1(new_n283), .B2(new_n236), .ZN(new_n284));
  INV_X1    g098(.A(new_n253), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n279), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n279), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n247), .A2(new_n253), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT86), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n278), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n232), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n290), .B1(new_n278), .B2(new_n289), .ZN(new_n293));
  OAI211_X1 g107(.A(KEYINPUT87), .B(new_n266), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n265), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n293), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n232), .A3(new_n291), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT87), .B1(new_n297), .B2(new_n266), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n188), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n266), .B1(new_n292), .B2(new_n293), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n303), .A2(new_n187), .A3(new_n265), .A4(new_n294), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n304), .A2(new_n300), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n308), .B(KEYINPUT82), .Z(new_n309));
  NOR2_X1   g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G217), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(G234), .B2(new_n266), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G953), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(G221), .A2(G234), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT73), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT68), .B(G953), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G221), .A4(G234), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G137), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n320), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n324), .B1(new_n320), .B2(new_n323), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n191), .B2(G128), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n237), .A2(KEYINPUT23), .A3(G119), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n329), .B(new_n330), .C1(G119), .C2(new_n237), .ZN(new_n331));
  XNOR2_X1  g145(.A(G119), .B(G128), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT24), .B(G110), .Z(new_n333));
  AOI22_X1  g147(.A1(new_n331), .A2(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n246), .A2(KEYINPUT16), .A3(G140), .ZN(new_n335));
  XNOR2_X1  g149(.A(G125), .B(G140), .ZN(new_n336));
  AOI211_X1 g150(.A(new_n239), .B(new_n335), .C1(KEYINPUT16), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(KEYINPUT16), .ZN(new_n338));
  INV_X1    g152(.A(new_n335), .ZN(new_n339));
  AOI21_X1  g153(.A(G146), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n334), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G125), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n246), .A2(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G146), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n335), .B1(new_n336), .B2(KEYINPUT16), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(G146), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n331), .A2(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT74), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n341), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n351), .B1(new_n341), .B2(new_n350), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n327), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT16), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n339), .B1(new_n345), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n239), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n347), .A2(G146), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n360), .A2(new_n334), .B1(new_n348), .B2(new_n349), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n327), .B1(new_n361), .B2(new_n351), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n314), .B1(new_n364), .B2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n341), .A2(new_n350), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT74), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n352), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n362), .B1(new_n368), .B2(new_n327), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT25), .A3(new_n266), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n313), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n312), .A2(G902), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT75), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n355), .A2(new_n363), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT76), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT11), .ZN(new_n379));
  INV_X1    g193(.A(G134), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(G137), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(G137), .ZN(new_n382));
  INV_X1    g196(.A(G137), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT11), .A3(G134), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G131), .ZN(new_n386));
  INV_X1    g200(.A(G131), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(new_n384), .A3(new_n387), .A4(new_n382), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT67), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n249), .A2(new_n248), .ZN(new_n391));
  XNOR2_X1  g205(.A(G143), .B(G146), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n252), .B(new_n390), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n390), .B1(new_n250), .B2(new_n252), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n389), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n382), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n380), .A2(G137), .ZN(new_n398));
  OAI21_X1  g212(.A(G131), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n399), .A2(new_n388), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n245), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n252), .B1(new_n391), .B2(new_n392), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT64), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n250), .A2(KEYINPUT64), .A3(new_n252), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n389), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n407), .A2(new_n401), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n202), .B(new_n402), .C1(new_n408), .C2(KEYINPUT30), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n199), .A2(new_n201), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n396), .A2(new_n410), .A3(new_n401), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G237), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n321), .A2(G210), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT27), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT26), .B(G101), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n407), .A2(new_n401), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n202), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n396), .A2(KEYINPUT28), .A3(new_n410), .A4(new_n401), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT28), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n411), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n423), .A2(new_n424), .A3(new_n417), .A4(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n417), .A3(new_n421), .A4(new_n422), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT69), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT29), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n419), .A2(new_n427), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n426), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n411), .A2(KEYINPUT70), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n396), .A2(new_n434), .A3(new_n410), .A4(new_n401), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n396), .A2(new_n401), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT71), .B1(new_n436), .B2(new_n202), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT71), .ZN(new_n438));
  AOI211_X1 g252(.A(new_n438), .B(new_n410), .C1(new_n396), .C2(new_n401), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n433), .B(new_n435), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n432), .B1(new_n440), .B2(KEYINPUT28), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n418), .A2(new_n430), .ZN(new_n442));
  AOI21_X1  g256(.A(G902), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n431), .B1(new_n443), .B2(KEYINPUT72), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT72), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n445), .B(G902), .C1(new_n441), .C2(new_n442), .ZN(new_n446));
  OAI21_X1  g260(.A(G472), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n409), .A2(new_n417), .A3(new_n411), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT31), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n409), .A2(KEYINPUT31), .A3(new_n417), .A4(new_n411), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n417), .B1(new_n423), .B2(new_n426), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(G472), .A2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT32), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n453), .B1(new_n450), .B2(new_n451), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n458), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n378), .B1(new_n447), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  OAI21_X1  g280(.A(G221), .B1(new_n466), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n321), .A2(G227), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT77), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G140), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n241), .B(new_n475), .C1(new_n234), .C2(new_n244), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n220), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT10), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n213), .B(new_n215), .C1(new_n394), .C2(new_n395), .ZN(new_n480));
  INV_X1    g294(.A(new_n389), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n245), .A2(KEYINPUT10), .A3(new_n220), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT78), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n478), .B1(new_n283), .B2(new_n236), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n220), .A2(new_n486), .B1(new_n477), .B2(new_n478), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n487), .A2(KEYINPUT78), .A3(new_n481), .A4(new_n480), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n245), .A2(new_n220), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n212), .A2(new_n219), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n283), .B2(new_n475), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n389), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n494));
  NOR2_X1   g308(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n493), .B2(new_n495), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n489), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT80), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT80), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n489), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n474), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n473), .B1(new_n485), .B2(new_n488), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n487), .A2(new_n480), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n389), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n469), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n489), .A2(new_n497), .A3(new_n500), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n500), .B1(new_n489), .B2(new_n497), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n473), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(KEYINPUT81), .A3(new_n506), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(G469), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G469), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n503), .A2(new_n497), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n474), .B1(new_n489), .B2(new_n505), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n514), .B(new_n266), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(G469), .A2(G902), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n468), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n315), .A2(new_n317), .A3(G214), .A4(new_n413), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n235), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n321), .A2(G143), .A3(G214), .A4(new_n413), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G131), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT89), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n528), .A3(G131), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(new_n523), .A3(new_n387), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n526), .A2(new_n527), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n360), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n528), .B1(new_n524), .B2(G131), .ZN(new_n533));
  AOI211_X1 g347(.A(KEYINPUT89), .B(new_n387), .C1(new_n522), .C2(new_n523), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT17), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G113), .B(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n203), .ZN(new_n538));
  AND2_X1   g352(.A1(KEYINPUT18), .A2(G131), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n336), .A2(new_n239), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n524), .A2(new_n539), .B1(new_n346), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n524), .A2(new_n539), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n536), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n538), .B1(new_n536), .B2(new_n544), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n266), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G475), .ZN(new_n549));
  NOR2_X1   g363(.A1(G475), .A2(G902), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT91), .ZN(new_n551));
  INV_X1    g365(.A(new_n538), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n336), .A2(KEYINPUT19), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT19), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT90), .B1(new_n555), .B2(G146), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT90), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n557), .B(new_n239), .C1(new_n553), .C2(new_n554), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n359), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n533), .A2(new_n534), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n560), .B2(new_n530), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n552), .B1(new_n561), .B2(new_n543), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n551), .B1(new_n545), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n545), .A2(new_n562), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT92), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT20), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT92), .ZN(new_n568));
  INV_X1    g382(.A(new_n551), .ZN(new_n569));
  AND4_X1   g383(.A1(new_n568), .A2(new_n564), .A3(new_n566), .A4(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n549), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(G234), .A2(G237), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(G952), .A3(new_n255), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT95), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n318), .A2(G902), .A3(new_n572), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT21), .B(G898), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n235), .A2(G128), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n237), .A2(G143), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(new_n380), .ZN(new_n582));
  XNOR2_X1  g396(.A(G116), .B(G122), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n206), .ZN(new_n584));
  INV_X1    g398(.A(G122), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT14), .B1(new_n585), .B2(G116), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT14), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n189), .A3(G122), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(G116), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n586), .A2(new_n588), .A3(KEYINPUT93), .A4(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n590), .B(G107), .C1(KEYINPUT93), .C2(new_n588), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n582), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n579), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n593), .A2(KEYINPUT13), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n580), .B1(new_n593), .B2(KEYINPUT13), .ZN(new_n595));
  OAI21_X1  g409(.A(G134), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n581), .A2(new_n380), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n583), .B(new_n206), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n466), .A2(new_n311), .A3(G953), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n592), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n592), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n266), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n603), .A2(KEYINPUT94), .ZN(new_n604));
  INV_X1    g418(.A(G478), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(KEYINPUT15), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(KEYINPUT94), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n603), .B2(new_n606), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n571), .A2(new_n578), .A3(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n310), .A2(new_n465), .A3(new_n520), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  NAND2_X1  g426(.A1(new_n455), .A2(new_n456), .ZN(new_n613));
  OAI21_X1  g427(.A(G472), .B1(new_n461), .B2(G902), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n377), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n468), .B(new_n615), .C1(new_n513), .C2(new_n519), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n564), .A2(new_n569), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n568), .B1(new_n545), .B2(new_n562), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n617), .B1(KEYINPUT20), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n565), .A2(new_n566), .A3(new_n563), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n619), .A2(new_n620), .B1(G475), .B2(new_n548), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n601), .A2(new_n602), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(KEYINPUT33), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(KEYINPUT33), .ZN(new_n624));
  OAI211_X1 g438(.A(G478), .B(new_n266), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  AOI211_X1 g442(.A(new_n309), .B(new_n578), .C1(new_n299), .C2(new_n304), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n616), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  AOI21_X1  g446(.A(new_n309), .B1(new_n299), .B2(new_n304), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n617), .A2(KEYINPUT20), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n563), .A2(new_n566), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n609), .B(new_n549), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n578), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n633), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n616), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  AND2_X1   g456(.A1(new_n613), .A2(new_n614), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT25), .B1(new_n369), .B2(new_n266), .ZN(new_n644));
  AND4_X1   g458(.A1(KEYINPUT25), .A2(new_n355), .A3(new_n363), .A4(new_n266), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n312), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n366), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n373), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n310), .A2(new_n520), .A3(new_n610), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  INV_X1    g468(.A(new_n650), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n447), .B2(new_n464), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n576), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(KEYINPUT96), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(KEYINPUT96), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n575), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n636), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n656), .A2(new_n520), .A3(new_n633), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XOR2_X1   g478(.A(new_n661), .B(KEYINPUT39), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n520), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n666), .B(KEYINPUT40), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT99), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n307), .A2(KEYINPUT38), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT38), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n305), .B2(new_n306), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n412), .A2(new_n417), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n678), .B(new_n266), .C1(new_n417), .C2(new_n440), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G472), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT97), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n679), .A2(KEYINPUT97), .A3(G472), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n460), .A3(new_n462), .A4(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n309), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n655), .ZN(new_n686));
  INV_X1    g500(.A(new_n609), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n621), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n673), .B1(new_n677), .B2(new_n688), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n677), .A2(new_n673), .A3(new_n688), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n670), .B(new_n672), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  NAND2_X1  g506(.A1(new_n625), .A2(new_n626), .ZN(new_n693));
  INV_X1    g507(.A(new_n661), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n571), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n656), .A2(new_n520), .A3(new_n633), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n489), .A2(new_n505), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n700), .A2(new_n473), .B1(new_n503), .B2(new_n497), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n701), .B2(G902), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n467), .A3(new_n517), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT100), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT100), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n702), .A2(new_n705), .A3(new_n517), .A4(new_n467), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n704), .A2(KEYINPUT101), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT101), .B1(new_n704), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n465), .A2(new_n628), .A3(new_n629), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n699), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n704), .A2(new_n706), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n704), .A2(KEYINPUT101), .A3(new_n706), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n633), .A2(new_n628), .A3(new_n638), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n716), .A2(KEYINPUT102), .A3(new_n465), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n711), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT41), .B(G113), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT103), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(G15));
  OAI211_X1 g537(.A(new_n639), .B(new_n465), .C1(new_n707), .C2(new_n708), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  AND3_X1   g539(.A1(new_n633), .A2(new_n706), .A3(new_n704), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n610), .A3(new_n656), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  OAI21_X1  g542(.A(KEYINPUT104), .B1(new_n621), .B2(new_n687), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n571), .A2(new_n730), .A3(new_n609), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n729), .A2(new_n633), .A3(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n450), .A2(new_n451), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n437), .A2(new_n439), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n433), .A2(new_n435), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT28), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n417), .B1(new_n736), .B2(new_n426), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n456), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n377), .A2(new_n738), .A3(new_n614), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(new_n638), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n732), .B(new_n740), .C1(new_n707), .C2(new_n708), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NAND3_X1  g556(.A1(new_n738), .A2(new_n614), .A3(new_n650), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT105), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n738), .A2(new_n650), .A3(new_n614), .A4(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n695), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n633), .A2(new_n704), .A3(new_n706), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT106), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n726), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  NOR2_X1   g568(.A1(new_n468), .A2(new_n309), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n305), .B2(new_n306), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n518), .B(KEYINPUT107), .Z(new_n758));
  NAND2_X1  g572(.A1(new_n511), .A2(new_n506), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n517), .B(new_n758), .C1(new_n759), .C2(new_n514), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n696), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n455), .A2(new_n762), .A3(new_n459), .ZN(new_n763));
  INV_X1    g577(.A(new_n459), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT108), .B1(new_n461), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n462), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT109), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n763), .A2(new_n462), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n447), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n377), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n773), .A3(new_n377), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n761), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n465), .A2(new_n757), .A3(new_n696), .A4(new_n760), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT42), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n387), .ZN(G33));
  NAND4_X1  g595(.A1(new_n465), .A2(new_n757), .A3(new_n662), .A4(new_n760), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  OR3_X1    g597(.A1(new_n571), .A2(KEYINPUT43), .A3(new_n627), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n621), .A2(new_n693), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT43), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n643), .A2(new_n655), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(KEYINPUT44), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n309), .B1(new_n305), .B2(new_n306), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n787), .A2(new_n788), .ZN(new_n794));
  OAI22_X1  g608(.A1(new_n792), .A2(new_n793), .B1(KEYINPUT44), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n758), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n508), .A2(new_n512), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(G469), .B1(new_n759), .B2(new_n798), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n796), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT111), .B1(new_n802), .B2(KEYINPUT46), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT46), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n800), .B1(new_n797), .B2(new_n798), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n796), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n803), .A2(new_n517), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n467), .A3(new_n665), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n795), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(new_n383), .ZN(G39));
  NAND2_X1  g626(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n809), .A2(new_n467), .A3(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n809), .A2(new_n467), .B1(new_n815), .B2(new_n813), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n464), .A2(new_n696), .A3(new_n447), .A4(new_n378), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n791), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  INV_X1    g634(.A(G952), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n255), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT122), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n726), .A2(new_n747), .A3(new_n751), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n751), .B1(new_n726), .B2(new_n747), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n663), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n650), .A2(new_n468), .A3(new_n661), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n684), .A2(new_n760), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n732), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n697), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT52), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n830), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n753), .A2(new_n832), .A3(new_n833), .A4(new_n663), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n621), .A2(KEYINPUT114), .A3(new_n627), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n571), .A2(new_n693), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n621), .A2(new_n609), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n685), .A2(new_n305), .A3(new_n306), .A4(new_n638), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n616), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n741), .A2(new_n842), .A3(new_n652), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n611), .A2(new_n724), .A3(new_n727), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n720), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n609), .A2(new_n661), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n846), .B(new_n549), .C1(new_n635), .C2(new_n634), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n513), .B2(new_n519), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n656), .A3(new_n757), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n747), .A2(new_n760), .A3(new_n757), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n782), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n775), .B2(new_n779), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n835), .A2(new_n854), .A3(KEYINPUT53), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  INV_X1    g670(.A(new_n761), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n770), .A2(new_n773), .A3(new_n377), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n773), .B1(new_n770), .B2(new_n377), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n851), .B1(new_n860), .B2(new_n778), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n720), .A3(new_n843), .A4(new_n844), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n831), .A2(new_n834), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n856), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n855), .A2(new_n864), .A3(KEYINPUT115), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n835), .A2(new_n854), .A3(new_n866), .A4(KEYINPUT53), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n865), .A2(KEYINPUT54), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n855), .A2(new_n864), .A3(KEYINPUT116), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n870), .B(new_n856), .C1(new_n862), .C2(new_n863), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT54), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n575), .A2(new_n784), .A3(new_n786), .A4(new_n739), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n791), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT117), .Z(new_n876));
  AND2_X1   g690(.A1(new_n702), .A2(new_n517), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n877), .A2(new_n468), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n817), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n704), .A2(new_n706), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n881), .B2(new_n791), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n791), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n744), .A2(new_n746), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n787), .A2(new_n575), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n684), .A2(new_n378), .A3(new_n574), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n571), .A2(new_n693), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  INV_X1    g707(.A(new_n677), .ZN(new_n894));
  NOR2_X1   g708(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n712), .A2(new_n685), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n894), .A2(new_n896), .A3(new_n874), .A4(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n874), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n674), .B2(new_n676), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n895), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n893), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n879), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n885), .A2(new_n887), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n858), .A2(new_n859), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n905), .A2(KEYINPUT48), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT48), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n885), .A2(new_n628), .A3(new_n889), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n821), .B(G953), .C1(new_n874), .C2(new_n726), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n904), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n898), .A2(new_n901), .A3(KEYINPUT119), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT119), .B1(new_n898), .B2(new_n901), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n892), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n892), .B(new_n918), .C1(new_n914), .C2(new_n915), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n919), .A3(new_n879), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n913), .B1(new_n893), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n823), .B1(new_n873), .B2(new_n921), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n785), .A2(new_n684), .A3(new_n378), .A4(new_n756), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n877), .B(KEYINPUT49), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n894), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT123), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n920), .A2(new_n893), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n909), .A2(new_n912), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n879), .B2(new_n903), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n932), .A2(new_n868), .A3(new_n872), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n928), .B(new_n925), .C1(new_n933), .C2(new_n823), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n927), .A2(new_n934), .ZN(G75));
  NAND2_X1  g749(.A1(new_n869), .A2(new_n871), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n266), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(G210), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n233), .A2(new_n260), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(new_n258), .Z(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT55), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n938), .B2(new_n939), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n321), .A2(G952), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(G51));
  XNOR2_X1  g760(.A(new_n936), .B(KEYINPUT54), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n758), .B(KEYINPUT57), .ZN(new_n948));
  OAI22_X1  g762(.A1(new_n947), .A2(new_n948), .B1(new_n516), .B2(new_n515), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n937), .A2(new_n806), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(G54));
  NAND3_X1  g765(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  INV_X1    g766(.A(new_n564), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n945), .ZN(G60));
  NOR2_X1   g770(.A1(new_n623), .A2(new_n624), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n873), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT59), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n945), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n958), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n947), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n962), .A2(new_n965), .ZN(G63));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT60), .Z(new_n968));
  NAND4_X1  g782(.A1(new_n869), .A2(new_n648), .A3(new_n871), .A4(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n869), .A2(new_n871), .A3(new_n968), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n963), .B(new_n969), .C1(new_n970), .C2(new_n369), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT61), .B1(new_n969), .B2(KEYINPUT124), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G66));
  INV_X1    g787(.A(new_n577), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n255), .B1(new_n974), .B2(G224), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n845), .B2(new_n321), .ZN(new_n976));
  INV_X1    g790(.A(G898), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n940), .B1(new_n977), .B2(new_n318), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n976), .B(new_n978), .ZN(G69));
  INV_X1    g793(.A(new_n811), .ZN(new_n980));
  INV_X1    g794(.A(new_n732), .ZN(new_n981));
  OR3_X1    g795(.A1(new_n810), .A2(new_n981), .A3(new_n906), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n753), .A2(new_n663), .A3(new_n697), .ZN(new_n983));
  INV_X1    g797(.A(new_n782), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n983), .A2(new_n780), .A3(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n819), .A2(new_n980), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n986), .A2(new_n318), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n402), .B1(new_n408), .B2(KEYINPUT30), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(new_n555), .Z(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(G900), .B2(new_n318), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT127), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n666), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n992), .A2(new_n465), .A3(new_n791), .A4(new_n840), .ZN(new_n993));
  INV_X1    g807(.A(new_n983), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n691), .A2(KEYINPUT62), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT62), .B1(new_n691), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n819), .A2(new_n980), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n321), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n989), .B(KEYINPUT125), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1000), .B1(new_n999), .B2(new_n1002), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n991), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n321), .B1(G227), .B2(G900), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1006), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n991), .B(new_n1008), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(new_n986), .B2(new_n845), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n412), .A2(new_n417), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n678), .A2(new_n1012), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1016), .A2(new_n1014), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n865), .A2(new_n867), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(new_n963), .A3(new_n1018), .ZN(new_n1019));
  OR3_X1    g833(.A1(new_n997), .A2(new_n845), .A3(new_n998), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n678), .B1(new_n1020), .B2(new_n1012), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1019), .A2(new_n1021), .ZN(G57));
endmodule


