

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U545 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U546 ( .A(n689), .B(n688), .ZN(n719) );
  XNOR2_X1 U547 ( .A(KEYINPUT100), .B(KEYINPUT30), .ZN(n507) );
  XOR2_X1 U548 ( .A(G543), .B(KEYINPUT0), .Z(n508) );
  XOR2_X1 U549 ( .A(n760), .B(KEYINPUT94), .Z(n509) );
  INV_X1 U550 ( .A(n721), .ZN(n700) );
  INV_X1 U551 ( .A(G168), .ZN(n684) );
  NOR2_X1 U552 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U553 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n688) );
  INV_X1 U554 ( .A(KEYINPUT96), .ZN(n680) );
  XNOR2_X1 U555 ( .A(n729), .B(KEYINPUT32), .ZN(n752) );
  NAND2_X1 U556 ( .A1(n765), .A2(n674), .ZN(n721) );
  INV_X1 U557 ( .A(KEYINPUT103), .ZN(n747) );
  XNOR2_X1 U558 ( .A(n748), .B(n747), .ZN(n749) );
  NAND2_X1 U559 ( .A1(n761), .A2(n509), .ZN(n762) );
  NOR2_X1 U560 ( .A1(G651), .A2(n633), .ZN(n644) );
  XOR2_X1 U561 ( .A(KEYINPUT73), .B(n577), .Z(n909) );
  NOR2_X1 U562 ( .A1(n519), .A2(n518), .ZN(G160) );
  AND2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U564 ( .A1(n882), .A2(G113), .ZN(n513) );
  INV_X1 U565 ( .A(G2105), .ZN(n514) );
  AND2_X1 U566 ( .A1(G2104), .A2(n514), .ZN(n510) );
  XNOR2_X2 U567 ( .A(n510), .B(KEYINPUT64), .ZN(n886) );
  NAND2_X1 U568 ( .A1(n886), .A2(G101), .ZN(n511) );
  XOR2_X1 U569 ( .A(KEYINPUT23), .B(n511), .Z(n512) );
  NAND2_X1 U570 ( .A1(n513), .A2(n512), .ZN(n519) );
  NOR2_X1 U571 ( .A1(G2104), .A2(n514), .ZN(n883) );
  NAND2_X1 U572 ( .A1(G125), .A2(n883), .ZN(n517) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  XOR2_X2 U574 ( .A(KEYINPUT17), .B(n515), .Z(n888) );
  NAND2_X1 U575 ( .A1(G137), .A2(n888), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U577 ( .A1(G543), .A2(G651), .ZN(n636) );
  NAND2_X1 U578 ( .A1(n636), .A2(G89), .ZN(n520) );
  XNOR2_X1 U579 ( .A(n520), .B(KEYINPUT4), .ZN(n524) );
  XNOR2_X1 U580 ( .A(KEYINPUT66), .B(n508), .ZN(n633) );
  INV_X1 U581 ( .A(G651), .ZN(n526) );
  OR2_X1 U582 ( .A1(n633), .A2(n526), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n521), .B(KEYINPUT67), .ZN(n566) );
  INV_X1 U584 ( .A(n566), .ZN(n522) );
  INV_X1 U585 ( .A(n522), .ZN(n640) );
  NAND2_X1 U586 ( .A1(G76), .A2(n640), .ZN(n523) );
  NAND2_X1 U587 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n525), .B(KEYINPUT5), .ZN(n532) );
  NOR2_X1 U589 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n527), .Z(n637) );
  NAND2_X1 U591 ( .A1(G63), .A2(n637), .ZN(n529) );
  NAND2_X1 U592 ( .A1(G51), .A2(n644), .ZN(n528) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U594 ( .A(KEYINPUT6), .B(n530), .Z(n531) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n533), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U597 ( .A1(G138), .A2(n888), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(KEYINPUT88), .ZN(n536) );
  NAND2_X1 U599 ( .A1(n882), .A2(G114), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U601 ( .A1(G126), .A2(n883), .ZN(n538) );
  NAND2_X1 U602 ( .A1(G102), .A2(n886), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n540), .A2(n539), .ZN(G164) );
  NAND2_X1 U605 ( .A1(G91), .A2(n636), .ZN(n542) );
  NAND2_X1 U606 ( .A1(G78), .A2(n640), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U608 ( .A1(G65), .A2(n637), .ZN(n544) );
  NAND2_X1 U609 ( .A1(G53), .A2(n644), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(G299) );
  NAND2_X1 U612 ( .A1(G64), .A2(n637), .ZN(n548) );
  NAND2_X1 U613 ( .A1(G52), .A2(n644), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n640), .A2(G77), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT68), .ZN(n551) );
  NAND2_X1 U617 ( .A1(G90), .A2(n636), .ZN(n550) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(KEYINPUT69), .B(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(KEYINPUT9), .B(n553), .ZN(n554) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(G171) );
  AND2_X1 U622 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  NAND2_X1 U625 ( .A1(G88), .A2(n636), .ZN(n557) );
  NAND2_X1 U626 ( .A1(G75), .A2(n640), .ZN(n556) );
  NAND2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G62), .A2(n637), .ZN(n559) );
  NAND2_X1 U629 ( .A1(G50), .A2(n644), .ZN(n558) );
  NAND2_X1 U630 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U631 ( .A(KEYINPUT83), .B(n560), .Z(n561) );
  NOR2_X1 U632 ( .A1(n562), .A2(n561), .ZN(G166) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U635 ( .A(n563), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U636 ( .A(G223), .ZN(n825) );
  NAND2_X1 U637 ( .A1(n825), .A2(G567), .ZN(n564) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U639 ( .A1(n637), .A2(G56), .ZN(n565) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n565), .Z(n573) );
  NAND2_X1 U641 ( .A1(n566), .A2(G68), .ZN(n567) );
  XNOR2_X1 U642 ( .A(n567), .B(KEYINPUT71), .ZN(n570) );
  NAND2_X1 U643 ( .A1(n636), .A2(G81), .ZN(n568) );
  XOR2_X1 U644 ( .A(KEYINPUT12), .B(n568), .Z(n569) );
  NOR2_X1 U645 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U646 ( .A(n571), .B(KEYINPUT13), .ZN(n572) );
  NOR2_X1 U647 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U648 ( .A(n574), .B(KEYINPUT72), .ZN(n576) );
  NAND2_X1 U649 ( .A1(G43), .A2(n644), .ZN(n575) );
  NAND2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  INV_X1 U651 ( .A(n909), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n578), .A2(G860), .ZN(G153) );
  INV_X1 U653 ( .A(G171), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G92), .A2(n636), .ZN(n580) );
  NAND2_X1 U656 ( .A1(G66), .A2(n637), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U658 ( .A(KEYINPUT74), .B(n581), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G79), .A2(n640), .ZN(n583) );
  NAND2_X1 U660 ( .A1(G54), .A2(n644), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n586), .Z(n587) );
  XNOR2_X1 U664 ( .A(KEYINPUT75), .B(n587), .ZN(n918) );
  INV_X1 U665 ( .A(G868), .ZN(n654) );
  NAND2_X1 U666 ( .A1(n918), .A2(n654), .ZN(n588) );
  NAND2_X1 U667 ( .A1(n589), .A2(n588), .ZN(G284) );
  NOR2_X1 U668 ( .A1(G286), .A2(n654), .ZN(n591) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n590) );
  NOR2_X1 U670 ( .A1(n591), .A2(n590), .ZN(G297) );
  INV_X1 U671 ( .A(G559), .ZN(n595) );
  NOR2_X1 U672 ( .A1(G860), .A2(n595), .ZN(n592) );
  XNOR2_X1 U673 ( .A(n592), .B(KEYINPUT76), .ZN(n593) );
  NOR2_X1 U674 ( .A1(n918), .A2(n593), .ZN(n594) );
  XOR2_X1 U675 ( .A(KEYINPUT16), .B(n594), .Z(G148) );
  INV_X1 U676 ( .A(n918), .ZN(n618) );
  NAND2_X1 U677 ( .A1(n595), .A2(n618), .ZN(n596) );
  NAND2_X1 U678 ( .A1(n596), .A2(G868), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n909), .A2(n654), .ZN(n597) );
  NAND2_X1 U680 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G123), .A2(n883), .ZN(n599) );
  XOR2_X1 U682 ( .A(KEYINPUT18), .B(n599), .Z(n604) );
  NAND2_X1 U683 ( .A1(G111), .A2(n882), .ZN(n601) );
  NAND2_X1 U684 ( .A1(G99), .A2(n886), .ZN(n600) );
  NAND2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U686 ( .A(KEYINPUT77), .B(n602), .Z(n603) );
  NOR2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n888), .A2(G135), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n606), .A2(n605), .ZN(n969) );
  XOR2_X1 U690 ( .A(G2096), .B(KEYINPUT78), .Z(n607) );
  XNOR2_X1 U691 ( .A(n969), .B(n607), .ZN(n609) );
  INV_X1 U692 ( .A(G2100), .ZN(n608) );
  NAND2_X1 U693 ( .A1(n609), .A2(n608), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G93), .A2(n636), .ZN(n611) );
  NAND2_X1 U695 ( .A1(G80), .A2(n640), .ZN(n610) );
  NAND2_X1 U696 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U697 ( .A(n612), .B(KEYINPUT79), .ZN(n614) );
  NAND2_X1 U698 ( .A1(G67), .A2(n637), .ZN(n613) );
  NAND2_X1 U699 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U700 ( .A1(n644), .A2(G55), .ZN(n615) );
  XOR2_X1 U701 ( .A(KEYINPUT80), .B(n615), .Z(n616) );
  OR2_X1 U702 ( .A1(n617), .A2(n616), .ZN(n655) );
  NAND2_X1 U703 ( .A1(G559), .A2(n618), .ZN(n619) );
  XNOR2_X1 U704 ( .A(n619), .B(n909), .ZN(n652) );
  NOR2_X1 U705 ( .A1(G860), .A2(n652), .ZN(n620) );
  XOR2_X1 U706 ( .A(KEYINPUT81), .B(n620), .Z(n621) );
  XOR2_X1 U707 ( .A(n655), .B(n621), .Z(G145) );
  NAND2_X1 U708 ( .A1(G72), .A2(n640), .ZN(n623) );
  NAND2_X1 U709 ( .A1(G47), .A2(n644), .ZN(n622) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U711 ( .A1(G85), .A2(n636), .ZN(n624) );
  XNOR2_X1 U712 ( .A(KEYINPUT65), .B(n624), .ZN(n625) );
  NOR2_X1 U713 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U714 ( .A1(n637), .A2(G60), .ZN(n627) );
  NAND2_X1 U715 ( .A1(n628), .A2(n627), .ZN(G290) );
  NAND2_X1 U716 ( .A1(G49), .A2(n644), .ZN(n630) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U718 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U719 ( .A(KEYINPUT82), .B(n631), .ZN(n632) );
  NOR2_X1 U720 ( .A1(n637), .A2(n632), .ZN(n635) );
  NAND2_X1 U721 ( .A1(G87), .A2(n633), .ZN(n634) );
  NAND2_X1 U722 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U723 ( .A1(G86), .A2(n636), .ZN(n639) );
  NAND2_X1 U724 ( .A1(G61), .A2(n637), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n640), .A2(G73), .ZN(n641) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(n641), .Z(n642) );
  NOR2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n644), .A2(G48), .ZN(n645) );
  NAND2_X1 U730 ( .A1(n646), .A2(n645), .ZN(G305) );
  XNOR2_X1 U731 ( .A(G166), .B(G290), .ZN(n649) );
  XNOR2_X1 U732 ( .A(n655), .B(G305), .ZN(n647) );
  XNOR2_X1 U733 ( .A(G288), .B(n647), .ZN(n648) );
  XNOR2_X1 U734 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U735 ( .A(KEYINPUT19), .B(n650), .ZN(n651) );
  XNOR2_X1 U736 ( .A(n651), .B(G299), .ZN(n834) );
  XNOR2_X1 U737 ( .A(n652), .B(n834), .ZN(n653) );
  NAND2_X1 U738 ( .A1(n653), .A2(G868), .ZN(n657) );
  NAND2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n658) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U745 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U747 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NAND2_X1 U748 ( .A1(G108), .A2(G120), .ZN(n662) );
  NOR2_X1 U749 ( .A1(G237), .A2(n662), .ZN(n663) );
  NAND2_X1 U750 ( .A1(G69), .A2(n663), .ZN(n831) );
  NAND2_X1 U751 ( .A1(G567), .A2(n831), .ZN(n664) );
  XNOR2_X1 U752 ( .A(n664), .B(KEYINPUT86), .ZN(n671) );
  NOR2_X1 U753 ( .A1(G220), .A2(G219), .ZN(n666) );
  XNOR2_X1 U754 ( .A(KEYINPUT22), .B(KEYINPUT84), .ZN(n665) );
  XNOR2_X1 U755 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U756 ( .A1(n667), .A2(G96), .ZN(n668) );
  NOR2_X1 U757 ( .A1(G218), .A2(n668), .ZN(n669) );
  XNOR2_X1 U758 ( .A(KEYINPUT85), .B(n669), .ZN(n832) );
  NAND2_X1 U759 ( .A1(G2106), .A2(n832), .ZN(n670) );
  NAND2_X1 U760 ( .A1(n671), .A2(n670), .ZN(n833) );
  NAND2_X1 U761 ( .A1(G661), .A2(G483), .ZN(n672) );
  XOR2_X1 U762 ( .A(KEYINPUT87), .B(n672), .Z(n673) );
  NOR2_X1 U763 ( .A1(n833), .A2(n673), .ZN(n830) );
  NAND2_X1 U764 ( .A1(n830), .A2(G36), .ZN(G176) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  XOR2_X1 U766 ( .A(G1981), .B(G305), .Z(n906) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n765) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n764) );
  INV_X1 U769 ( .A(n764), .ZN(n674) );
  NAND2_X1 U770 ( .A1(G8), .A2(n721), .ZN(n759) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n741) );
  NAND2_X1 U772 ( .A1(n741), .A2(KEYINPUT33), .ZN(n675) );
  NOR2_X1 U773 ( .A1(n759), .A2(n675), .ZN(n676) );
  XOR2_X1 U774 ( .A(KEYINPUT104), .B(n676), .Z(n677) );
  NAND2_X1 U775 ( .A1(n906), .A2(n677), .ZN(n750) );
  XNOR2_X1 U776 ( .A(KEYINPUT25), .B(G2078), .ZN(n937) );
  NOR2_X1 U777 ( .A1(n721), .A2(n937), .ZN(n679) );
  INV_X1 U778 ( .A(G1961), .ZN(n983) );
  NOR2_X1 U779 ( .A1(n700), .A2(n983), .ZN(n678) );
  NOR2_X1 U780 ( .A1(n679), .A2(n678), .ZN(n715) );
  NOR2_X1 U781 ( .A1(G171), .A2(n715), .ZN(n687) );
  NOR2_X1 U782 ( .A1(G2084), .A2(n721), .ZN(n731) );
  NOR2_X1 U783 ( .A1(G1966), .A2(n759), .ZN(n681) );
  XNOR2_X1 U784 ( .A(n681), .B(n680), .ZN(n734) );
  NAND2_X1 U785 ( .A1(n734), .A2(G8), .ZN(n682) );
  NOR2_X1 U786 ( .A1(n731), .A2(n682), .ZN(n683) );
  XNOR2_X1 U787 ( .A(n683), .B(n507), .ZN(n685) );
  NOR2_X1 U788 ( .A1(n687), .A2(n686), .ZN(n689) );
  AND2_X1 U789 ( .A1(n700), .A2(G1996), .ZN(n691) );
  XOR2_X1 U790 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n690) );
  XNOR2_X1 U791 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U792 ( .A1(n721), .A2(G1341), .ZN(n692) );
  NAND2_X1 U793 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U794 ( .A1(n909), .A2(n694), .ZN(n698) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n721), .ZN(n696) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n700), .ZN(n695) );
  NAND2_X1 U797 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U798 ( .A1(n699), .A2(n918), .ZN(n697) );
  NAND2_X1 U799 ( .A1(n698), .A2(n697), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n918), .A2(n699), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n700), .A2(G2072), .ZN(n701) );
  XOR2_X1 U802 ( .A(KEYINPUT27), .B(n701), .Z(n704) );
  NAND2_X1 U803 ( .A1(G1956), .A2(n721), .ZN(n702) );
  XOR2_X1 U804 ( .A(KEYINPUT97), .B(n702), .Z(n703) );
  NAND2_X1 U805 ( .A1(n704), .A2(n703), .ZN(n710) );
  NOR2_X1 U806 ( .A1(n710), .A2(G299), .ZN(n705) );
  NOR2_X1 U807 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U808 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U809 ( .A(KEYINPUT99), .B(n709), .ZN(n713) );
  NAND2_X1 U810 ( .A1(G299), .A2(n710), .ZN(n711) );
  XOR2_X1 U811 ( .A(KEYINPUT28), .B(n711), .Z(n712) );
  XNOR2_X1 U812 ( .A(n714), .B(KEYINPUT29), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n715), .A2(G171), .ZN(n716) );
  NAND2_X1 U814 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n719), .A2(n718), .ZN(n730) );
  AND2_X1 U816 ( .A1(G286), .A2(G8), .ZN(n720) );
  NAND2_X1 U817 ( .A1(n730), .A2(n720), .ZN(n728) );
  INV_X1 U818 ( .A(G8), .ZN(n726) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n759), .ZN(n723) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n721), .ZN(n722) );
  NOR2_X1 U821 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U822 ( .A1(n724), .A2(G303), .ZN(n725) );
  OR2_X1 U823 ( .A1(n726), .A2(n725), .ZN(n727) );
  AND2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U825 ( .A(n730), .B(KEYINPUT102), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n731), .A2(G8), .ZN(n732) );
  XOR2_X1 U827 ( .A(KEYINPUT95), .B(n732), .Z(n733) );
  AND2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n751) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n915) );
  INV_X1 U831 ( .A(n759), .ZN(n737) );
  NAND2_X1 U832 ( .A1(n915), .A2(n737), .ZN(n742) );
  INV_X1 U833 ( .A(n742), .ZN(n738) );
  AND2_X1 U834 ( .A1(n751), .A2(n738), .ZN(n739) );
  NAND2_X1 U835 ( .A1(n752), .A2(n739), .ZN(n746) );
  INV_X1 U836 ( .A(KEYINPUT33), .ZN(n744) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n740) );
  NOR2_X1 U838 ( .A1(n741), .A2(n740), .ZN(n923) );
  OR2_X1 U839 ( .A1(n742), .A2(n923), .ZN(n743) );
  AND2_X1 U840 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U841 ( .A1(n746), .A2(n745), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n763) );
  NAND2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n755) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n753) );
  NAND2_X1 U845 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n756), .A2(n759), .ZN(n761) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n757) );
  XOR2_X1 U849 ( .A(n757), .B(KEYINPUT24), .Z(n758) );
  NOR2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  OR2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n799) );
  XNOR2_X1 U852 ( .A(G1986), .B(G290), .ZN(n917) );
  NOR2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n810) );
  NAND2_X1 U854 ( .A1(n917), .A2(n810), .ZN(n797) );
  NAND2_X1 U855 ( .A1(G131), .A2(n888), .ZN(n767) );
  NAND2_X1 U856 ( .A1(G95), .A2(n886), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n771) );
  NAND2_X1 U858 ( .A1(G107), .A2(n882), .ZN(n769) );
  NAND2_X1 U859 ( .A1(G119), .A2(n883), .ZN(n768) );
  NAND2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U862 ( .A(n772), .B(KEYINPUT91), .ZN(n879) );
  NAND2_X1 U863 ( .A1(G1991), .A2(n879), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G117), .A2(n882), .ZN(n774) );
  NAND2_X1 U865 ( .A1(G129), .A2(n883), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n886), .A2(G105), .ZN(n775) );
  XOR2_X1 U868 ( .A(KEYINPUT38), .B(n775), .Z(n776) );
  NOR2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n888), .A2(G141), .ZN(n778) );
  NAND2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n865) );
  NAND2_X1 U872 ( .A1(G1996), .A2(n865), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U874 ( .A(KEYINPUT92), .B(n782), .Z(n965) );
  XNOR2_X1 U875 ( .A(n810), .B(KEYINPUT93), .ZN(n783) );
  NOR2_X1 U876 ( .A1(n965), .A2(n783), .ZN(n802) );
  INV_X1 U877 ( .A(n802), .ZN(n795) );
  XNOR2_X1 U878 ( .A(G2067), .B(KEYINPUT37), .ZN(n808) );
  NAND2_X1 U879 ( .A1(G104), .A2(n886), .ZN(n784) );
  XOR2_X1 U880 ( .A(KEYINPUT89), .B(n784), .Z(n786) );
  NAND2_X1 U881 ( .A1(n888), .A2(G140), .ZN(n785) );
  NAND2_X1 U882 ( .A1(n786), .A2(n785), .ZN(n788) );
  XNOR2_X1 U883 ( .A(KEYINPUT90), .B(KEYINPUT34), .ZN(n787) );
  XNOR2_X1 U884 ( .A(n788), .B(n787), .ZN(n793) );
  NAND2_X1 U885 ( .A1(G116), .A2(n882), .ZN(n790) );
  NAND2_X1 U886 ( .A1(G128), .A2(n883), .ZN(n789) );
  NAND2_X1 U887 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U888 ( .A(KEYINPUT35), .B(n791), .Z(n792) );
  NOR2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U890 ( .A(KEYINPUT36), .B(n794), .ZN(n896) );
  NOR2_X1 U891 ( .A1(n808), .A2(n896), .ZN(n976) );
  NAND2_X1 U892 ( .A1(n810), .A2(n976), .ZN(n806) );
  AND2_X1 U893 ( .A1(n795), .A2(n806), .ZN(n796) );
  AND2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n813) );
  XOR2_X1 U896 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n805) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n865), .ZN(n961) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n879), .ZN(n968) );
  NOR2_X1 U900 ( .A1(n800), .A2(n968), .ZN(n801) );
  NOR2_X1 U901 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U902 ( .A1(n961), .A2(n803), .ZN(n804) );
  XNOR2_X1 U903 ( .A(n805), .B(n804), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n808), .A2(n896), .ZN(n973) );
  NAND2_X1 U906 ( .A1(n809), .A2(n973), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U909 ( .A(KEYINPUT40), .B(n814), .ZN(G329) );
  XNOR2_X1 U910 ( .A(G2430), .B(G2454), .ZN(n823) );
  XNOR2_X1 U911 ( .A(KEYINPUT106), .B(G2435), .ZN(n821) );
  XOR2_X1 U912 ( .A(G2451), .B(G2427), .Z(n816) );
  XNOR2_X1 U913 ( .A(G2438), .B(G2446), .ZN(n815) );
  XNOR2_X1 U914 ( .A(n816), .B(n815), .ZN(n817) );
  XOR2_X1 U915 ( .A(n817), .B(G2443), .Z(n819) );
  XNOR2_X1 U916 ( .A(G1348), .B(G1341), .ZN(n818) );
  XNOR2_X1 U917 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U918 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U919 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n824), .A2(G14), .ZN(n901) );
  XNOR2_X1 U921 ( .A(KEYINPUT107), .B(n901), .ZN(G401) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n825), .ZN(G217) );
  NAND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n826) );
  XOR2_X1 U924 ( .A(KEYINPUT108), .B(n826), .Z(n827) );
  NAND2_X1 U925 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n828) );
  XOR2_X1 U927 ( .A(KEYINPUT109), .B(n828), .Z(n829) );
  NAND2_X1 U928 ( .A1(n830), .A2(n829), .ZN(G188) );
  XOR2_X1 U929 ( .A(G120), .B(KEYINPUT110), .Z(G236) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(KEYINPUT111), .B(n833), .ZN(G319) );
  XNOR2_X1 U936 ( .A(G286), .B(n909), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n918), .B(G171), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  NOR2_X1 U940 ( .A1(G37), .A2(n838), .ZN(G397) );
  XNOR2_X1 U941 ( .A(G1996), .B(G2474), .ZN(n848) );
  XOR2_X1 U942 ( .A(G1956), .B(G1961), .Z(n840) );
  XNOR2_X1 U943 ( .A(G1991), .B(G1981), .ZN(n839) );
  XNOR2_X1 U944 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U945 ( .A(G1966), .B(G1971), .Z(n842) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1976), .ZN(n841) );
  XNOR2_X1 U947 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U948 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U949 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n845) );
  XNOR2_X1 U950 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U952 ( .A(G2100), .B(G2096), .Z(n850) );
  XNOR2_X1 U953 ( .A(KEYINPUT42), .B(G2678), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U955 ( .A(KEYINPUT43), .B(G2090), .Z(n852) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U957 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U958 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U959 ( .A(G2084), .B(G2078), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n856), .B(n855), .ZN(G227) );
  NAND2_X1 U961 ( .A1(G124), .A2(n883), .ZN(n857) );
  XNOR2_X1 U962 ( .A(n857), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U963 ( .A1(G136), .A2(n888), .ZN(n858) );
  XOR2_X1 U964 ( .A(KEYINPUT113), .B(n858), .Z(n859) );
  NAND2_X1 U965 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G112), .A2(n882), .ZN(n862) );
  NAND2_X1 U967 ( .A1(G100), .A2(n886), .ZN(n861) );
  NAND2_X1 U968 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U969 ( .A1(n864), .A2(n863), .ZN(G162) );
  XNOR2_X1 U970 ( .A(G160), .B(n865), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n866), .B(n969), .ZN(n878) );
  XOR2_X1 U972 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n876) );
  NAND2_X1 U973 ( .A1(G139), .A2(n888), .ZN(n868) );
  NAND2_X1 U974 ( .A1(G103), .A2(n886), .ZN(n867) );
  NAND2_X1 U975 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G115), .A2(n882), .ZN(n870) );
  NAND2_X1 U977 ( .A1(G127), .A2(n883), .ZN(n869) );
  NAND2_X1 U978 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U979 ( .A(KEYINPUT115), .B(n871), .ZN(n872) );
  XNOR2_X1 U980 ( .A(KEYINPUT47), .B(n872), .ZN(n873) );
  NOR2_X1 U981 ( .A1(n874), .A2(n873), .ZN(n954) );
  XNOR2_X1 U982 ( .A(n954), .B(G162), .ZN(n875) );
  XNOR2_X1 U983 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U984 ( .A(n878), .B(n877), .ZN(n881) );
  XNOR2_X1 U985 ( .A(n879), .B(G164), .ZN(n880) );
  XNOR2_X1 U986 ( .A(n881), .B(n880), .ZN(n895) );
  NAND2_X1 U987 ( .A1(G118), .A2(n882), .ZN(n885) );
  NAND2_X1 U988 ( .A1(G130), .A2(n883), .ZN(n884) );
  NAND2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n893) );
  NAND2_X1 U990 ( .A1(G106), .A2(n886), .ZN(n887) );
  XNOR2_X1 U991 ( .A(n887), .B(KEYINPUT114), .ZN(n890) );
  NAND2_X1 U992 ( .A1(G142), .A2(n888), .ZN(n889) );
  NAND2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U994 ( .A(n891), .B(KEYINPUT45), .Z(n892) );
  NOR2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(n895), .B(n894), .Z(n897) );
  XOR2_X1 U997 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U998 ( .A1(G37), .A2(n898), .ZN(G395) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n899) );
  XOR2_X1 U1000 ( .A(KEYINPUT49), .B(n899), .Z(n900) );
  NAND2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n902) );
  NOR2_X1 U1002 ( .A1(G397), .A2(n902), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n903), .ZN(n904) );
  NOR2_X1 U1004 ( .A1(n904), .A2(G395), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n905), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1006 ( .A(G308), .ZN(G225) );
  INV_X1 U1007 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1008 ( .A(G16), .B(KEYINPUT56), .Z(n928) );
  XNOR2_X1 U1009 ( .A(G1966), .B(G168), .ZN(n907) );
  NAND2_X1 U1010 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1011 ( .A(n908), .B(KEYINPUT57), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(G301), .B(G1961), .ZN(n911) );
  XNOR2_X1 U1013 ( .A(n909), .B(G1341), .ZN(n910) );
  NOR2_X1 U1014 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n926) );
  NAND2_X1 U1016 ( .A1(G1971), .A2(G303), .ZN(n914) );
  NAND2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(G1956), .B(G299), .ZN(n916) );
  NOR2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n920) );
  XOR2_X1 U1020 ( .A(G1348), .B(n918), .Z(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n953) );
  XNOR2_X1 U1026 ( .A(G2084), .B(G34), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n929), .B(KEYINPUT54), .ZN(n945) );
  XNOR2_X1 U1028 ( .A(G2090), .B(G35), .ZN(n942) );
  XNOR2_X1 U1029 ( .A(G1996), .B(G32), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(G33), .B(G2072), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n936) );
  XOR2_X1 U1032 ( .A(G1991), .B(G25), .Z(n932) );
  NAND2_X1 U1033 ( .A1(n932), .A2(G28), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(G26), .B(G2067), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1037 ( .A(G27), .B(n937), .Z(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(KEYINPUT53), .B(n940), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1041 ( .A(KEYINPUT120), .B(n943), .Z(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(KEYINPUT121), .B(n946), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n978) );
  XNOR2_X1 U1045 ( .A(n947), .B(n978), .ZN(n949) );
  INV_X1 U1046 ( .A(G29), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(G11), .A2(n950), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(KEYINPUT122), .B(n951), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n982) );
  XOR2_X1 U1051 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n959) );
  XOR2_X1 U1052 ( .A(G2072), .B(n954), .Z(n956) );
  XOR2_X1 U1053 ( .A(G164), .B(G2078), .Z(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(n957), .B(KEYINPUT50), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(n959), .B(n958), .ZN(n964) );
  XOR2_X1 U1057 ( .A(G2090), .B(G162), .Z(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1059 ( .A(KEYINPUT51), .B(n962), .Z(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(G2084), .B(G160), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(KEYINPUT52), .B(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n980), .A2(G29), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n1010) );
  XOR2_X1 U1072 ( .A(G16), .B(KEYINPUT123), .Z(n1008) );
  XNOR2_X1 U1073 ( .A(G5), .B(n983), .ZN(n998) );
  XOR2_X1 U1074 ( .A(G1981), .B(G6), .Z(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(G19), .B(G1341), .ZN(n985) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(n987), .B(KEYINPUT126), .ZN(n990) );
  XOR2_X1 U1079 ( .A(G1956), .B(KEYINPUT124), .Z(n988) );
  XNOR2_X1 U1080 ( .A(G20), .B(n988), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1082 ( .A(KEYINPUT59), .B(G1348), .Z(n991) );
  XNOR2_X1 U1083 ( .A(G4), .B(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1085 ( .A(KEYINPUT60), .B(n994), .Z(n996) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G21), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(G1976), .B(G23), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G22), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(G1986), .B(G24), .Z(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1006), .Z(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1011), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

