

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U548 ( .A(n680), .B(KEYINPUT64), .ZN(n682) );
  BUF_X2 U549 ( .A(n888), .Z(n513) );
  XOR2_X1 U550 ( .A(KEYINPUT17), .B(n516), .Z(n888) );
  INV_X2 U551 ( .A(n697), .ZN(n735) );
  INV_X1 U552 ( .A(n682), .ZN(n697) );
  NAND2_X1 U553 ( .A1(G160), .A2(G40), .ZN(n809) );
  NOR2_X1 U554 ( .A1(G164), .A2(G1384), .ZN(n810) );
  INV_X1 U555 ( .A(KEYINPUT28), .ZN(n686) );
  NOR2_X1 U556 ( .A1(n723), .A2(n722), .ZN(n725) );
  XNOR2_X1 U557 ( .A(n718), .B(KEYINPUT30), .ZN(n719) );
  INV_X1 U558 ( .A(KEYINPUT31), .ZN(n724) );
  INV_X1 U559 ( .A(KEYINPUT76), .ZN(n600) );
  INV_X1 U560 ( .A(KEYINPUT104), .ZN(n765) );
  XNOR2_X1 U561 ( .A(n600), .B(KEYINPUT15), .ZN(n601) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  NOR2_X1 U563 ( .A1(G651), .A2(n633), .ZN(n650) );
  INV_X1 U564 ( .A(G2105), .ZN(n514) );
  AND2_X4 U565 ( .A1(n514), .A2(G2104), .ZN(n887) );
  NAND2_X1 U566 ( .A1(n887), .A2(G102), .ZN(n515) );
  XNOR2_X1 U567 ( .A(n515), .B(KEYINPUT90), .ZN(n518) );
  NAND2_X1 U568 ( .A1(G138), .A2(n513), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n518), .A2(n517), .ZN(n523) );
  INV_X1 U570 ( .A(G2105), .ZN(n519) );
  NOR2_X1 U571 ( .A1(G2104), .A2(n519), .ZN(n883) );
  NAND2_X1 U572 ( .A1(G126), .A2(n883), .ZN(n521) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U574 ( .A1(G114), .A2(n884), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U576 ( .A1(n523), .A2(n522), .ZN(G164) );
  XNOR2_X1 U577 ( .A(KEYINPUT6), .B(KEYINPUT80), .ZN(n530) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  NAND2_X1 U579 ( .A1(n650), .A2(G51), .ZN(n528) );
  INV_X1 U580 ( .A(G651), .ZN(n532) );
  NOR2_X1 U581 ( .A1(G543), .A2(n532), .ZN(n525) );
  XNOR2_X1 U582 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n524) );
  XNOR2_X1 U583 ( .A(n525), .B(n524), .ZN(n642) );
  NAND2_X1 U584 ( .A1(n642), .A2(G63), .ZN(n526) );
  XOR2_X1 U585 ( .A(KEYINPUT79), .B(n526), .Z(n527) );
  NAND2_X1 U586 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U587 ( .A(n530), .B(n529), .Z(n539) );
  XNOR2_X1 U588 ( .A(KEYINPUT78), .B(KEYINPUT5), .ZN(n537) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U590 ( .A1(n645), .A2(G89), .ZN(n531) );
  XNOR2_X1 U591 ( .A(n531), .B(KEYINPUT4), .ZN(n535) );
  OR2_X1 U592 ( .A1(n532), .A2(n633), .ZN(n533) );
  XOR2_X2 U593 ( .A(KEYINPUT66), .B(n533), .Z(n640) );
  NAND2_X1 U594 ( .A1(G76), .A2(n640), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U596 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n540), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U599 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U600 ( .A1(G101), .A2(n887), .ZN(n541) );
  XNOR2_X1 U601 ( .A(n541), .B(KEYINPUT65), .ZN(n542) );
  XNOR2_X1 U602 ( .A(n542), .B(KEYINPUT23), .ZN(n544) );
  NAND2_X1 U603 ( .A1(G113), .A2(n884), .ZN(n543) );
  NAND2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G137), .A2(n513), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G125), .A2(n883), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X2 U608 ( .A1(n548), .A2(n547), .ZN(G160) );
  NAND2_X1 U609 ( .A1(G85), .A2(n645), .ZN(n550) );
  NAND2_X1 U610 ( .A1(G60), .A2(n642), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n650), .A2(G47), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G72), .A2(n640), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U615 ( .A1(n554), .A2(n553), .ZN(G290) );
  NAND2_X1 U616 ( .A1(G64), .A2(n642), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G52), .A2(n650), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U619 ( .A(KEYINPUT68), .B(n557), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n645), .A2(G90), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G77), .A2(n640), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n560), .Z(n561) );
  NOR2_X1 U624 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U625 ( .A1(G111), .A2(n884), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G99), .A2(n887), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G135), .A2(n513), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n883), .A2(G123), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT18), .B(n565), .Z(n566) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT82), .ZN(n971) );
  XNOR2_X1 U634 ( .A(n971), .B(G2096), .ZN(n571) );
  OR2_X1 U635 ( .A1(G2100), .A2(n571), .ZN(G156) );
  INV_X1 U636 ( .A(G57), .ZN(G237) );
  NAND2_X1 U637 ( .A1(n645), .A2(G88), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G75), .A2(n640), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G62), .A2(n642), .ZN(n575) );
  NAND2_X1 U641 ( .A1(G50), .A2(n650), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(G166) );
  NAND2_X1 U644 ( .A1(G94), .A2(G452), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n829) );
  NAND2_X1 U649 ( .A1(n829), .A2(G567), .ZN(n580) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  NAND2_X1 U651 ( .A1(n650), .A2(G43), .ZN(n581) );
  XNOR2_X1 U652 ( .A(KEYINPUT74), .B(n581), .ZN(n592) );
  XNOR2_X1 U653 ( .A(KEYINPUT73), .B(KEYINPUT13), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G81), .A2(n645), .ZN(n582) );
  XNOR2_X1 U655 ( .A(n582), .B(KEYINPUT72), .ZN(n583) );
  XNOR2_X1 U656 ( .A(n583), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G68), .A2(n640), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n587), .B(n586), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n642), .A2(G56), .ZN(n588) );
  XOR2_X1 U661 ( .A(KEYINPUT14), .B(n588), .Z(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n993) );
  INV_X1 U664 ( .A(G860), .ZN(n624) );
  OR2_X1 U665 ( .A1(n993), .A2(n624), .ZN(G153) );
  NAND2_X1 U666 ( .A1(n650), .A2(G54), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n642), .A2(G66), .ZN(n594) );
  NAND2_X1 U668 ( .A1(G79), .A2(n640), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U670 ( .A1(G92), .A2(n645), .ZN(n595) );
  XNOR2_X1 U671 ( .A(KEYINPUT75), .B(n595), .ZN(n596) );
  NOR2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n602) );
  XNOR2_X2 U674 ( .A(n602), .B(n601), .ZN(n1003) );
  INV_X1 U675 ( .A(n1003), .ZN(n622) );
  NOR2_X1 U676 ( .A1(G868), .A2(n622), .ZN(n604) );
  INV_X1 U677 ( .A(G868), .ZN(n661) );
  NOR2_X1 U678 ( .A1(G171), .A2(n661), .ZN(n603) );
  NOR2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U680 ( .A(KEYINPUT77), .B(n605), .ZN(G284) );
  NAND2_X1 U681 ( .A1(G91), .A2(n645), .ZN(n606) );
  XNOR2_X1 U682 ( .A(n606), .B(KEYINPUT70), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n642), .A2(G65), .ZN(n608) );
  NAND2_X1 U684 ( .A1(G78), .A2(n640), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G53), .A2(n650), .ZN(n609) );
  XNOR2_X1 U687 ( .A(KEYINPUT71), .B(n609), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G299) );
  NOR2_X1 U690 ( .A1(G286), .A2(n661), .ZN(n614) );
  XOR2_X1 U691 ( .A(KEYINPUT81), .B(n614), .Z(n616) );
  NOR2_X1 U692 ( .A1(G868), .A2(G299), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n616), .A2(n615), .ZN(G297) );
  NAND2_X1 U694 ( .A1(n624), .A2(G559), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n617), .A2(n622), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n618), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U697 ( .A1(G868), .A2(n993), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(G868), .ZN(n619) );
  NOR2_X1 U699 ( .A1(G559), .A2(n619), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(G282) );
  NAND2_X1 U701 ( .A1(n622), .A2(G559), .ZN(n623) );
  XOR2_X1 U702 ( .A(n993), .B(n623), .Z(n658) );
  NAND2_X1 U703 ( .A1(n624), .A2(n658), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G93), .A2(n645), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G67), .A2(n642), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G55), .A2(n650), .ZN(n627) );
  XNOR2_X1 U708 ( .A(KEYINPUT83), .B(n627), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G80), .A2(n640), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n660) );
  XNOR2_X1 U712 ( .A(n632), .B(n660), .ZN(G145) );
  NAND2_X1 U713 ( .A1(G87), .A2(n633), .ZN(n634) );
  XNOR2_X1 U714 ( .A(n634), .B(KEYINPUT84), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G49), .A2(n650), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n642), .A2(n637), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G73), .A2(n640), .ZN(n641) );
  XNOR2_X1 U721 ( .A(n641), .B(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G61), .A2(n642), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G86), .A2(n645), .ZN(n646) );
  XNOR2_X1 U725 ( .A(KEYINPUT85), .B(n646), .ZN(n647) );
  NOR2_X1 U726 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U727 ( .A(n649), .B(KEYINPUT86), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n650), .A2(G48), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(G305) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(G288), .ZN(n657) );
  INV_X1 U731 ( .A(G299), .ZN(n1000) );
  XNOR2_X1 U732 ( .A(n1000), .B(G305), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n653), .B(n660), .ZN(n654) );
  XNOR2_X1 U734 ( .A(G166), .B(n654), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n655), .B(G290), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n657), .B(n656), .ZN(n906) );
  XNOR2_X1 U737 ( .A(n658), .B(n906), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n659), .A2(G868), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U741 ( .A(KEYINPUT87), .B(n664), .Z(G295) );
  NAND2_X1 U742 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n666), .ZN(n668) );
  XNOR2_X1 U745 ( .A(KEYINPUT88), .B(KEYINPUT21), .ZN(n667) );
  XNOR2_X1 U746 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U747 ( .A1(G2072), .A2(n669), .ZN(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n671) );
  NAND2_X1 U750 ( .A1(G132), .A2(G82), .ZN(n670) );
  XNOR2_X1 U751 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U752 ( .A1(n672), .A2(G218), .ZN(n673) );
  NAND2_X1 U753 ( .A1(G96), .A2(n673), .ZN(n834) );
  NAND2_X1 U754 ( .A1(n834), .A2(G2106), .ZN(n677) );
  NAND2_X1 U755 ( .A1(G120), .A2(G69), .ZN(n674) );
  NOR2_X1 U756 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U757 ( .A1(G108), .A2(n675), .ZN(n835) );
  NAND2_X1 U758 ( .A1(n835), .A2(G567), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n677), .A2(n676), .ZN(n916) );
  NAND2_X1 U760 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U761 ( .A1(n916), .A2(n678), .ZN(n833) );
  NAND2_X1 U762 ( .A1(n833), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  INV_X1 U764 ( .A(n809), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n679), .A2(n810), .ZN(n680) );
  NAND2_X1 U766 ( .A1(G8), .A2(n682), .ZN(n681) );
  XNOR2_X2 U767 ( .A(n681), .B(KEYINPUT98), .ZN(n768) );
  NOR2_X1 U768 ( .A1(n768), .A2(G1966), .ZN(n729) );
  NAND2_X1 U769 ( .A1(G2072), .A2(n697), .ZN(n683) );
  XNOR2_X1 U770 ( .A(n683), .B(KEYINPUT27), .ZN(n685) );
  XNOR2_X1 U771 ( .A(G1956), .B(KEYINPUT99), .ZN(n927) );
  NOR2_X1 U772 ( .A1(n697), .A2(n927), .ZN(n684) );
  NOR2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n705) );
  NOR2_X1 U774 ( .A1(n705), .A2(n1000), .ZN(n687) );
  XNOR2_X1 U775 ( .A(n687), .B(n686), .ZN(n709) );
  NAND2_X1 U776 ( .A1(G2067), .A2(n697), .ZN(n689) );
  NAND2_X1 U777 ( .A1(n735), .A2(G1348), .ZN(n688) );
  NAND2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U779 ( .A1(n1003), .A2(n690), .ZN(n704) );
  NAND2_X1 U780 ( .A1(n1003), .A2(G1348), .ZN(n691) );
  NAND2_X1 U781 ( .A1(KEYINPUT26), .A2(n691), .ZN(n692) );
  NOR2_X1 U782 ( .A1(G1341), .A2(n692), .ZN(n693) );
  NOR2_X1 U783 ( .A1(n697), .A2(n693), .ZN(n702) );
  NAND2_X1 U784 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n695) );
  NAND2_X1 U785 ( .A1(G2067), .A2(n1003), .ZN(n694) );
  NAND2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U788 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n698) );
  NOR2_X1 U789 ( .A1(n993), .A2(n698), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U792 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U793 ( .A1(n705), .A2(n1000), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U795 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U796 ( .A(KEYINPUT29), .B(n710), .Z(n714) );
  AND2_X1 U797 ( .A1(n735), .A2(G1961), .ZN(n712) );
  XNOR2_X1 U798 ( .A(KEYINPUT25), .B(G2078), .ZN(n946) );
  NOR2_X1 U799 ( .A1(n735), .A2(n946), .ZN(n711) );
  NOR2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U801 ( .A1(G171), .A2(n715), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n727) );
  NOR2_X1 U803 ( .A1(G171), .A2(n715), .ZN(n723) );
  NOR2_X1 U804 ( .A1(n735), .A2(G2084), .ZN(n730) );
  INV_X1 U805 ( .A(n730), .ZN(n716) );
  NAND2_X1 U806 ( .A1(G8), .A2(n716), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n729), .A2(n717), .ZN(n720) );
  INV_X1 U808 ( .A(KEYINPUT100), .ZN(n718) );
  XNOR2_X1 U809 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U810 ( .A1(G168), .A2(n721), .ZN(n722) );
  XNOR2_X1 U811 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U812 ( .A1(n727), .A2(n726), .ZN(n734) );
  XNOR2_X1 U813 ( .A(KEYINPUT101), .B(n734), .ZN(n728) );
  NOR2_X1 U814 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U815 ( .A1(G8), .A2(n730), .ZN(n731) );
  NAND2_X1 U816 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U817 ( .A(n733), .B(KEYINPUT102), .ZN(n757) );
  NAND2_X1 U818 ( .A1(n734), .A2(G286), .ZN(n740) );
  NOR2_X1 U819 ( .A1(n768), .A2(G1971), .ZN(n737) );
  NOR2_X1 U820 ( .A1(n735), .A2(G2090), .ZN(n736) );
  NOR2_X1 U821 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U822 ( .A1(n738), .A2(G303), .ZN(n739) );
  NAND2_X1 U823 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U824 ( .A1(G8), .A2(n741), .ZN(n742) );
  XNOR2_X1 U825 ( .A(n742), .B(KEYINPUT32), .ZN(n758) );
  NAND2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  AND2_X1 U827 ( .A1(n758), .A2(n1011), .ZN(n743) );
  NAND2_X1 U828 ( .A1(n757), .A2(n743), .ZN(n748) );
  INV_X1 U829 ( .A(n1011), .ZN(n746) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n1008) );
  NOR2_X1 U832 ( .A1(n744), .A2(n1008), .ZN(n745) );
  OR2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n747) );
  AND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n768), .A2(n749), .ZN(n750) );
  NOR2_X1 U836 ( .A1(KEYINPUT33), .A2(n750), .ZN(n751) );
  XNOR2_X1 U837 ( .A(n751), .B(KEYINPUT103), .ZN(n756) );
  OR2_X1 U838 ( .A1(G1981), .A2(G305), .ZN(n767) );
  NAND2_X1 U839 ( .A1(G1981), .A2(G305), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n767), .A2(n752), .ZN(n997) );
  NAND2_X1 U841 ( .A1(KEYINPUT33), .A2(n1008), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n768), .A2(n753), .ZN(n754) );
  NOR2_X1 U843 ( .A1(n997), .A2(n754), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n764) );
  NAND2_X1 U845 ( .A1(n757), .A2(n758), .ZN(n761) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n768), .A2(n762), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n766) );
  XNOR2_X1 U851 ( .A(n766), .B(n765), .ZN(n817) );
  XOR2_X1 U852 ( .A(n767), .B(KEYINPUT24), .Z(n770) );
  INV_X1 U853 ( .A(n768), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n770), .A2(n769), .ZN(n815) );
  XNOR2_X1 U855 ( .A(G2067), .B(KEYINPUT37), .ZN(n771) );
  XNOR2_X1 U856 ( .A(n771), .B(KEYINPUT91), .ZN(n811) );
  NAND2_X1 U857 ( .A1(G104), .A2(n887), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G140), .A2(n513), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n774), .ZN(n781) );
  NAND2_X1 U861 ( .A1(n884), .A2(G116), .ZN(n775) );
  XNOR2_X1 U862 ( .A(n775), .B(KEYINPUT92), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G128), .A2(n883), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U865 ( .A(KEYINPUT35), .B(n778), .ZN(n779) );
  XNOR2_X1 U866 ( .A(KEYINPUT93), .B(n779), .ZN(n780) );
  NOR2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U868 ( .A(n782), .B(KEYINPUT36), .Z(n783) );
  XNOR2_X1 U869 ( .A(KEYINPUT94), .B(n783), .ZN(n879) );
  NOR2_X1 U870 ( .A1(n811), .A2(n879), .ZN(n973) );
  NAND2_X1 U871 ( .A1(G105), .A2(n887), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT38), .ZN(n791) );
  NAND2_X1 U873 ( .A1(G129), .A2(n883), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G117), .A2(n884), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G141), .A2(n513), .ZN(n787) );
  XNOR2_X1 U877 ( .A(KEYINPUT95), .B(n787), .ZN(n788) );
  NOR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U880 ( .A(KEYINPUT96), .B(n792), .ZN(n880) );
  NOR2_X1 U881 ( .A1(G1996), .A2(n880), .ZN(n793) );
  XOR2_X1 U882 ( .A(KEYINPUT105), .B(n793), .Z(n977) );
  NOR2_X1 U883 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G95), .A2(n887), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G131), .A2(n513), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G119), .A2(n883), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G107), .A2(n884), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n902) );
  NOR2_X1 U891 ( .A1(G1991), .A2(n902), .ZN(n969) );
  NOR2_X1 U892 ( .A1(n800), .A2(n969), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G1996), .A2(n880), .ZN(n801) );
  XOR2_X1 U894 ( .A(KEYINPUT97), .B(n801), .Z(n803) );
  NAND2_X1 U895 ( .A1(G1991), .A2(n902), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n820) );
  NOR2_X1 U897 ( .A1(n804), .A2(n820), .ZN(n805) );
  XNOR2_X1 U898 ( .A(n805), .B(KEYINPUT106), .ZN(n806) );
  NOR2_X1 U899 ( .A1(n977), .A2(n806), .ZN(n807) );
  XNOR2_X1 U900 ( .A(n807), .B(KEYINPUT39), .ZN(n808) );
  NOR2_X1 U901 ( .A1(n973), .A2(n808), .ZN(n813) );
  NOR2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n822) );
  NAND2_X1 U903 ( .A1(n811), .A2(n879), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n822), .A2(n819), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U906 ( .A(KEYINPUT107), .B(n814), .ZN(n818) );
  AND2_X1 U907 ( .A1(n815), .A2(n818), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n827) );
  INV_X1 U909 ( .A(n818), .ZN(n825) );
  XOR2_X1 U910 ( .A(G1986), .B(G290), .Z(n1001) );
  INV_X1 U911 ( .A(n819), .ZN(n821) );
  NOR2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n975) );
  NAND2_X1 U913 ( .A1(n1001), .A2(n975), .ZN(n823) );
  NAND2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n824) );
  OR2_X1 U915 ( .A1(n825), .A2(n824), .ZN(n826) );
  AND2_X1 U916 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U917 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U918 ( .A(G171), .ZN(G301) );
  NAND2_X1 U919 ( .A1(n829), .A2(G2106), .ZN(n830) );
  XOR2_X1 U920 ( .A(KEYINPUT109), .B(n830), .Z(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U925 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  INV_X1 U927 ( .A(G132), .ZN(G219) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G82), .ZN(G220) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U933 ( .A(G1341), .B(G2454), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n836), .B(G2430), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n837), .B(G1348), .ZN(n843) );
  XOR2_X1 U936 ( .A(G2443), .B(G2427), .Z(n839) );
  XNOR2_X1 U937 ( .A(G2438), .B(G2446), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n841) );
  XOR2_X1 U939 ( .A(G2451), .B(G2435), .Z(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n844), .A2(G14), .ZN(n845) );
  XOR2_X1 U943 ( .A(KEYINPUT108), .B(n845), .Z(G401) );
  XOR2_X1 U944 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2067), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2090), .B(G2072), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U951 ( .A(G2084), .B(G2078), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1991), .B(G1956), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1981), .B(G1966), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U956 ( .A(G1986), .B(G1976), .Z(n857) );
  XNOR2_X1 U957 ( .A(G1961), .B(G1971), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U960 ( .A(KEYINPUT111), .B(G2474), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U962 ( .A(G1996), .B(KEYINPUT41), .Z(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G124), .A2(n883), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT44), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n865), .B(KEYINPUT112), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G112), .A2(n884), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G100), .A2(n887), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G136), .A2(n513), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U972 ( .A1(n871), .A2(n870), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G103), .A2(n887), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G139), .A2(n513), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G127), .A2(n883), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G115), .A2(n884), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n964) );
  XNOR2_X1 U981 ( .A(n879), .B(n964), .ZN(n882) );
  XNOR2_X1 U982 ( .A(G160), .B(n880), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n882), .B(n881), .ZN(n896) );
  NAND2_X1 U984 ( .A1(G130), .A2(n883), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G118), .A2(n884), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U987 ( .A1(G106), .A2(n887), .ZN(n890) );
  NAND2_X1 U988 ( .A1(G142), .A2(n513), .ZN(n889) );
  NAND2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U990 ( .A(KEYINPUT45), .B(n891), .ZN(n892) );
  XNOR2_X1 U991 ( .A(KEYINPUT113), .B(n892), .ZN(n893) );
  NOR2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U993 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U994 ( .A(G164), .B(G162), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n904) );
  XOR2_X1 U996 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n900) );
  XNOR2_X1 U997 ( .A(n971), .B(KEYINPUT48), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(n993), .B(n906), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(G171), .B(n1003), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1005 ( .A(G286), .B(n909), .Z(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G397) );
  OR2_X1 U1007 ( .A1(n916), .A2(G401), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(n916), .ZN(G319) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1016 ( .A(G1971), .B(G22), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(G23), .B(G1976), .ZN(n917) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n920) );
  XOR2_X1 U1019 ( .A(G1986), .B(G24), .Z(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n922) );
  XOR2_X1 U1021 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n921) );
  XNOR2_X1 U1022 ( .A(n922), .B(n921), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G21), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G5), .B(G1961), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n939) );
  XOR2_X1 U1027 ( .A(G1981), .B(G6), .Z(n929) );
  XNOR2_X1 U1028 ( .A(n927), .B(G20), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(G19), .B(G1341), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(KEYINPUT124), .B(n932), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(G1348), .B(KEYINPUT59), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(n933), .B(G4), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1036 ( .A(KEYINPUT60), .B(n936), .Z(n937) );
  XNOR2_X1 U1037 ( .A(KEYINPUT125), .B(n937), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1039 ( .A(KEYINPUT61), .B(n940), .Z(n941) );
  NOR2_X1 U1040 ( .A1(G16), .A2(n941), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(KEYINPUT127), .B(n942), .ZN(n992) );
  XOR2_X1 U1042 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n960) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n955) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n943) );
  NAND2_X1 U1045 ( .A1(n943), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G2072), .B(G33), .ZN(n945) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n944) );
  NOR2_X1 U1048 ( .A1(n945), .A2(n944), .ZN(n950) );
  XOR2_X1 U1049 ( .A(n946), .B(G27), .Z(n948) );
  XNOR2_X1 U1050 ( .A(G2067), .B(G26), .ZN(n947) );
  NOR2_X1 U1051 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1052 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n953), .ZN(n954) );
  NOR2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1056 ( .A(G2084), .B(G34), .Z(n956) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n956), .ZN(n957) );
  NAND2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(n960), .B(n959), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(G29), .A2(n961), .ZN(n962) );
  XOR2_X1 U1061 ( .A(KEYINPUT118), .B(n962), .Z(n963) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n963), .ZN(n990) );
  XOR2_X1 U1063 ( .A(G2072), .B(n964), .Z(n966) );
  XOR2_X1 U1064 ( .A(G164), .B(G2078), .Z(n965) );
  NOR2_X1 U1065 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1066 ( .A(KEYINPUT50), .B(n967), .Z(n983) );
  XOR2_X1 U1067 ( .A(G2084), .B(G160), .Z(n968) );
  NOR2_X1 U1068 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n980) );
  XOR2_X1 U1072 ( .A(G2090), .B(G162), .Z(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(n978), .B(KEYINPUT51), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(KEYINPUT115), .B(n981), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1078 ( .A(n984), .B(KEYINPUT52), .Z(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT116), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(KEYINPUT55), .A2(n986), .ZN(n988) );
  INV_X1 U1081 ( .A(G29), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n1023) );
  XNOR2_X1 U1085 ( .A(G301), .B(G1961), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n993), .B(G1341), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n1017) );
  XOR2_X1 U1088 ( .A(G168), .B(G1966), .Z(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1090 ( .A(KEYINPUT57), .B(n998), .Z(n999) );
  XNOR2_X1 U1091 ( .A(KEYINPUT120), .B(n999), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(n1000), .B(G1956), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G1348), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1015) );
  XOR2_X1 U1097 ( .A(n1008), .B(KEYINPUT121), .Z(n1010) );
  XOR2_X1 U1098 ( .A(G166), .B(G1971), .Z(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT122), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(G16), .B(KEYINPUT119), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT56), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(n1021), .B(KEYINPUT123), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(n1024), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

