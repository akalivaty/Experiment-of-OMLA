

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722;

  AND2_X1 U370 ( .A1(n392), .A2(n634), .ZN(n349) );
  BUF_X1 U371 ( .A(n654), .Z(n350) );
  XNOR2_X1 U372 ( .A(n438), .B(n437), .ZN(n524) );
  XNOR2_X1 U373 ( .A(n479), .B(n414), .ZN(n703) );
  XNOR2_X1 U374 ( .A(n454), .B(n453), .ZN(n690) );
  XOR2_X1 U375 ( .A(KEYINPUT65), .B(G101), .Z(n475) );
  XOR2_X1 U376 ( .A(G104), .B(G107), .Z(n454) );
  INV_X1 U377 ( .A(G953), .ZN(n708) );
  XNOR2_X2 U378 ( .A(n603), .B(n604), .ZN(n605) );
  NAND2_X2 U379 ( .A1(n413), .A2(n591), .ZN(n412) );
  NAND2_X1 U380 ( .A1(n349), .A2(n574), .ZN(n391) );
  NOR2_X2 U381 ( .A1(n402), .A2(n520), .ZN(n401) );
  XNOR2_X2 U382 ( .A(n561), .B(KEYINPUT1), .ZN(n638) );
  NOR2_X1 U383 ( .A1(n567), .A2(n566), .ZN(n568) );
  AND2_X1 U384 ( .A1(n596), .A2(n411), .ZN(n410) );
  NOR2_X1 U385 ( .A1(n717), .A2(n722), .ZN(n569) );
  XNOR2_X1 U386 ( .A(n568), .B(KEYINPUT40), .ZN(n722) );
  XNOR2_X1 U387 ( .A(n690), .B(n404), .ZN(n485) );
  XNOR2_X1 U388 ( .A(n484), .B(n483), .ZN(n691) );
  XNOR2_X1 U389 ( .A(n447), .B(n446), .ZN(n484) );
  XNOR2_X1 U390 ( .A(n473), .B(G134), .ZN(n442) );
  XOR2_X1 U391 ( .A(G122), .B(G116), .Z(n482) );
  XOR2_X1 U392 ( .A(G125), .B(G146), .Z(n479) );
  XNOR2_X2 U393 ( .A(n391), .B(n390), .ZN(n374) );
  XNOR2_X1 U394 ( .A(n704), .B(n353), .ZN(n459) );
  XNOR2_X1 U395 ( .A(G119), .B(KEYINPUT96), .ZN(n446) );
  XOR2_X1 U396 ( .A(G113), .B(KEYINPUT3), .Z(n447) );
  XNOR2_X1 U397 ( .A(n441), .B(n442), .ZN(n704) );
  XNOR2_X1 U398 ( .A(n488), .B(n487), .ZN(n489) );
  INV_X1 U399 ( .A(KEYINPUT84), .ZN(n487) );
  XNOR2_X1 U400 ( .A(n418), .B(G140), .ZN(n414) );
  XOR2_X1 U401 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n418) );
  XNOR2_X1 U402 ( .A(n462), .B(n461), .ZN(n561) );
  XNOR2_X1 U403 ( .A(n460), .B(G469), .ZN(n461) );
  INV_X1 U404 ( .A(KEYINPUT69), .ZN(n460) );
  OR2_X1 U405 ( .A1(G902), .A2(G237), .ZN(n486) );
  INV_X1 U406 ( .A(KEYINPUT48), .ZN(n390) );
  AND2_X1 U407 ( .A1(n721), .A2(KEYINPUT44), .ZN(n505) );
  NOR2_X1 U408 ( .A1(G237), .A2(G953), .ZN(n433) );
  XOR2_X1 U409 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n429) );
  XNOR2_X1 U410 ( .A(G113), .B(G122), .ZN(n431) );
  XOR2_X1 U411 ( .A(G131), .B(G104), .Z(n432) );
  XNOR2_X1 U412 ( .A(n705), .B(KEYINPUT87), .ZN(n394) );
  XOR2_X1 U413 ( .A(KEYINPUT108), .B(n507), .Z(n656) );
  NOR2_X1 U414 ( .A1(n522), .A2(n524), .ZN(n507) );
  NOR2_X1 U415 ( .A1(n640), .A2(n553), .ZN(n376) );
  XNOR2_X1 U416 ( .A(n451), .B(n450), .ZN(n537) );
  NOR2_X1 U417 ( .A1(G902), .A2(n608), .ZN(n450) );
  XNOR2_X1 U418 ( .A(G119), .B(G110), .ZN(n416) );
  XNOR2_X1 U419 ( .A(KEYINPUT23), .B(KEYINPUT100), .ZN(n417) );
  XNOR2_X1 U420 ( .A(n370), .B(n369), .ZN(n368) );
  XNOR2_X1 U421 ( .A(KEYINPUT24), .B(G128), .ZN(n370) );
  XNOR2_X1 U422 ( .A(G137), .B(KEYINPUT99), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n419) );
  XNOR2_X1 U424 ( .A(n366), .B(KEYINPUT66), .ZN(n365) );
  NAND2_X1 U425 ( .A1(n708), .A2(G234), .ZN(n364) );
  INV_X1 U426 ( .A(KEYINPUT8), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n691), .B(n406), .ZN(n405) );
  XNOR2_X1 U428 ( .A(n352), .B(n485), .ZN(n403) );
  XNOR2_X1 U429 ( .A(n480), .B(n476), .ZN(n406) );
  XNOR2_X1 U430 ( .A(n563), .B(n562), .ZN(n651) );
  INV_X1 U431 ( .A(KEYINPUT41), .ZN(n562) );
  NOR2_X1 U432 ( .A1(n657), .A2(n656), .ZN(n563) );
  XNOR2_X1 U433 ( .A(n548), .B(n547), .ZN(n567) );
  XNOR2_X1 U434 ( .A(n546), .B(KEYINPUT39), .ZN(n547) );
  XNOR2_X1 U435 ( .A(KEYINPUT34), .B(KEYINPUT72), .ZN(n499) );
  NAND2_X1 U436 ( .A1(n397), .A2(n396), .ZN(n395) );
  INV_X1 U437 ( .A(n561), .ZN(n396) );
  XNOR2_X1 U438 ( .A(n560), .B(n358), .ZN(n397) );
  XNOR2_X1 U439 ( .A(n470), .B(n469), .ZN(n551) );
  BUF_X1 U440 ( .A(n537), .Z(n647) );
  AND2_X2 U441 ( .A1(n410), .A2(n412), .ZN(n685) );
  XOR2_X1 U442 ( .A(n459), .B(n458), .Z(n683) );
  NAND2_X1 U443 ( .A1(n685), .A2(G210), .ZN(n385) );
  XOR2_X1 U444 ( .A(KEYINPUT4), .B(KEYINPUT81), .Z(n472) );
  XOR2_X1 U445 ( .A(KEYINPUT97), .B(KEYINPUT17), .Z(n476) );
  AND2_X1 U446 ( .A1(n374), .A2(n409), .ZN(n590) );
  NAND2_X1 U447 ( .A1(G237), .A2(G234), .ZN(n493) );
  NOR2_X1 U448 ( .A1(n553), .A2(n552), .ZN(n559) );
  OR2_X1 U449 ( .A1(n551), .A2(n640), .ZN(n552) );
  XNOR2_X1 U450 ( .A(n449), .B(G116), .ZN(n398) );
  NOR2_X1 U451 ( .A1(n636), .A2(n373), .ZN(n372) );
  INV_X1 U452 ( .A(n635), .ZN(n373) );
  XNOR2_X1 U453 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U454 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n481) );
  XNOR2_X1 U455 ( .A(G107), .B(KEYINPUT106), .ZN(n420) );
  XOR2_X1 U456 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n421) );
  XNOR2_X1 U457 ( .A(n351), .B(n434), .ZN(n435) );
  XNOR2_X1 U458 ( .A(G902), .B(KEYINPUT15), .ZN(n463) );
  INV_X1 U459 ( .A(KEYINPUT70), .ZN(n404) );
  NOR2_X1 U460 ( .A1(n638), .A2(n408), .ZN(n407) );
  INV_X1 U461 ( .A(n641), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U463 ( .A(KEYINPUT22), .B(KEYINPUT73), .ZN(n509) );
  AND2_X1 U464 ( .A1(n545), .A2(n377), .ZN(n580) );
  NAND2_X1 U465 ( .A1(n551), .A2(n376), .ZN(n375) );
  BUF_X1 U466 ( .A(n550), .Z(n583) );
  XNOR2_X1 U467 ( .A(n492), .B(n491), .ZN(n399) );
  XNOR2_X1 U468 ( .A(KEYINPUT19), .B(KEYINPUT79), .ZN(n491) );
  INV_X1 U469 ( .A(n647), .ZN(n389) );
  NAND2_X1 U470 ( .A1(n511), .A2(n638), .ZN(n532) );
  XNOR2_X1 U471 ( .A(n415), .B(n703), .ZN(n599) );
  XNOR2_X1 U472 ( .A(n367), .B(n363), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n371), .B(n368), .ZN(n367) );
  INV_X1 U474 ( .A(n395), .ZN(n575) );
  XNOR2_X1 U475 ( .A(n503), .B(KEYINPUT82), .ZN(n504) );
  INV_X1 U476 ( .A(KEYINPUT35), .ZN(n503) );
  NOR2_X1 U477 ( .A1(n395), .A2(n399), .ZN(n625) );
  XNOR2_X1 U478 ( .A(n386), .B(KEYINPUT110), .ZN(n720) );
  NOR2_X1 U479 ( .A1(n532), .A2(n387), .ZN(n386) );
  NAND2_X1 U480 ( .A1(n389), .A2(n388), .ZN(n387) );
  INV_X1 U481 ( .A(n551), .ZN(n388) );
  NOR2_X1 U482 ( .A1(n522), .A2(n521), .ZN(n627) );
  NOR2_X1 U483 ( .A1(n561), .A2(n637), .ZN(n544) );
  XNOR2_X1 U484 ( .A(n683), .B(n360), .ZN(n379) );
  INV_X1 U485 ( .A(KEYINPUT56), .ZN(n381) );
  NAND2_X1 U486 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U487 ( .A(n385), .B(n359), .ZN(n384) );
  XOR2_X1 U488 ( .A(n432), .B(n431), .Z(n351) );
  XOR2_X1 U489 ( .A(n477), .B(n478), .Z(n352) );
  XOR2_X1 U490 ( .A(n475), .B(G146), .Z(n353) );
  INV_X1 U491 ( .A(n636), .ZN(n409) );
  AND2_X1 U492 ( .A1(n394), .A2(n589), .ZN(n355) );
  AND2_X1 U493 ( .A1(n512), .A2(n407), .ZN(n356) );
  XOR2_X1 U494 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n357) );
  XNOR2_X1 U495 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n358) );
  XNOR2_X1 U496 ( .A(n405), .B(n403), .ZN(n679) );
  XNOR2_X1 U497 ( .A(n398), .B(n459), .ZN(n608) );
  XOR2_X1 U498 ( .A(n679), .B(n682), .Z(n359) );
  NOR2_X1 U499 ( .A1(G952), .A2(n708), .ZN(n689) );
  INV_X1 U500 ( .A(n689), .ZN(n383) );
  XNOR2_X1 U501 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n360) );
  XNOR2_X2 U502 ( .A(n362), .B(n504), .ZN(n721) );
  XNOR2_X1 U503 ( .A(n598), .B(n599), .ZN(n600) );
  XNOR2_X1 U504 ( .A(n609), .B(n610), .ZN(n611) );
  XNOR2_X2 U505 ( .A(n361), .B(n357), .ZN(n668) );
  NAND2_X1 U506 ( .A1(n525), .A2(n554), .ZN(n361) );
  NAND2_X1 U507 ( .A1(n695), .A2(n595), .ZN(n596) );
  XNOR2_X2 U508 ( .A(n400), .B(KEYINPUT45), .ZN(n695) );
  NOR2_X2 U509 ( .A1(n501), .A2(n502), .ZN(n362) );
  NAND2_X1 U510 ( .A1(n419), .A2(G221), .ZN(n363) );
  XNOR2_X1 U511 ( .A(n416), .B(n417), .ZN(n371) );
  NAND2_X2 U512 ( .A1(n374), .A2(n372), .ZN(n705) );
  NAND2_X1 U513 ( .A1(n551), .A2(n506), .ZN(n637) );
  NOR2_X1 U514 ( .A1(n561), .A2(n375), .ZN(n377) );
  AND2_X1 U515 ( .A1(n378), .A2(n383), .ZN(G54) );
  XNOR2_X1 U516 ( .A(n380), .B(n379), .ZN(n378) );
  NAND2_X1 U517 ( .A1(n685), .A2(G469), .ZN(n380) );
  NAND2_X1 U518 ( .A1(n355), .A2(n695), .ZN(n413) );
  XNOR2_X1 U519 ( .A(n382), .B(n381), .ZN(G51) );
  NOR2_X1 U520 ( .A1(n720), .A2(n719), .ZN(n516) );
  XNOR2_X1 U521 ( .A(n393), .B(KEYINPUT75), .ZN(n392) );
  NAND2_X1 U522 ( .A1(n588), .A2(n587), .ZN(n393) );
  NOR2_X1 U523 ( .A1(n399), .A2(n497), .ZN(n498) );
  NAND2_X1 U524 ( .A1(n401), .A2(n519), .ZN(n400) );
  NAND2_X1 U525 ( .A1(n518), .A2(n536), .ZN(n402) );
  NAND2_X1 U526 ( .A1(n511), .A2(n356), .ZN(n513) );
  NAND2_X1 U527 ( .A1(n412), .A2(n596), .ZN(n674) );
  INV_X1 U528 ( .A(n597), .ZN(n411) );
  NOR2_X1 U529 ( .A1(n638), .A2(n637), .ZN(n525) );
  BUF_X1 U530 ( .A(n651), .Z(n669) );
  XNOR2_X1 U531 ( .A(n445), .B(n444), .ZN(n448) );
  XNOR2_X1 U532 ( .A(n448), .B(n484), .ZN(n449) );
  INV_X1 U533 ( .A(KEYINPUT88), .ZN(n546) );
  XNOR2_X1 U534 ( .A(KEYINPUT63), .B(KEYINPUT93), .ZN(n612) );
  NAND2_X1 U535 ( .A1(G217), .A2(n419), .ZN(n426) );
  XNOR2_X1 U536 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U537 ( .A(n422), .B(KEYINPUT105), .Z(n424) );
  XNOR2_X2 U538 ( .A(G128), .B(G143), .ZN(n473) );
  XNOR2_X1 U539 ( .A(n482), .B(n442), .ZN(n423) );
  XNOR2_X1 U540 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U541 ( .A(n426), .B(n425), .ZN(n684) );
  NOR2_X1 U542 ( .A1(n684), .A2(G902), .ZN(n427) );
  XNOR2_X1 U543 ( .A(n427), .B(G478), .ZN(n523) );
  INV_X1 U544 ( .A(n523), .ZN(n522) );
  XNOR2_X1 U545 ( .A(G143), .B(KEYINPUT104), .ZN(n428) );
  XNOR2_X1 U546 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U547 ( .A(n703), .B(n430), .Z(n436) );
  XNOR2_X1 U548 ( .A(n433), .B(KEYINPUT78), .ZN(n443) );
  NAND2_X1 U549 ( .A1(G214), .A2(n443), .ZN(n434) );
  XNOR2_X1 U550 ( .A(n436), .B(n435), .ZN(n602) );
  NOR2_X1 U551 ( .A1(G902), .A2(n602), .ZN(n438) );
  XNOR2_X1 U552 ( .A(KEYINPUT13), .B(G475), .ZN(n437) );
  NAND2_X1 U553 ( .A1(n522), .A2(n524), .ZN(n581) );
  XOR2_X1 U554 ( .A(n581), .B(KEYINPUT83), .Z(n502) );
  INV_X1 U555 ( .A(G472), .ZN(n451) );
  XOR2_X1 U556 ( .A(G131), .B(KEYINPUT68), .Z(n440) );
  XNOR2_X1 U557 ( .A(G137), .B(KEYINPUT4), .ZN(n439) );
  XNOR2_X1 U558 ( .A(n440), .B(n439), .ZN(n441) );
  NAND2_X1 U559 ( .A1(n443), .A2(G210), .ZN(n445) );
  XOR2_X1 U560 ( .A(KEYINPUT5), .B(KEYINPUT102), .Z(n444) );
  XNOR2_X1 U561 ( .A(KEYINPUT6), .B(KEYINPUT107), .ZN(n452) );
  XNOR2_X1 U562 ( .A(n537), .B(n452), .ZN(n554) );
  XNOR2_X1 U563 ( .A(G110), .B(KEYINPUT95), .ZN(n453) );
  XOR2_X1 U564 ( .A(G140), .B(KEYINPUT80), .Z(n456) );
  NAND2_X1 U565 ( .A1(G227), .A2(n708), .ZN(n455) );
  XNOR2_X1 U566 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U567 ( .A(n485), .B(n457), .ZN(n458) );
  NOR2_X1 U568 ( .A1(G902), .A2(n683), .ZN(n462) );
  XNOR2_X1 U569 ( .A(n463), .B(KEYINPUT94), .ZN(n597) );
  NAND2_X1 U570 ( .A1(G234), .A2(n597), .ZN(n464) );
  XNOR2_X1 U571 ( .A(KEYINPUT20), .B(n464), .ZN(n466) );
  NAND2_X1 U572 ( .A1(n466), .A2(G221), .ZN(n465) );
  XOR2_X1 U573 ( .A(KEYINPUT21), .B(n465), .Z(n506) );
  NOR2_X1 U574 ( .A1(G902), .A2(n599), .ZN(n470) );
  XOR2_X1 U575 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n468) );
  NAND2_X1 U576 ( .A1(n466), .A2(G217), .ZN(n467) );
  XNOR2_X1 U577 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U578 ( .A1(G214), .A2(n486), .ZN(n653) );
  NAND2_X1 U579 ( .A1(G224), .A2(n708), .ZN(n471) );
  XNOR2_X1 U580 ( .A(n472), .B(n471), .ZN(n478) );
  INV_X1 U581 ( .A(n473), .ZN(n474) );
  XNOR2_X1 U582 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X1 U583 ( .A(n479), .B(KEYINPUT18), .ZN(n480) );
  NAND2_X1 U584 ( .A1(n679), .A2(n597), .ZN(n490) );
  NAND2_X1 U585 ( .A1(n486), .A2(G210), .ZN(n488) );
  XNOR2_X2 U586 ( .A(n490), .B(n489), .ZN(n550) );
  NAND2_X1 U587 ( .A1(n653), .A2(n550), .ZN(n492) );
  XOR2_X1 U588 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n494) );
  XNOR2_X1 U589 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U590 ( .A1(G952), .A2(n495), .ZN(n667) );
  NOR2_X1 U591 ( .A1(G953), .A2(n667), .ZN(n543) );
  NAND2_X1 U592 ( .A1(G902), .A2(n495), .ZN(n540) );
  OR2_X1 U593 ( .A1(n708), .A2(G898), .ZN(n694) );
  NOR2_X1 U594 ( .A1(n540), .A2(n694), .ZN(n496) );
  NOR2_X1 U595 ( .A1(n543), .A2(n496), .ZN(n497) );
  XNOR2_X1 U596 ( .A(n498), .B(KEYINPUT0), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n527), .B(KEYINPUT98), .ZN(n529) );
  NAND2_X1 U598 ( .A1(n668), .A2(n529), .ZN(n500) );
  XNOR2_X1 U599 ( .A(n500), .B(n499), .ZN(n501) );
  NOR2_X1 U600 ( .A1(KEYINPUT90), .A2(n505), .ZN(n520) );
  NAND2_X1 U601 ( .A1(KEYINPUT90), .A2(n721), .ZN(n514) );
  INV_X1 U602 ( .A(n506), .ZN(n640) );
  NOR2_X1 U603 ( .A1(n640), .A2(n656), .ZN(n508) );
  NAND2_X1 U604 ( .A1(n527), .A2(n508), .ZN(n510) );
  INV_X1 U605 ( .A(n554), .ZN(n512) );
  XNOR2_X1 U606 ( .A(KEYINPUT109), .B(n551), .ZN(n641) );
  XOR2_X1 U607 ( .A(KEYINPUT32), .B(n513), .Z(n719) );
  NAND2_X1 U608 ( .A1(n514), .A2(n516), .ZN(n515) );
  NAND2_X1 U609 ( .A1(n515), .A2(KEYINPUT44), .ZN(n519) );
  NOR2_X1 U610 ( .A1(KEYINPUT44), .A2(n721), .ZN(n517) );
  NAND2_X1 U611 ( .A1(n517), .A2(n516), .ZN(n518) );
  INV_X1 U612 ( .A(n524), .ZN(n521) );
  INV_X1 U613 ( .A(n627), .ZN(n566) );
  NOR2_X1 U614 ( .A1(n524), .A2(n523), .ZN(n629) );
  INV_X1 U615 ( .A(n629), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n566), .A2(n549), .ZN(n576) );
  INV_X1 U617 ( .A(n576), .ZN(n658) );
  NAND2_X1 U618 ( .A1(n525), .A2(n647), .ZN(n526) );
  XNOR2_X1 U619 ( .A(n526), .B(KEYINPUT103), .ZN(n649) );
  NAND2_X1 U620 ( .A1(n649), .A2(n527), .ZN(n528) );
  XNOR2_X1 U621 ( .A(KEYINPUT31), .B(n528), .ZN(n630) );
  NAND2_X1 U622 ( .A1(n544), .A2(n529), .ZN(n530) );
  NOR2_X1 U623 ( .A1(n647), .A2(n530), .ZN(n617) );
  NOR2_X1 U624 ( .A1(n630), .A2(n617), .ZN(n531) );
  NOR2_X1 U625 ( .A1(n658), .A2(n531), .ZN(n535) );
  NOR2_X1 U626 ( .A1(n554), .A2(n532), .ZN(n533) );
  XNOR2_X1 U627 ( .A(n533), .B(KEYINPUT89), .ZN(n534) );
  NOR2_X1 U628 ( .A1(n641), .A2(n534), .ZN(n614) );
  NOR2_X1 U629 ( .A1(n535), .A2(n614), .ZN(n536) );
  XOR2_X1 U630 ( .A(n550), .B(KEYINPUT38), .Z(n654) );
  INV_X1 U631 ( .A(KEYINPUT30), .ZN(n539) );
  NAND2_X1 U632 ( .A1(n537), .A2(n653), .ZN(n538) );
  XNOR2_X1 U633 ( .A(n539), .B(n538), .ZN(n545) );
  OR2_X1 U634 ( .A1(n708), .A2(n540), .ZN(n541) );
  NOR2_X1 U635 ( .A1(G900), .A2(n541), .ZN(n542) );
  NOR2_X1 U636 ( .A1(n543), .A2(n542), .ZN(n553) );
  NAND2_X1 U637 ( .A1(n350), .A2(n580), .ZN(n548) );
  OR2_X1 U638 ( .A1(n549), .A2(n567), .ZN(n635) );
  NAND2_X1 U639 ( .A1(n554), .A2(n559), .ZN(n556) );
  NAND2_X1 U640 ( .A1(n627), .A2(n653), .ZN(n555) );
  NOR2_X1 U641 ( .A1(n556), .A2(n555), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n638), .A2(n570), .ZN(n557) );
  XOR2_X1 U643 ( .A(KEYINPUT43), .B(n557), .Z(n558) );
  NOR2_X1 U644 ( .A1(n583), .A2(n558), .ZN(n636) );
  XOR2_X1 U645 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n565) );
  NAND2_X1 U646 ( .A1(n559), .A2(n647), .ZN(n560) );
  NAND2_X1 U647 ( .A1(n653), .A2(n654), .ZN(n657) );
  NAND2_X1 U648 ( .A1(n575), .A2(n651), .ZN(n564) );
  XNOR2_X1 U649 ( .A(n565), .B(n564), .ZN(n717) );
  XNOR2_X1 U650 ( .A(n569), .B(KEYINPUT46), .ZN(n574) );
  NAND2_X1 U651 ( .A1(n570), .A2(n583), .ZN(n571) );
  XOR2_X1 U652 ( .A(KEYINPUT36), .B(n571), .Z(n573) );
  INV_X1 U653 ( .A(n638), .ZN(n572) );
  NAND2_X1 U654 ( .A1(n573), .A2(n572), .ZN(n634) );
  INV_X1 U655 ( .A(KEYINPUT76), .ZN(n579) );
  NOR2_X1 U656 ( .A1(n579), .A2(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U657 ( .A1(n625), .A2(n576), .ZN(n577) );
  XNOR2_X1 U658 ( .A(n578), .B(n577), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n579), .A2(KEYINPUT47), .ZN(n586) );
  INV_X1 U660 ( .A(n580), .ZN(n582) );
  NOR2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n624) );
  XNOR2_X1 U663 ( .A(KEYINPUT86), .B(n624), .ZN(n585) );
  AND2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U665 ( .A1(KEYINPUT85), .A2(n590), .ZN(n589) );
  INV_X1 U666 ( .A(KEYINPUT2), .ZN(n591) );
  INV_X1 U667 ( .A(n590), .ZN(n594) );
  XOR2_X1 U668 ( .A(n635), .B(KEYINPUT85), .Z(n592) );
  NAND2_X1 U669 ( .A1(n592), .A2(KEYINPUT2), .ZN(n593) );
  NOR2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U671 ( .A1(G217), .A2(n685), .ZN(n598) );
  NOR2_X2 U672 ( .A1(n600), .A2(n689), .ZN(n601) );
  XNOR2_X1 U673 ( .A(n601), .B(KEYINPUT122), .ZN(G66) );
  XOR2_X1 U674 ( .A(n602), .B(KEYINPUT59), .Z(n604) );
  NAND2_X1 U675 ( .A1(n685), .A2(G475), .ZN(n603) );
  NOR2_X2 U676 ( .A1(n605), .A2(n689), .ZN(n607) );
  XNOR2_X1 U677 ( .A(KEYINPUT60), .B(KEYINPUT64), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n607), .B(n606), .ZN(G60) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT62), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G472), .A2(n685), .ZN(n609) );
  NOR2_X2 U681 ( .A1(n611), .A2(n689), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n613), .B(n612), .ZN(G57) );
  XOR2_X1 U683 ( .A(G101), .B(n614), .Z(G3) );
  XOR2_X1 U684 ( .A(G104), .B(KEYINPUT113), .Z(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n627), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n616), .B(n615), .ZN(G6) );
  XNOR2_X1 U687 ( .A(G107), .B(KEYINPUT27), .ZN(n621) );
  XOR2_X1 U688 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n619) );
  NAND2_X1 U689 ( .A1(n617), .A2(n629), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n621), .B(n620), .ZN(G9) );
  XOR2_X1 U692 ( .A(G128), .B(KEYINPUT29), .Z(n623) );
  NAND2_X1 U693 ( .A1(n625), .A2(n629), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n623), .B(n622), .ZN(G30) );
  XNOR2_X1 U695 ( .A(G143), .B(n624), .ZN(G45) );
  NAND2_X1 U696 ( .A1(n625), .A2(n627), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n626), .B(G146), .ZN(G48) );
  NAND2_X1 U698 ( .A1(n630), .A2(n627), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(G113), .ZN(G15) );
  XOR2_X1 U700 ( .A(G116), .B(KEYINPUT115), .Z(n632) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U702 ( .A(n632), .B(n631), .ZN(G18) );
  XOR2_X1 U703 ( .A(G125), .B(KEYINPUT37), .Z(n633) );
  XNOR2_X1 U704 ( .A(n634), .B(n633), .ZN(G27) );
  XNOR2_X1 U705 ( .A(G134), .B(n635), .ZN(G36) );
  XOR2_X1 U706 ( .A(G140), .B(n636), .Z(G42) );
  NAND2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U708 ( .A(KEYINPUT50), .B(n639), .ZN(n645) );
  XOR2_X1 U709 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n643) );
  NAND2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U712 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U714 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U715 ( .A(n650), .B(KEYINPUT51), .ZN(n652) );
  NAND2_X1 U716 ( .A1(n652), .A2(n669), .ZN(n664) );
  NOR2_X1 U717 ( .A1(n350), .A2(n653), .ZN(n655) );
  NOR2_X1 U718 ( .A1(n656), .A2(n655), .ZN(n660) );
  NOR2_X1 U719 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U720 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U721 ( .A(KEYINPUT117), .B(n661), .ZN(n662) );
  NAND2_X1 U722 ( .A1(n662), .A2(n668), .ZN(n663) );
  NAND2_X1 U723 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U724 ( .A(KEYINPUT52), .B(n665), .Z(n666) );
  NOR2_X1 U725 ( .A1(n667), .A2(n666), .ZN(n672) );
  NAND2_X1 U726 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U727 ( .A(KEYINPUT118), .B(n670), .Z(n671) );
  NOR2_X1 U728 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U729 ( .A(KEYINPUT119), .B(n673), .Z(n675) );
  NAND2_X1 U730 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U731 ( .A(KEYINPUT120), .B(n676), .ZN(n677) );
  NOR2_X1 U732 ( .A1(n677), .A2(G953), .ZN(n678) );
  XNOR2_X1 U733 ( .A(n678), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U734 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n681) );
  XNOR2_X1 U735 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n680) );
  XNOR2_X1 U736 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U737 ( .A(n684), .B(KEYINPUT121), .Z(n687) );
  NAND2_X1 U738 ( .A1(n685), .A2(G478), .ZN(n686) );
  XNOR2_X1 U739 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U740 ( .A1(n689), .A2(n688), .ZN(G63) );
  XNOR2_X1 U741 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U742 ( .A(n692), .B(G101), .ZN(n693) );
  NAND2_X1 U743 ( .A1(n694), .A2(n693), .ZN(n702) );
  NAND2_X1 U744 ( .A1(n708), .A2(n695), .ZN(n699) );
  NAND2_X1 U745 ( .A1(G953), .A2(G224), .ZN(n696) );
  XNOR2_X1 U746 ( .A(KEYINPUT61), .B(n696), .ZN(n697) );
  NAND2_X1 U747 ( .A1(n697), .A2(G898), .ZN(n698) );
  NAND2_X1 U748 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U749 ( .A(n700), .B(KEYINPUT123), .ZN(n701) );
  XNOR2_X1 U750 ( .A(n702), .B(n701), .ZN(G69) );
  XOR2_X1 U751 ( .A(n704), .B(n703), .Z(n710) );
  XOR2_X1 U752 ( .A(KEYINPUT87), .B(KEYINPUT124), .Z(n706) );
  XNOR2_X1 U753 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U754 ( .A(n710), .B(n707), .ZN(n709) );
  NAND2_X1 U755 ( .A1(n709), .A2(n708), .ZN(n715) );
  XNOR2_X1 U756 ( .A(G227), .B(n710), .ZN(n711) );
  NAND2_X1 U757 ( .A1(n711), .A2(G900), .ZN(n712) );
  NAND2_X1 U758 ( .A1(G953), .A2(n712), .ZN(n713) );
  XOR2_X1 U759 ( .A(KEYINPUT125), .B(n713), .Z(n714) );
  NAND2_X1 U760 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U761 ( .A(KEYINPUT126), .B(n716), .ZN(G72) );
  XNOR2_X1 U762 ( .A(n717), .B(G137), .ZN(n718) );
  XNOR2_X1 U763 ( .A(n718), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U764 ( .A(G119), .B(n719), .Z(G21) );
  XOR2_X1 U765 ( .A(G110), .B(n720), .Z(G12) );
  XOR2_X1 U766 ( .A(n721), .B(G122), .Z(G24) );
  XOR2_X1 U767 ( .A(n722), .B(G131), .Z(G33) );
endmodule

