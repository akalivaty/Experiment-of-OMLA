//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  INV_X1    g000(.A(G64gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(G57gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(G57gat), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n203), .A2(new_n204), .B1(new_n207), .B2(KEYINPUT9), .ZN(new_n208));
  XNOR2_X1  g007(.A(G71gat), .B(G78gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G231gat), .A2(G233gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G127gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n218), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G8gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n212), .B2(new_n211), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n217), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(G183gat), .B(G211gat), .Z(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n225), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G120gat), .B(G148gat), .Z(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT103), .ZN(new_n233));
  XNOR2_X1  g032(.A(G176gat), .B(G204gat), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n233), .B(new_n234), .Z(new_n235));
  XOR2_X1   g034(.A(G99gat), .B(G106gat), .Z(new_n236));
  INV_X1    g035(.A(G85gat), .ZN(new_n237));
  INV_X1    g036(.A(G92gat), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT7), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT7), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(G85gat), .A3(G92gat), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n236), .A2(KEYINPUT98), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT97), .B(G92gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(G99gat), .A2(G106gat), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n243), .A2(new_n237), .B1(KEYINPUT8), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n236), .A2(KEYINPUT98), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n246), .A2(new_n247), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n210), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n246), .A2(new_n247), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n247), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n211), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT10), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT100), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT100), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n250), .A2(new_n253), .A3(new_n257), .A4(new_n254), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n250), .A2(new_n254), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n235), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n250), .A2(new_n253), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(new_n262), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT101), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT101), .B1(new_n264), .B2(new_n262), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT102), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT102), .B1(new_n267), .B2(new_n268), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n263), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n262), .B(KEYINPUT104), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n259), .B1(new_n255), .B2(KEYINPUT100), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n274), .B1(new_n275), .B2(new_n258), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n235), .B1(new_n269), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n251), .A2(new_n252), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT99), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT15), .ZN(new_n282));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(KEYINPUT91), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(KEYINPUT91), .B2(new_n283), .ZN(new_n285));
  NAND2_X1  g084(.A1(G29gat), .A2(G36gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT92), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n289));
  NOR3_X1   g088(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n290), .B(KEYINPUT93), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n289), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n283), .A2(KEYINPUT15), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(new_n288), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n285), .A3(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(KEYINPUT94), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(KEYINPUT94), .ZN(new_n300));
  AOI211_X1 g099(.A(KEYINPUT17), .B(new_n293), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT17), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n298), .B(KEYINPUT94), .ZN(new_n303));
  INV_X1    g102(.A(new_n293), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n281), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G190gat), .B(G218gat), .Z(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n293), .B1(new_n299), .B2(new_n300), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G232gat), .A2(G233gat), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n310), .A2(new_n280), .B1(KEYINPUT41), .B2(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n306), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n308), .B1(new_n306), .B2(new_n312), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n311), .A2(KEYINPUT41), .ZN(new_n315));
  XNOR2_X1  g114(.A(G134gat), .B(G162gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OR3_X1    g117(.A1(new_n313), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n313), .B2(new_n314), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n231), .A2(new_n279), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT105), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n231), .A2(new_n279), .A3(new_n321), .A4(KEYINPUT105), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT90), .ZN(new_n327));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT26), .ZN(new_n330));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT26), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n331), .C1(new_n334), .C2(new_n329), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT27), .B(G183gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT67), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT67), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(G183gat), .ZN(new_n340));
  INV_X1    g139(.A(G183gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(KEYINPUT27), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n338), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(G190gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n337), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n336), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(new_n344), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n335), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT24), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n341), .A2(new_n347), .ZN(new_n354));
  NAND3_X1  g153(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n329), .A2(KEYINPUT23), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT64), .ZN(new_n358));
  OAI22_X1  g157(.A1(new_n358), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT64), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n357), .B(new_n332), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n356), .B1(new_n362), .B2(KEYINPUT65), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n364));
  INV_X1    g163(.A(new_n332), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(KEYINPUT23), .B2(new_n329), .ZN(new_n366));
  INV_X1    g165(.A(new_n329), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n360), .A2(KEYINPUT64), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n364), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n351), .B1(new_n363), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n362), .A2(new_n351), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n353), .A2(KEYINPUT66), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n353), .A2(KEYINPUT66), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(new_n354), .A3(new_n355), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n350), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n328), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n380));
  XNOR2_X1  g179(.A(G211gat), .B(G218gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT75), .ZN(new_n382));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT22), .ZN(new_n384));
  INV_X1    g183(.A(G211gat), .ZN(new_n385));
  INV_X1    g184(.A(G218gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n387), .B(new_n383), .C1(new_n381), .C2(KEYINPUT75), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n377), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT68), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT28), .B1(new_n336), .B2(new_n347), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n341), .A2(KEYINPUT27), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n339), .A2(G183gat), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT67), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT67), .B1(new_n395), .B2(new_n396), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n394), .B1(new_n399), .B2(new_n345), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n393), .B1(new_n400), .B2(new_n335), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n350), .A2(KEYINPUT68), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n392), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n328), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT78), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n406), .B(new_n328), .C1(new_n378), .C2(KEYINPUT29), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n380), .A2(new_n391), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n403), .A2(new_n328), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n378), .A2(new_n404), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n389), .A2(KEYINPUT76), .A3(new_n390), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT76), .B1(new_n389), .B2(new_n390), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n411), .B(new_n412), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT89), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n419));
  INV_X1    g218(.A(new_n417), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n408), .A2(new_n415), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n416), .B2(KEYINPUT37), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n327), .B1(new_n427), .B2(KEYINPUT38), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n425), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT38), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n411), .A2(new_n412), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n413), .A2(new_n414), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n380), .A2(new_n405), .A3(new_n407), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(new_n391), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n432), .B1(new_n437), .B2(KEYINPUT37), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G141gat), .ZN(new_n440));
  INV_X1    g239(.A(G148gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G141gat), .A2(G148gat), .ZN(new_n443));
  AND2_X1   g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(G155gat), .A2(G162gat), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n442), .B(new_n443), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(KEYINPUT80), .A2(G155gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(KEYINPUT80), .A2(G155gat), .ZN(new_n449));
  OAI21_X1  g248(.A(G162gat), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n446), .B1(new_n450), .B2(KEYINPUT2), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT79), .B1(new_n444), .B2(new_n445), .ZN(new_n452));
  INV_X1    g251(.A(G162gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n227), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT79), .ZN(new_n455));
  NAND2_X1  g254(.A1(G155gat), .A2(G162gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(G141gat), .A2(G148gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(G141gat), .A2(G148gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(KEYINPUT2), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n452), .A2(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT81), .B1(new_n451), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n452), .A2(new_n457), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n461), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n454), .A2(new_n456), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n227), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n453), .B1(new_n469), .B2(new_n447), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT2), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n460), .B(new_n467), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n466), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT70), .ZN(new_n475));
  AND2_X1   g274(.A1(G113gat), .A2(G120gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(G113gat), .A2(G120gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G113gat), .ZN(new_n479));
  INV_X1    g278(.A(G120gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G113gat), .A2(G120gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(KEYINPUT70), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G127gat), .B(G134gat), .ZN(new_n484));
  AND2_X1   g283(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n485));
  NOR2_X1   g284(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n478), .A2(new_n483), .A3(new_n484), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n216), .A2(G134gat), .ZN(new_n489));
  INV_X1    g288(.A(G134gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G127gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n491), .A3(KEYINPUT69), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT1), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n481), .A2(new_n493), .A3(new_n482), .ZN(new_n494));
  OR3_X1    g293(.A1(new_n490), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n463), .A2(new_n474), .A3(KEYINPUT4), .A4(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT3), .B1(new_n451), .B2(new_n462), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n488), .A2(new_n496), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT3), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n466), .A2(new_n472), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n466), .A2(new_n472), .A3(new_n496), .A4(new_n488), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n498), .A2(new_n503), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n500), .B1(new_n462), .B2(new_n451), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT82), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n505), .ZN(new_n511));
  INV_X1    g310(.A(new_n504), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n466), .A2(new_n472), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(KEYINPUT82), .A3(new_n500), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n508), .A2(new_n515), .A3(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT83), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT83), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n508), .A2(new_n515), .A3(new_n518), .A4(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n463), .A2(new_n474), .A3(new_n506), .A4(new_n497), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n503), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n526), .A2(KEYINPUT5), .A3(new_n512), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G1gat), .B(G29gat), .Z(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G57gat), .B(G85gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(KEYINPUT6), .A3(new_n535), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n517), .A2(new_n519), .B1(new_n525), .B2(new_n527), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT6), .B1(new_n537), .B2(new_n534), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n529), .A2(new_n535), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n408), .A2(new_n415), .A3(new_n425), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n439), .A2(new_n536), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI211_X1 g342(.A(KEYINPUT90), .B(new_n431), .C1(new_n422), .C2(new_n426), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n429), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n388), .A2(new_n381), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n409), .B1(new_n388), .B2(new_n381), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT3), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(new_n463), .B2(new_n474), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n391), .B1(new_n502), .B2(new_n410), .ZN(new_n551));
  INV_X1    g350(.A(G228gat), .ZN(new_n552));
  INV_X1    g351(.A(G233gat), .ZN(new_n553));
  OAI22_X1  g352(.A1(new_n550), .A2(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT29), .B1(new_n389), .B2(new_n390), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n513), .B1(new_n556), .B2(KEYINPUT3), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n502), .A2(new_n410), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n555), .B(new_n557), .C1(new_n558), .C2(new_n434), .ZN(new_n559));
  INV_X1    g358(.A(G22gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n554), .B2(new_n559), .ZN(new_n563));
  OAI21_X1  g362(.A(G78gat), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(new_n206), .A3(new_n561), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G50gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT87), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G106gat), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n564), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n564), .B2(new_n566), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n525), .A2(new_n503), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n512), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n511), .A2(new_n514), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n504), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(KEYINPUT39), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT39), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n578), .A3(new_n512), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n534), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT40), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n577), .A2(KEYINPUT40), .A3(new_n534), .A4(new_n579), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n539), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n416), .A2(new_n430), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(KEYINPUT30), .A3(new_n541), .ZN(new_n586));
  OR3_X1    g385(.A1(new_n416), .A2(KEYINPUT30), .A3(new_n430), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n572), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n546), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n392), .A2(new_n401), .A3(new_n497), .A4(new_n402), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT72), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n346), .A2(new_n349), .ZN(new_n595));
  INV_X1    g394(.A(new_n335), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT68), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI211_X1 g396(.A(new_n393), .B(new_n335), .C1(new_n346), .C2(new_n349), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n599), .A2(KEYINPUT72), .A3(new_n497), .A4(new_n392), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n403), .A2(new_n500), .ZN(new_n601));
  NAND2_X1  g400(.A1(G227gat), .A2(G233gat), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n594), .A2(new_n600), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT32), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n600), .A3(new_n601), .ZN(new_n610));
  INV_X1    g409(.A(new_n602), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT33), .B1(new_n610), .B2(new_n611), .ZN(new_n613));
  XOR2_X1   g412(.A(G15gat), .B(G43gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT73), .ZN(new_n615));
  XOR2_X1   g414(.A(G71gat), .B(G99gat), .Z(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n612), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  AOI221_X4 g418(.A(new_n609), .B1(KEYINPUT33), .B2(new_n617), .C1(new_n610), .C2(new_n611), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n608), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n610), .A2(new_n611), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n618), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n612), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n620), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n607), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n621), .A2(KEYINPUT36), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT36), .B1(new_n621), .B2(new_n628), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n540), .A2(new_n536), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n632), .A2(KEYINPUT86), .A3(new_n588), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT86), .B1(new_n632), .B2(new_n588), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n572), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n631), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n572), .A2(new_n621), .A3(new_n628), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n633), .B2(new_n634), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT35), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n540), .A2(new_n536), .ZN(new_n641));
  INV_X1    g440(.A(new_n588), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT35), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n638), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n591), .A2(new_n637), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n223), .B1(new_n301), .B2(new_n305), .ZN(new_n646));
  NAND2_X1  g445(.A1(G229gat), .A2(G233gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n310), .A2(new_n222), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT18), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n310), .B2(new_n222), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n309), .A2(KEYINPUT95), .A3(new_n223), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n648), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n647), .B(KEYINPUT13), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n646), .A2(KEYINPUT18), .A3(new_n647), .A4(new_n648), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n651), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G113gat), .B(G141gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G197gat), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT11), .B(G169gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT12), .Z(new_n664));
  NAND2_X1  g463(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n651), .A2(new_n657), .A3(new_n666), .A4(new_n658), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT96), .B1(new_n645), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n640), .A2(new_n644), .ZN(new_n671));
  INV_X1    g470(.A(new_n634), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n632), .A2(KEYINPUT86), .A3(new_n588), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n636), .A3(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n629), .A2(new_n630), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n428), .A2(new_n542), .A3(new_n544), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n674), .B(new_n675), .C1(new_n676), .C2(new_n589), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT96), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n679), .A3(new_n668), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n326), .B1(new_n670), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n641), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n642), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(G8gat), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n684), .A2(KEYINPUT106), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n687), .B2(new_n692), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n688), .A2(new_n689), .B1(new_n686), .B2(new_n693), .ZN(G1325gat));
  AND2_X1   g493(.A1(new_n621), .A2(new_n628), .ZN(new_n695));
  AOI21_X1  g494(.A(G15gat), .B1(new_n681), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n631), .A2(G15gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT107), .Z(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n681), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n636), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n645), .B2(new_n321), .ZN(new_n704));
  INV_X1    g503(.A(new_n321), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n674), .A2(new_n675), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n428), .A2(new_n542), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n589), .B1(new_n707), .B2(new_n545), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n639), .A2(KEYINPUT35), .B1(new_n638), .B2(new_n643), .ZN(new_n710));
  OAI211_X1 g509(.A(KEYINPUT44), .B(new_n705), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n231), .A2(new_n278), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n668), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(new_n641), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT108), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n712), .A2(new_n718), .A3(new_n641), .A4(new_n715), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(G29gat), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n713), .A2(new_n705), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n670), .B2(new_n680), .ZN(new_n722));
  INV_X1    g521(.A(G29gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(new_n723), .A3(new_n641), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n720), .A2(new_n726), .A3(new_n727), .ZN(G1328gat));
  INV_X1    g527(.A(G36gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n722), .A2(new_n729), .A3(new_n642), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n730), .A2(KEYINPUT46), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(KEYINPUT46), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n704), .A2(new_n711), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n733), .A2(new_n588), .A3(new_n714), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n731), .B(new_n732), .C1(new_n729), .C2(new_n734), .ZN(G1329gat));
  INV_X1    g534(.A(G43gat), .ZN(new_n736));
  NOR4_X1   g535(.A1(new_n733), .A2(new_n736), .A3(new_n675), .A4(new_n714), .ZN(new_n737));
  AOI21_X1  g536(.A(G43gat), .B1(new_n722), .B2(new_n695), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT47), .B1(new_n737), .B2(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1330gat));
  INV_X1    g542(.A(G50gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n722), .A2(new_n744), .A3(new_n636), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n704), .A2(new_n636), .A3(new_n711), .A4(new_n715), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G50gat), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1331gat));
  INV_X1    g549(.A(new_n231), .ZN(new_n751));
  NOR4_X1   g550(.A1(new_n751), .A2(new_n705), .A3(new_n668), .A4(new_n279), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n678), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n632), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n588), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  AND2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n756), .B2(new_n757), .ZN(G1333gat));
  OAI21_X1  g559(.A(G71gat), .B1(new_n753), .B2(new_n675), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n695), .A2(new_n205), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n753), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g563(.A1(new_n753), .A2(new_n572), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(new_n206), .ZN(G1335gat));
  AOI21_X1  g565(.A(new_n321), .B1(new_n671), .B2(new_n677), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n231), .A2(new_n668), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(KEYINPUT51), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n641), .A2(new_n278), .A3(new_n237), .ZN(new_n775));
  INV_X1    g574(.A(new_n768), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n279), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n733), .A2(new_n632), .A3(new_n778), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n774), .A2(new_n775), .B1(new_n779), .B2(new_n237), .ZN(G1336gat));
  NOR3_X1   g579(.A1(new_n279), .A2(G92gat), .A3(new_n588), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n771), .B2(new_n772), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n704), .A2(new_n642), .A3(new_n711), .A4(new_n777), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n243), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n785), .A2(new_n786), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n784), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n785), .A2(new_n792), .A3(new_n788), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n785), .B2(new_n788), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n793), .A2(new_n794), .A3(new_n783), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(G1337gat));
  INV_X1    g596(.A(G99gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n695), .A2(new_n798), .A3(new_n278), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n733), .A2(new_n675), .A3(new_n778), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n774), .A2(new_n799), .B1(new_n800), .B2(new_n798), .ZN(G1338gat));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n279), .A2(G106gat), .A3(new_n572), .ZN(new_n803));
  INV_X1    g602(.A(new_n772), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT51), .B1(new_n767), .B2(new_n768), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n802), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n704), .A2(new_n636), .A3(new_n711), .A4(new_n777), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G106gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n802), .B1(new_n773), .B2(new_n803), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT53), .B1(new_n773), .B2(new_n803), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n807), .A2(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n807), .A2(KEYINPUT112), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n816), .ZN(G1339gat));
  NAND2_X1  g616(.A1(new_n261), .A2(new_n262), .ZN(new_n818));
  INV_X1    g617(.A(new_n274), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n818), .B(KEYINPUT54), .C1(new_n819), .C2(new_n261), .ZN(new_n820));
  INV_X1    g619(.A(new_n235), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n276), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(new_n823), .A3(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n273), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT113), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n273), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n820), .A2(new_n823), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n826), .A2(new_n668), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n655), .A2(new_n656), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n647), .B1(new_n646), .B2(new_n648), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n663), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n278), .A2(new_n667), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n705), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  AND4_X1   g636(.A1(new_n667), .A2(new_n319), .A3(new_n320), .A4(new_n835), .ZN(new_n838));
  AND4_X1   g637(.A1(new_n828), .A2(new_n838), .A3(new_n826), .A4(new_n831), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n751), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n322), .A2(new_n668), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n636), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n842), .A2(new_n641), .A3(new_n588), .A4(new_n695), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(new_n479), .A3(new_n669), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n632), .B1(new_n840), .B2(new_n841), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n638), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n588), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n668), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n844), .B1(new_n848), .B2(new_n479), .ZN(G1340gat));
  NAND4_X1  g648(.A1(new_n846), .A2(new_n480), .A3(new_n588), .A4(new_n278), .ZN(new_n850));
  OAI21_X1  g649(.A(G120gat), .B1(new_n843), .B2(new_n279), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(G1341gat));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n216), .A3(new_n231), .ZN(new_n855));
  OAI21_X1  g654(.A(G127gat), .B1(new_n843), .B2(new_n751), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  NAND4_X1  g656(.A1(new_n846), .A2(new_n490), .A3(new_n588), .A4(new_n705), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n843), .B2(new_n321), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(G1343gat));
  NOR3_X1   g661(.A1(new_n631), .A2(new_n632), .A3(new_n642), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n840), .A2(new_n841), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n636), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  INV_X1    g667(.A(new_n825), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n830), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n829), .A2(KEYINPUT116), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n869), .B(new_n668), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n705), .B1(new_n873), .B2(new_n836), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n751), .B1(new_n874), .B2(new_n839), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n868), .B(new_n572), .C1(new_n875), .C2(new_n841), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n668), .B(new_n863), .C1(new_n867), .C2(new_n876), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(G141gat), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n631), .A2(new_n572), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n866), .A2(new_n641), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n668), .A2(new_n440), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT117), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n588), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT58), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n845), .A2(KEYINPUT118), .A3(new_n879), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT118), .B1(new_n845), .B2(new_n879), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n588), .A4(new_n882), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT58), .B1(new_n877), .B2(G141gat), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n880), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n845), .A2(KEYINPUT118), .A3(new_n879), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n588), .A3(new_n882), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT119), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n890), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n885), .A2(new_n897), .ZN(G1344gat));
  NAND2_X1  g697(.A1(new_n863), .A2(new_n278), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n324), .A2(new_n669), .A3(new_n325), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n875), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n636), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n868), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n866), .A2(new_n636), .A3(new_n865), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT59), .B1(new_n905), .B2(new_n441), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n441), .A2(KEYINPUT59), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n863), .B1(new_n867), .B2(new_n876), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n279), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n279), .A2(G148gat), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n893), .A2(new_n588), .A3(new_n894), .A4(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(KEYINPUT120), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(KEYINPUT120), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G1345gat));
  NAND2_X1  g714(.A1(new_n469), .A2(new_n447), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n893), .A2(new_n894), .ZN(new_n917));
  OR4_X1    g716(.A1(new_n916), .A2(new_n917), .A3(new_n642), .A4(new_n751), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n908), .B2(new_n751), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1346gat));
  OAI21_X1  g719(.A(G162gat), .B1(new_n908), .B2(new_n321), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n705), .A2(new_n453), .A3(new_n588), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n917), .B2(new_n922), .ZN(G1347gat));
  NAND2_X1  g722(.A1(new_n638), .A2(new_n642), .ZN(new_n924));
  AOI211_X1 g723(.A(new_n641), .B(new_n924), .C1(new_n840), .C2(new_n841), .ZN(new_n925));
  INV_X1    g724(.A(G169gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n668), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT121), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n641), .A2(new_n588), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(new_n695), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n842), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n669), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n932), .ZN(G1348gat));
  OAI21_X1  g732(.A(G176gat), .B1(new_n931), .B2(new_n279), .ZN(new_n934));
  INV_X1    g733(.A(G176gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n925), .A2(new_n935), .A3(new_n278), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1349gat));
  NAND3_X1  g736(.A1(new_n842), .A2(new_n231), .A3(new_n930), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT123), .B1(new_n938), .B2(G183gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n231), .A2(new_n399), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n925), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n925), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n842), .A2(new_n705), .A3(new_n930), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(G190gat), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(KEYINPUT125), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(KEYINPUT125), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n947), .A2(KEYINPUT125), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n925), .A2(new_n347), .A3(new_n705), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n925), .A2(KEYINPUT124), .A3(new_n347), .A4(new_n705), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n951), .A2(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n950), .A2(new_n957), .ZN(G1351gat));
  NAND4_X1  g757(.A1(new_n866), .A2(new_n632), .A3(new_n642), .A4(new_n879), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT126), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n668), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n675), .A2(new_n929), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n903), .B2(new_n904), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n668), .A2(G197gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  XNOR2_X1  g764(.A(KEYINPUT127), .B(G204gat), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n959), .A2(new_n279), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n963), .A2(new_n278), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n966), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n960), .A2(new_n385), .A3(new_n231), .ZN(new_n972));
  INV_X1    g771(.A(new_n962), .ZN(new_n973));
  INV_X1    g772(.A(new_n904), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT57), .B1(new_n901), .B2(new_n636), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n231), .B(new_n973), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  NAND3_X1  g778(.A1(new_n960), .A2(new_n386), .A3(new_n705), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n963), .A2(new_n705), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n386), .ZN(G1355gat));
endmodule


