//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  AND3_X1   g002(.A1(KEYINPUT76), .A2(G125), .A3(G140), .ZN(new_n189));
  AOI21_X1  g003(.A(G140), .B1(KEYINPUT76), .B2(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT16), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT77), .B1(new_n193), .B2(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT77), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n195), .A2(new_n196), .A3(new_n192), .A4(G125), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n191), .A2(new_n194), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n191), .A2(new_n194), .A3(G146), .A4(new_n197), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT24), .B(G110), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT72), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G119), .B(G128), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n200), .A2(new_n201), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT75), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT73), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(G128), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(KEYINPUT23), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT23), .B1(new_n213), .B2(G119), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT73), .B1(new_n213), .B2(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n216), .A3(KEYINPUT74), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G110), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT74), .B1(new_n212), .B2(new_n216), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n207), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n219), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n221), .A2(KEYINPUT75), .A3(G110), .A4(new_n217), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n206), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G125), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G140), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n193), .A2(new_n225), .A3(new_n199), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n204), .A2(new_n205), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n212), .A2(new_n216), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G110), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n201), .B(new_n226), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G137), .ZN(new_n232));
  INV_X1    g046(.A(G221), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n233), .A2(new_n187), .A3(G953), .ZN(new_n234));
  XOR2_X1   g048(.A(new_n232), .B(new_n234), .Z(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n230), .A3(new_n235), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  AOI21_X1  g054(.A(G902), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n239), .A2(new_n240), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n188), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n243), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n237), .A2(new_n245), .A3(new_n238), .A4(new_n241), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n237), .A2(new_n238), .ZN(new_n247));
  AOI21_X1  g061(.A(G902), .B1(new_n187), .B2(G217), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n244), .A2(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G472), .A2(G902), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(G101), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n199), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n199), .A2(G143), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n262), .A2(new_n213), .B1(KEYINPUT1), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n261), .A3(new_n265), .A4(G128), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(G137), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT11), .A3(G134), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(G137), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n270), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n271), .A2(G134), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n269), .A2(G137), .ZN(new_n277));
  OAI21_X1  g091(.A(G131), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n267), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n270), .A2(new_n274), .A3(new_n272), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G131), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n275), .ZN(new_n283));
  AND2_X1   g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT64), .B1(new_n262), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(G143), .B(G146), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n284), .ZN(new_n289));
  NOR2_X1   g103(.A1(KEYINPUT0), .A2(G128), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n286), .A2(new_n289), .B1(new_n262), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n283), .B1(new_n292), .B2(KEYINPUT65), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n262), .A2(new_n291), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n288), .B1(new_n287), .B2(new_n284), .ZN(new_n295));
  AND4_X1   g109(.A1(new_n288), .A2(new_n259), .A3(new_n261), .A4(new_n284), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n280), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n302));
  INV_X1    g116(.A(G113), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT2), .A2(G113), .ZN(new_n307));
  XNOR2_X1  g121(.A(G116), .B(G119), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(new_n306), .B2(new_n307), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n300), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n263), .A2(KEYINPUT1), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n287), .B2(G128), .ZN(new_n316));
  INV_X1    g130(.A(new_n266), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n262), .A2(new_n213), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n319), .A2(KEYINPUT67), .A3(new_n315), .A4(new_n266), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n279), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n292), .A2(new_n283), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n311), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n258), .B1(new_n313), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n323), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(KEYINPUT28), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n257), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT30), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n267), .A2(new_n279), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n297), .A2(new_n298), .B1(new_n275), .B2(new_n282), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n286), .A2(new_n289), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT65), .A3(new_n294), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n312), .B(new_n328), .C1(new_n333), .C2(KEYINPUT30), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n325), .A2(new_n257), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT31), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n334), .A2(KEYINPUT31), .A3(new_n335), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n327), .B(KEYINPUT68), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n335), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT31), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n334), .A2(KEYINPUT31), .A3(new_n335), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT68), .B1(new_n344), .B2(new_n327), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n251), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT32), .ZN(new_n347));
  INV_X1    g161(.A(new_n251), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n323), .B1(new_n333), .B2(new_n311), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n326), .B1(new_n349), .B2(KEYINPUT28), .ZN(new_n350));
  OAI22_X1  g164(.A1(new_n337), .A2(new_n336), .B1(new_n350), .B2(new_n256), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT68), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n348), .B1(new_n353), .B2(new_n338), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT32), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n358));
  INV_X1    g172(.A(G902), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n321), .A2(new_n322), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n312), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n361), .A2(new_n323), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(new_n258), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n257), .B1(new_n258), .B2(new_n323), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT29), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n359), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n297), .A2(new_n298), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n332), .A3(new_n283), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n311), .B1(new_n368), .B2(new_n280), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT28), .B1(new_n369), .B2(new_n325), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n370), .A2(new_n364), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n370), .B2(new_n364), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT29), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT70), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n334), .A2(new_n323), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(new_n257), .ZN(new_n377));
  AOI211_X1 g191(.A(KEYINPUT70), .B(new_n256), .C1(new_n334), .C2(new_n323), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n366), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G472), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n358), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n366), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n376), .A2(new_n257), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT70), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n376), .A2(new_n375), .A3(new_n257), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n370), .A2(new_n364), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT69), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n370), .A2(new_n364), .A3(new_n371), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n383), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT71), .A3(G472), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n382), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n250), .B1(new_n357), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n252), .A2(G143), .A3(G214), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(G143), .B1(new_n252), .B2(G214), .ZN(new_n399));
  OAI21_X1  g213(.A(G131), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT17), .ZN(new_n401));
  INV_X1    g215(.A(G237), .ZN(new_n402));
  INV_X1    g216(.A(G953), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G214), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n260), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n273), .A3(new_n397), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(KEYINPUT17), .B(G131), .C1(new_n398), .C2(new_n399), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n407), .A2(new_n200), .A3(new_n201), .A4(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G113), .B(G122), .ZN(new_n410));
  INV_X1    g224(.A(G104), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(KEYINPUT18), .A2(G131), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n405), .A2(new_n397), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT18), .B(G131), .C1(new_n398), .C2(new_n399), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT76), .A2(G125), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n192), .ZN(new_n417));
  NAND3_X1  g231(.A1(KEYINPUT76), .A2(G125), .A3(G140), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(G146), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n419), .A2(new_n420), .A3(new_n226), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n420), .B1(new_n419), .B2(new_n226), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n414), .B(new_n415), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n409), .A2(new_n412), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n412), .B1(new_n409), .B2(new_n423), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n359), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G475), .ZN(new_n427));
  NOR2_X1   g241(.A1(G475), .A2(G902), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n417), .A2(KEYINPUT19), .A3(new_n418), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n193), .A2(new_n225), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n431), .A3(new_n199), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n201), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n400), .A2(new_n406), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n201), .A2(KEYINPUT87), .A3(new_n432), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n412), .B1(new_n438), .B2(new_n423), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n428), .B1(new_n439), .B2(new_n424), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(KEYINPUT20), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n436), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT87), .B1(new_n201), .B2(new_n432), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n423), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n412), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n409), .A2(new_n423), .A3(new_n412), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n442), .B1(new_n449), .B2(new_n428), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n427), .B1(new_n441), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT9), .B(G234), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(G217), .A3(new_n403), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT88), .B(new_n457), .C1(new_n213), .C2(G143), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n213), .A2(G143), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n260), .A2(G128), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT88), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n456), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n461), .A2(new_n457), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n457), .B1(new_n213), .B2(G143), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT88), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(KEYINPUT89), .A3(new_n459), .A4(new_n458), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n463), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G134), .ZN(new_n471));
  XNOR2_X1  g285(.A(G116), .B(G122), .ZN(new_n472));
  INV_X1    g286(.A(G107), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G116), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(G122), .ZN(new_n476));
  INV_X1    g290(.A(G122), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(G116), .ZN(new_n478));
  OAI21_X1  g292(.A(G107), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n461), .A2(new_n459), .A3(new_n269), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n471), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n485), .A2(new_n477), .A3(G116), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n473), .B(new_n486), .C1(new_n485), .C2(new_n472), .ZN(new_n487));
  INV_X1    g301(.A(new_n481), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n269), .B1(new_n461), .B2(new_n459), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n474), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n455), .B1(new_n484), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n482), .B1(new_n470), .B2(G134), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n494), .A2(new_n491), .A3(new_n454), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n359), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G478), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n496), .B(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n403), .A2(G952), .ZN(new_n500));
  NAND2_X1  g314(.A1(G234), .A2(G237), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(G902), .A3(G953), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT21), .B(G898), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n451), .A2(new_n499), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(G214), .B1(G237), .B2(G902), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT3), .B1(new_n411), .B2(G107), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT3), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n473), .A3(G104), .ZN(new_n513));
  INV_X1    g327(.A(G101), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n411), .A2(G107), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n511), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n411), .A2(G107), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n473), .A2(G104), .ZN(new_n518));
  OAI21_X1  g332(.A(G101), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n521));
  OR2_X1    g335(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g336(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n522), .A2(G116), .A3(new_n209), .A4(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n525));
  NAND2_X1  g339(.A1(new_n209), .A2(G116), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n475), .A2(G119), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n524), .B(G113), .C1(new_n525), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n520), .A2(new_n521), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n511), .A2(new_n513), .A3(new_n515), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT4), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(G101), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n309), .B2(new_n310), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(G101), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n535), .A2(KEYINPUT4), .A3(new_n516), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n530), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT82), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n539), .B(new_n530), .C1(new_n534), .C2(new_n536), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(KEYINPUT6), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n537), .A2(new_n544), .A3(new_n540), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n403), .A2(G224), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n546), .B(KEYINPUT83), .Z(new_n547));
  AOI21_X1  g361(.A(new_n224), .B1(new_n331), .B2(new_n294), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n264), .A2(new_n224), .A3(new_n266), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n547), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n297), .A2(G125), .ZN(new_n552));
  INV_X1    g366(.A(new_n547), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n549), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n543), .A2(new_n545), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n548), .B2(new_n550), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n552), .A2(KEYINPUT7), .A3(new_n547), .A4(new_n549), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT85), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n516), .A2(new_n519), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n309), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT84), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT5), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n564), .B1(new_n528), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n308), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(G113), .A3(new_n567), .A4(new_n524), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n529), .A2(new_n521), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n563), .A2(new_n568), .B1(new_n569), .B2(new_n562), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n539), .A2(KEYINPUT8), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT8), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n538), .A2(KEYINPUT82), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n538), .A2(KEYINPUT82), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n561), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n563), .A2(new_n568), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n569), .A2(new_n562), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n539), .B(KEYINPUT8), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(KEYINPUT85), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n560), .A2(new_n542), .A3(new_n577), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n556), .A2(new_n359), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(G210), .B1(G237), .B2(G902), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n556), .A2(new_n583), .A3(new_n359), .A4(new_n585), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n510), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n233), .B1(new_n453), .B2(new_n359), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n266), .A2(KEYINPUT79), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT79), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n287), .A2(new_n593), .A3(new_n265), .A4(G128), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n264), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n520), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n283), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n535), .A2(KEYINPUT4), .A3(new_n516), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n292), .A2(new_n600), .A3(new_n533), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n318), .A2(KEYINPUT10), .A3(new_n320), .A4(new_n520), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n598), .A2(new_n599), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(G110), .B(G140), .ZN(new_n604));
  INV_X1    g418(.A(G227), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(G953), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n604), .B(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT80), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n283), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n603), .A2(KEYINPUT80), .A3(new_n608), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n562), .A2(new_n264), .A3(new_n266), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n596), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT12), .B1(new_n617), .B2(new_n283), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT12), .ZN(new_n619));
  AOI211_X1 g433(.A(new_n619), .B(new_n599), .C1(new_n596), .C2(new_n616), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n603), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n607), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n615), .A2(G469), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(G469), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n603), .B(new_n608), .C1(new_n618), .C2(new_n620), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n608), .B1(new_n613), .B2(new_n603), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n625), .B(new_n359), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n625), .A2(new_n359), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n624), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n508), .A2(new_n589), .A3(new_n591), .A4(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n396), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  AND3_X1   g450(.A1(new_n632), .A2(new_n249), .A3(new_n591), .ZN(new_n637));
  AOI21_X1  g451(.A(G902), .B1(new_n353), .B2(new_n338), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n637), .B(new_n346), .C1(new_n381), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT90), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n510), .B(new_n507), .C1(new_n587), .C2(new_n588), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n496), .A2(KEYINPUT91), .A3(new_n497), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT91), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n460), .A2(new_n462), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n464), .B1(new_n644), .B2(KEYINPUT89), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n269), .B1(new_n645), .B2(new_n463), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n492), .B(new_n455), .C1(new_n646), .C2(new_n482), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n454), .B1(new_n494), .B2(new_n491), .ZN(new_n648));
  AOI21_X1  g462(.A(G902), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n643), .B1(new_n649), .B2(G478), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT33), .B1(new_n493), .B2(new_n495), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n647), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n497), .A2(G902), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n642), .A2(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n440), .A2(KEYINPUT20), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n449), .A2(new_n442), .A3(new_n428), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n657), .A2(new_n658), .B1(G475), .B2(new_n426), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n656), .A2(new_n659), .A3(KEYINPUT92), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT92), .ZN(new_n661));
  INV_X1    g475(.A(new_n653), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n652), .B1(new_n647), .B2(new_n648), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n655), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT91), .B1(new_n496), .B2(new_n497), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n649), .A2(new_n643), .A3(G478), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n661), .B1(new_n667), .B2(new_n451), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n641), .B1(new_n660), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT93), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT93), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n641), .B(new_n671), .C1(new_n660), .C2(new_n668), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n353), .A2(new_n338), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n359), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G472), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT90), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n346), .A4(new_n637), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n640), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT34), .B(G104), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G6));
  XOR2_X1   g495(.A(new_n507), .B(KEYINPUT94), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n589), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n659), .A2(new_n499), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n640), .A2(new_n678), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT35), .B(G107), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G9));
  NAND2_X1  g502(.A1(new_n244), .A2(new_n246), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n231), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n248), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT95), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT95), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n689), .A2(new_n695), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n633), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n354), .B1(new_n675), .B2(G472), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT37), .B(G110), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G12));
  NOR3_X1   g516(.A1(new_n380), .A2(new_n358), .A3(new_n381), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT71), .B1(new_n393), .B2(G472), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n355), .B1(new_n674), .B2(new_n251), .ZN(new_n705));
  AOI211_X1 g519(.A(KEYINPUT32), .B(new_n348), .C1(new_n353), .C2(new_n338), .ZN(new_n706));
  OAI22_X1  g520(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(G900), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n503), .B1(new_n505), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n684), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n689), .A2(new_n695), .A3(new_n692), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n695), .B1(new_n689), .B2(new_n692), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n613), .A2(new_n603), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n607), .ZN(new_n715));
  AOI21_X1  g529(.A(G902), .B1(new_n715), .B2(new_n626), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n630), .B1(new_n716), .B2(new_n625), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n590), .B1(new_n717), .B2(new_n624), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n713), .A2(new_n589), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n707), .A2(new_n710), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G128), .ZN(G30));
  XNOR2_X1  g535(.A(new_n649), .B(new_n498), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n693), .A2(new_n510), .A3(new_n722), .A4(new_n659), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n587), .A2(new_n588), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT38), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT96), .B(KEYINPUT39), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n709), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n718), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n726), .B1(KEYINPUT40), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n362), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n359), .B1(new_n731), .B2(new_n256), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n257), .B1(new_n334), .B2(new_n323), .ZN(new_n733));
  OAI21_X1  g547(.A(G472), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n357), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n730), .B(new_n735), .C1(KEYINPUT40), .C2(new_n729), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  NOR3_X1   g551(.A1(new_n656), .A2(new_n659), .A3(new_n709), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n707), .A2(new_n719), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  OAI21_X1  g554(.A(new_n359), .B1(new_n627), .B2(new_n628), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n591), .A3(new_n629), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n707), .A2(new_n673), .A3(new_n249), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT41), .B(G113), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT97), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n745), .B(new_n747), .ZN(G15));
  INV_X1    g562(.A(new_n684), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n744), .A2(new_n589), .A3(new_n682), .A4(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n396), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT98), .B(G116), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G18));
  INV_X1    g568(.A(new_n589), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n743), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n713), .A2(new_n756), .A3(new_n508), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n707), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT99), .B(G119), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G21));
  NAND4_X1  g574(.A1(new_n724), .A2(new_n509), .A3(new_n499), .A4(new_n451), .ZN(new_n761));
  INV_X1    g575(.A(new_n682), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n761), .A2(new_n743), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n363), .A2(new_n326), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n344), .B1(new_n256), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n251), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n676), .A2(new_n763), .A3(new_n249), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  AND2_X1   g582(.A1(new_n676), .A2(new_n766), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n693), .A3(new_n738), .A4(new_n756), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  INV_X1    g585(.A(KEYINPUT100), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n623), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT100), .B(new_n607), .C1(new_n621), .C2(new_n622), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(G469), .A3(new_n615), .A4(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n590), .B1(new_n717), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n587), .A2(new_n509), .A3(new_n588), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n776), .A2(new_n738), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n707), .A2(new_n249), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n396), .A2(KEYINPUT42), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G131), .ZN(G33));
  NAND3_X1  g599(.A1(new_n776), .A2(new_n710), .A3(new_n778), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n250), .B(new_n786), .C1(new_n357), .C2(new_n395), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n269), .ZN(G36));
  AND2_X1   g602(.A1(new_n615), .A2(new_n623), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(KEYINPUT45), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n773), .A2(KEYINPUT45), .A3(new_n615), .A4(new_n774), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(G469), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n631), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(KEYINPUT101), .A3(new_n629), .ZN(new_n794));
  INV_X1    g608(.A(new_n792), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n630), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(KEYINPUT46), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT101), .B1(new_n793), .B2(new_n629), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n591), .B(new_n728), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n699), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n656), .A2(new_n451), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT43), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n693), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n778), .B1(new_n804), .B2(KEYINPUT44), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n799), .B(new_n805), .C1(KEYINPUT44), .C2(new_n804), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n271), .ZN(G39));
  OAI21_X1  g621(.A(new_n591), .B1(new_n797), .B2(new_n798), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n347), .A2(new_n356), .B1(new_n382), .B2(new_n394), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n777), .A2(new_n249), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n812), .A2(new_n813), .A3(new_n738), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  AND2_X1   g630(.A1(new_n357), .A2(new_n734), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n744), .A2(new_n778), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n250), .A3(new_n502), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n451), .A3(new_n667), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT107), .Z(new_n822));
  AND4_X1   g636(.A1(new_n249), .A2(new_n769), .A3(new_n503), .A4(new_n802), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n725), .A2(new_n509), .A3(new_n743), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT50), .Z(new_n826));
  AND4_X1   g640(.A1(new_n503), .A2(new_n802), .A3(new_n744), .A4(new_n778), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n693), .A3(new_n769), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n822), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT108), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n822), .A2(new_n826), .A3(KEYINPUT108), .A4(new_n828), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n742), .A2(new_n629), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT102), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n590), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n810), .A2(new_n811), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n823), .A2(new_n778), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n831), .A2(new_n832), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT109), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n823), .A2(new_n756), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n660), .A2(new_n668), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n500), .B1(new_n820), .B2(new_n845), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n844), .A2(KEYINPUT111), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT111), .B1(new_n844), .B2(new_n846), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT48), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n396), .A2(new_n827), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(KEYINPUT48), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n851), .B(new_n852), .Z(new_n853));
  NAND3_X1  g667(.A1(new_n847), .A2(new_n848), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n829), .A2(new_n840), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n836), .A2(KEYINPUT110), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n836), .A2(KEYINPUT110), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n837), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n843), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n761), .A2(new_n693), .A3(new_n709), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(new_n776), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n735), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n770), .A2(new_n720), .A3(new_n863), .A4(new_n739), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT52), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n683), .A2(new_n659), .A3(new_n656), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n640), .A2(new_n678), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n745), .A2(new_n686), .A3(new_n867), .ZN(new_n868));
  AOI221_X4 g682(.A(new_n250), .B1(new_n750), .B2(new_n633), .C1(new_n357), .C2(new_n395), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n713), .A2(new_n756), .A3(new_n508), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n700), .B(new_n767), .C1(new_n813), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n779), .A2(new_n676), .A3(new_n693), .A4(new_n766), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT103), .ZN(new_n875));
  INV_X1    g689(.A(new_n709), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n659), .A2(new_n722), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n875), .B1(new_n778), .B2(new_n878), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n777), .A2(new_n877), .A3(KEYINPUT103), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n718), .B(new_n713), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n874), .B1(new_n813), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n787), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT42), .B1(new_n396), .B2(new_n779), .ZN(new_n885));
  AND4_X1   g699(.A1(KEYINPUT42), .A2(new_n707), .A3(new_n249), .A4(new_n779), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n883), .B(new_n884), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT104), .B1(new_n873), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n707), .B(new_n249), .C1(new_n751), .C2(new_n634), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n707), .A2(new_n757), .B1(new_n699), .B2(new_n698), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n767), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n745), .A2(new_n686), .A3(new_n867), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT104), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n787), .B1(new_n782), .B2(new_n783), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n883), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n865), .B1(new_n888), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n770), .A2(new_n720), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n898), .A2(KEYINPUT52), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(KEYINPUT53), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(KEYINPUT53), .B2(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  INV_X1    g716(.A(new_n865), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n873), .A2(new_n887), .A3(KEYINPUT104), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n882), .B(new_n787), .C1(new_n782), .C2(new_n783), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n894), .B1(new_n905), .B2(new_n893), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT105), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT105), .B1(new_n897), .B2(KEYINPUT53), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT106), .B(KEYINPUT54), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n865), .A2(new_n909), .A3(new_n899), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n893), .A3(new_n905), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n902), .A2(new_n915), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n860), .A2(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n834), .B(KEYINPUT49), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n725), .A2(new_n250), .A3(new_n510), .A4(new_n590), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n918), .A2(new_n817), .A3(new_n801), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(G75));
  NOR2_X1   g735(.A1(new_n403), .A2(G952), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n924), .A2(G902), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n925), .B2(G210), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n543), .A2(new_n545), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(new_n555), .Z(new_n928));
  XNOR2_X1  g742(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n923), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n926), .B2(new_n931), .ZN(G51));
  INV_X1    g747(.A(new_n912), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n924), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(KEYINPUT114), .A3(new_n915), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT114), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n924), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n630), .B(KEYINPUT57), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n628), .B2(new_n627), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n925), .A2(new_n795), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n922), .B1(new_n941), .B2(new_n942), .ZN(G54));
  NAND2_X1  g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT115), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n925), .A2(new_n449), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT116), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n449), .B1(new_n925), .B2(new_n945), .ZN(new_n950));
  NOR4_X1   g764(.A1(new_n948), .A2(new_n949), .A3(new_n922), .A4(new_n950), .ZN(G60));
  XOR2_X1   g765(.A(new_n654), .B(KEYINPUT117), .Z(new_n952));
  XNOR2_X1  g766(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n936), .A2(new_n938), .A3(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n957), .A2(KEYINPUT119), .A3(new_n923), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT119), .B1(new_n957), .B2(new_n923), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n952), .B1(new_n916), .B2(new_n955), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT60), .Z(new_n963));
  AND2_X1   g777(.A1(new_n924), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n691), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n965), .B(new_n923), .C1(new_n247), .C2(new_n964), .ZN(new_n966));
  XNOR2_X1  g780(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G66));
  INV_X1    g782(.A(new_n506), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n403), .B1(new_n969), .B2(G224), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n873), .B2(new_n403), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n927), .B1(G898), .B2(new_n403), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT121), .Z(new_n973));
  XNOR2_X1  g787(.A(new_n971), .B(new_n973), .ZN(G69));
  OAI21_X1  g788(.A(new_n328), .B1(new_n333), .B2(KEYINPUT30), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n429), .A2(new_n431), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n975), .B(new_n976), .Z(new_n977));
  AND3_X1   g791(.A1(new_n770), .A2(new_n720), .A3(new_n739), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n806), .A2(new_n979), .ZN(new_n980));
  OR4_X1    g794(.A1(new_n813), .A2(new_n799), .A3(new_n250), .A4(new_n761), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n980), .A2(new_n815), .A3(new_n895), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n403), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n708), .A2(G953), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT124), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n977), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n978), .A2(new_n736), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT122), .Z(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n667), .A2(new_n451), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n777), .B(new_n729), .C1(new_n991), .C2(new_n684), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n806), .B1(new_n396), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n989), .A2(new_n815), .A3(new_n990), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n403), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n986), .B1(new_n995), .B2(new_n977), .ZN(new_n996));
  OAI21_X1  g810(.A(G953), .B1(new_n605), .B2(new_n708), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT123), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n997), .B1(new_n986), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n996), .B(new_n999), .Z(G72));
  XNOR2_X1  g814(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n381), .A2(new_n359), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n994), .B2(new_n873), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n733), .ZN(new_n1005));
  INV_X1    g819(.A(new_n340), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1003), .B1(new_n387), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT127), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n901), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1005), .A2(new_n923), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1003), .B1(new_n982), .B2(new_n873), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT126), .Z(new_n1012));
  NOR2_X1   g826(.A1(new_n376), .A2(new_n256), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1010), .B1(new_n1012), .B2(new_n1013), .ZN(G57));
endmodule


