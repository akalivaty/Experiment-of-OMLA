//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n210));
  XNOR2_X1  g0010(.A(new_n209), .B(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(new_n203), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n203), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT66), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n207), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n211), .B1(new_n214), .B2(new_n216), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G107), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(KEYINPUT17), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n212), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n256), .B1(new_n253), .B2(G20), .ZN(new_n257));
  AOI211_X1 g0057(.A(new_n252), .B(new_n255), .C1(new_n257), .C2(KEYINPUT81), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n257), .A2(KEYINPUT81), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n258), .A2(new_n259), .B1(new_n256), .B2(new_n255), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n251), .A2(new_n212), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT78), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT70), .ZN(new_n264));
  INV_X1    g0064(.A(G20), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G159), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G58), .A2(G68), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n215), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G20), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT77), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G159), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n267), .B2(new_n268), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n265), .B1(new_n215), .B2(new_n271), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT77), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n263), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n270), .A2(KEYINPUT77), .A3(new_n273), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n278), .B1(new_n276), .B2(new_n277), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(KEYINPUT78), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT75), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n266), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT75), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n286), .A2(new_n291), .A3(new_n265), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT7), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n265), .A4(new_n290), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT76), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n284), .A2(new_n285), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT76), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT7), .A4(new_n265), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n294), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n280), .A2(new_n283), .B1(new_n300), .B2(G68), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n262), .B1(new_n301), .B2(KEYINPUT16), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n303));
  NAND3_X1  g0103(.A1(new_n288), .A2(new_n265), .A3(new_n290), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n293), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(KEYINPUT80), .A3(new_n295), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT80), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n307), .A3(new_n293), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n306), .A2(G68), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n281), .A2(new_n282), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n261), .B1(new_n302), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G41), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(G1), .A3(G13), .ZN(new_n314));
  INV_X1    g0114(.A(G223), .ZN(new_n315));
  INV_X1    g0115(.A(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G226), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G1698), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n317), .B(new_n319), .C1(new_n284), .C2(new_n285), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G87), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G41), .ZN(new_n323));
  INV_X1    g0123(.A(G45), .ZN(new_n324));
  AOI21_X1  g0124(.A(G1), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(new_n314), .A3(G274), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n314), .A2(G232), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(G190), .B2(new_n330), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n250), .B1(new_n312), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n292), .A2(new_n293), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n296), .A2(new_n299), .ZN(new_n336));
  OAI21_X1  g0136(.A(G68), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n283), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT78), .B1(new_n281), .B2(new_n282), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n337), .B(KEYINPUT16), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(new_n252), .A3(new_n311), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n341), .A2(new_n333), .A3(new_n250), .A4(new_n260), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n260), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n320), .A2(new_n321), .ZN(new_n345));
  INV_X1    g0145(.A(new_n314), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n326), .A2(new_n328), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(G179), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT82), .ZN(new_n350));
  OAI21_X1  g0150(.A(G169), .B1(new_n322), .B2(new_n329), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT18), .B1(new_n344), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT18), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n357), .B(new_n354), .C1(new_n341), .C2(new_n260), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n334), .A2(new_n343), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n288), .A2(new_n290), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G238), .A2(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G232), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(new_n361), .C1(new_n362), .C2(G1698), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n346), .C1(G107), .C2(new_n360), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n314), .A2(G244), .A3(new_n327), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n326), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(G179), .ZN(new_n367));
  INV_X1    g0167(.A(G169), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(new_n366), .ZN(new_n369));
  INV_X1    g0169(.A(new_n256), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n269), .B1(G20), .B2(G77), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT68), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n266), .B2(G20), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n265), .A2(KEYINPUT68), .A3(G33), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n262), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n255), .A2(new_n219), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n262), .B1(G1), .B2(new_n265), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n219), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n369), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n366), .A2(G200), .ZN(new_n385));
  INV_X1    g0185(.A(G190), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n382), .C1(new_n386), .C2(new_n366), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n388), .B(KEYINPUT72), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n375), .A2(new_n376), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT69), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT69), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n375), .A2(new_n392), .A3(new_n376), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(G77), .A3(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n262), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n396), .A2(KEYINPUT11), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT12), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n254), .B2(G68), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n255), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n380), .C2(new_n203), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n396), .B2(KEYINPUT11), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  AND2_X1   g0204(.A1(KEYINPUT74), .A2(G169), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n362), .A2(G1698), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n360), .B(new_n406), .C1(G226), .C2(G1698), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n266), .A2(new_n227), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n314), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n314), .A2(new_n327), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n326), .B1(new_n218), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT13), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n410), .A2(KEYINPUT13), .A3(new_n412), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n404), .B(new_n405), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n415), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(G179), .A3(new_n413), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n413), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n404), .B1(new_n420), .B2(new_n405), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n403), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(G200), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(G190), .A3(new_n413), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(new_n397), .A3(new_n402), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  OR3_X1    g0226(.A1(new_n359), .A2(new_n389), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n316), .A2(G222), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n360), .B(new_n428), .C1(new_n315), .C2(new_n316), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n346), .C1(G77), .C2(new_n360), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n326), .C1(new_n318), .C2(new_n411), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n386), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n391), .A2(new_n370), .A3(new_n393), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n269), .A2(G150), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(KEYINPUT71), .B1(G20), .B2(new_n204), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT71), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n437), .A3(new_n434), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n262), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n255), .A2(new_n201), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n380), .B2(new_n201), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT9), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n435), .A2(KEYINPUT71), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n204), .A2(G20), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n438), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n252), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT9), .ZN(new_n447));
  INV_X1    g0247(.A(new_n441), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n432), .B1(new_n442), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n431), .A2(G200), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n442), .A2(new_n449), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT73), .ZN(new_n454));
  INV_X1    g0254(.A(new_n432), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT10), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n450), .B(new_n451), .C1(new_n454), .C2(KEYINPUT10), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n446), .A2(new_n448), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n431), .A2(new_n368), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n461), .C1(G179), .C2(new_n431), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n458), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n427), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n254), .A2(G97), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n253), .A2(G33), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n262), .A2(new_n254), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n468), .B2(G97), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT83), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n306), .A2(G107), .A3(new_n308), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT6), .ZN(new_n472));
  INV_X1    g0272(.A(G107), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n227), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n473), .A2(KEYINPUT6), .A3(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n269), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n470), .B1(new_n480), .B2(new_n252), .ZN(new_n481));
  AOI211_X1 g0281(.A(KEYINPUT83), .B(new_n262), .C1(new_n471), .C2(new_n479), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n469), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT84), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n469), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n324), .A2(G1), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(G41), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n490));
  OAI211_X1 g0290(.A(G257), .B(new_n314), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT4), .B1(new_n297), .B2(new_n226), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G1698), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n220), .B1(new_n288), .B2(new_n290), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(G1698), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n495), .A2(new_n497), .B1(G33), .B2(G283), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n494), .B(new_n498), .C1(KEYINPUT4), .C2(new_n495), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n492), .B1(new_n499), .B2(new_n346), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n253), .A2(G45), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(KEYINPUT5), .B2(new_n323), .ZN(new_n502));
  INV_X1    g0302(.A(G274), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n213), .B2(new_n313), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n502), .B(new_n504), .C1(KEYINPUT5), .C2(new_n323), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(G179), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n505), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n507), .B(new_n492), .C1(new_n499), .C2(new_n346), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n508), .B2(new_n368), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n484), .A2(new_n486), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n483), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n500), .A2(new_n505), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G200), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(G190), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n228), .A2(new_n316), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n360), .A2(new_n517), .B1(G33), .B2(G294), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n360), .A2(G250), .A3(new_n316), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n346), .ZN(new_n521));
  OAI211_X1 g0321(.A(G264), .B(new_n314), .C1(new_n489), .C2(new_n490), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n505), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n368), .ZN(new_n524));
  XOR2_X1   g0324(.A(KEYINPUT87), .B(KEYINPUT22), .Z(new_n525));
  NAND4_X1  g0325(.A1(new_n525), .A2(new_n265), .A3(G87), .A4(new_n360), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n266), .A2(new_n244), .A3(G20), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT88), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n265), .B2(G107), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT23), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT23), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n528), .B(new_n531), .C1(new_n265), .C2(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n527), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n265), .B(G87), .C1(new_n284), .C2(new_n285), .ZN(new_n534));
  NOR2_X1   g0334(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n526), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT24), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n526), .A2(new_n533), .A3(new_n539), .A4(new_n536), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n262), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n255), .A2(new_n473), .ZN(new_n542));
  OR2_X1    g0342(.A1(new_n542), .A2(KEYINPUT25), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(KEYINPUT25), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n473), .C2(new_n467), .ZN(new_n545));
  OAI221_X1 g0345(.A(new_n524), .B1(G179), .B2(new_n523), .C1(new_n541), .C2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n541), .A2(new_n545), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n521), .A2(G190), .A3(new_n505), .A4(new_n522), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n505), .A2(new_n522), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n314), .B1(new_n518), .B2(new_n519), .ZN(new_n551));
  OAI21_X1  g0351(.A(G200), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT89), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n548), .A2(KEYINPUT89), .A3(new_n553), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n547), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n373), .A2(new_n254), .ZN(new_n559));
  XNOR2_X1  g0359(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n390), .B2(new_n227), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n360), .A2(new_n265), .A3(G68), .ZN(new_n563));
  AOI21_X1  g0363(.A(G20), .B1(new_n560), .B2(new_n408), .ZN(new_n564));
  NOR3_X1   g0364(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n559), .B1(new_n566), .B2(new_n252), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n468), .A2(new_n373), .ZN(new_n568));
  INV_X1    g0368(.A(G179), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n314), .A2(G250), .A3(new_n501), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT85), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT85), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n314), .A2(new_n572), .A3(G250), .A4(new_n501), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n504), .A2(new_n487), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n220), .A2(G1698), .ZN(new_n576));
  OAI221_X1 g0376(.A(new_n576), .B1(G238), .B2(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G116), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n314), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n567), .A2(new_n568), .B1(new_n569), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n580), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n368), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n577), .A2(new_n578), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n346), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n570), .A2(KEYINPUT85), .B1(new_n504), .B2(new_n487), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(G190), .A3(new_n573), .A4(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(G200), .B1(new_n575), .B2(new_n579), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n467), .A2(new_n225), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n559), .B(new_n590), .C1(new_n566), .C2(new_n252), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n581), .A2(new_n583), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT21), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n297), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G264), .A2(G1698), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n228), .B2(G1698), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n595), .B(new_n346), .C1(new_n297), .C2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G270), .B(new_n314), .C1(new_n489), .C2(new_n490), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n505), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G169), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n262), .A2(G116), .A3(new_n254), .A4(new_n466), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n255), .A2(new_n244), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G283), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n605), .B(new_n265), .C1(G33), .C2(new_n227), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n244), .A2(G20), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n252), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT20), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n604), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n593), .B1(new_n601), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n598), .A2(new_n505), .A3(new_n599), .A4(G179), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n611), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n608), .A2(new_n609), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n603), .B(new_n602), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(KEYINPUT21), .A3(G169), .A4(new_n600), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n613), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n618), .B1(G200), .B2(new_n600), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n386), .B2(new_n600), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n592), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n464), .A2(new_n516), .A3(new_n558), .A4(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n590), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n567), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT91), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n591), .A2(KEYINPUT91), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT90), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n585), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n575), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n579), .A2(KEYINPUT90), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(G200), .B1(G190), .B2(new_n580), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(new_n629), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n368), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n581), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n636), .A2(new_n509), .A3(new_n483), .A4(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n484), .A2(new_n486), .A3(new_n509), .A4(new_n592), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n556), .A2(new_n557), .B1(new_n620), .B2(new_n546), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n636), .A2(new_n638), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n644), .A2(new_n646), .A3(new_n510), .A4(new_n515), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(new_n647), .A3(new_n638), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n464), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n349), .A2(new_n351), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n344), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT18), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n344), .A2(new_n357), .A3(new_n650), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n341), .A2(new_n333), .A3(new_n260), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n342), .ZN(new_n657));
  INV_X1    g0457(.A(new_n384), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n425), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n422), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n654), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n458), .A2(new_n459), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n462), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n649), .A2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(new_n620), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n253), .A2(new_n265), .A3(G13), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n612), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n620), .A2(new_n622), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n674), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT92), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n558), .B1(new_n548), .B2(new_n673), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n546), .A2(new_n673), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT93), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n620), .A2(new_n672), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n547), .B2(new_n673), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT94), .Z(G399));
  NAND2_X1  g0491(.A1(new_n565), .A2(new_n244), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT95), .ZN(new_n693));
  INV_X1    g0493(.A(new_n208), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n693), .A2(new_n253), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n216), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  NAND4_X1  g0499(.A1(new_n516), .A2(new_n558), .A3(new_n623), .A4(new_n673), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  INV_X1    g0501(.A(new_n523), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n500), .A2(new_n702), .A3(new_n580), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT96), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n614), .B(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT97), .B(new_n701), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n600), .A2(new_n569), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n512), .A2(new_n523), .A3(new_n634), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n614), .B(KEYINPUT96), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n582), .A2(new_n523), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n701), .A2(KEYINPUT97), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n709), .A2(new_n710), .A3(new_n500), .A4(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n706), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT31), .B1(new_n713), .B2(new_n672), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n700), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n642), .A2(new_n640), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT98), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT98), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n642), .A2(new_n721), .A3(new_n640), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n639), .A2(new_n640), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n720), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n638), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n620), .A2(new_n546), .ZN(new_n727));
  INV_X1    g0527(.A(new_n557), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT89), .B1(new_n548), .B2(new_n553), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n645), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n726), .B1(new_n731), .B2(new_n516), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n672), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n648), .A2(new_n673), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n718), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n699), .B1(new_n738), .B2(G1), .ZN(G364));
  INV_X1    g0539(.A(G13), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n253), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n695), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n679), .B(new_n745), .C1(G330), .C2(new_n677), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n212), .B1(G20), .B2(new_n368), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT100), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n360), .A2(G355), .A3(new_n208), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G116), .B2(new_n208), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n286), .A2(new_n291), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n694), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n324), .B2(new_n697), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n248), .A2(G45), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n754), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT99), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n752), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n569), .A2(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n265), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n331), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G77), .A2(new_n767), .B1(new_n770), .B2(G107), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n265), .A2(new_n386), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n764), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n771), .B1(new_n202), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n265), .B1(new_n775), .B2(G190), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n227), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n772), .A2(new_n768), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n225), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n774), .A2(new_n297), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n765), .A2(new_n775), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G159), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  NAND3_X1  g0584(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n785), .A2(new_n386), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n787), .A2(new_n203), .B1(new_n789), .B2(new_n201), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n778), .A2(new_n594), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n793), .A2(new_n769), .B1(new_n766), .B2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n792), .B(new_n795), .C1(G329), .C2(new_n782), .ZN(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n297), .B1(new_n773), .B2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT33), .B(G317), .Z(new_n799));
  INV_X1    g0599(.A(G294), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n787), .A2(new_n799), .B1(new_n800), .B2(new_n776), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n798), .B(new_n801), .C1(G326), .C2(new_n788), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n780), .A2(new_n791), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n750), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n744), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n763), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n749), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n677), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n746), .A2(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n658), .A2(new_n673), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n387), .B1(new_n382), .B2(new_n673), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n384), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n735), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n648), .A2(new_n673), .A3(new_n813), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n717), .A2(G330), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n744), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n750), .A2(new_n747), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n744), .B1(G77), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n778), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n360), .B(new_n777), .C1(G107), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n769), .A2(new_n225), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G311), .B2(new_n782), .ZN(new_n827));
  INV_X1    g0627(.A(new_n773), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G294), .A2(new_n828), .B1(new_n767), .B2(G116), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n786), .A2(G283), .B1(new_n788), .B2(G303), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n825), .A2(new_n827), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n769), .A2(new_n203), .B1(new_n781), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G50), .B2(new_n824), .ZN(new_n834));
  INV_X1    g0634(.A(new_n755), .ZN(new_n835));
  INV_X1    g0635(.A(new_n776), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(G58), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G143), .A2(new_n828), .B1(new_n767), .B2(G159), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  INV_X1    g0639(.A(G150), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n789), .B2(new_n839), .C1(new_n840), .C2(new_n787), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT34), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n834), .B(new_n837), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n831), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT101), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n804), .B1(new_n845), .B2(new_n846), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n823), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n813), .B2(new_n748), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n820), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT102), .Z(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  NOR2_X1   g0653(.A1(new_n741), .A2(new_n253), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n403), .A2(new_n672), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n422), .A2(new_n425), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n403), .B(new_n672), .C1(new_n419), .C2(new_n421), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n813), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n700), .B2(new_n716), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n303), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n261), .B1(new_n302), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(new_n670), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n359), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n344), .B2(new_n355), .ZN(new_n867));
  INV_X1    g0667(.A(new_n670), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT105), .B1(new_n344), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT105), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n870), .B(new_n670), .C1(new_n341), .C2(new_n260), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n655), .B(new_n867), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n650), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n655), .B1(new_n863), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n874), .B2(new_n864), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n865), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n865), .B2(new_n876), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n860), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n865), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n655), .B(new_n651), .C1(new_n869), .C2(new_n871), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n866), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n869), .A2(new_n871), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n657), .A2(new_n652), .A3(new_n653), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n883), .A2(new_n872), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n881), .B1(new_n886), .B2(KEYINPUT38), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n880), .B(new_n859), .C1(new_n700), .C2(new_n716), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n879), .A2(new_n880), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT107), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n464), .A2(new_n717), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(G330), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n654), .A2(new_n670), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n810), .B(KEYINPUT104), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n816), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n858), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n877), .A2(new_n878), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n422), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n673), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT39), .B1(new_n877), .B2(new_n878), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT39), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n881), .C1(new_n886), .C2(KEYINPUT38), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n734), .A2(new_n464), .A3(new_n737), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n664), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n854), .B1(new_n894), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n910), .B2(new_n894), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n214), .A2(new_n244), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n478), .B(KEYINPUT103), .Z(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT35), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n916), .B2(new_n915), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT36), .Z(new_n919));
  NAND3_X1  g0719(.A1(new_n697), .A2(G77), .A3(new_n271), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(G50), .B2(new_n203), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(G1), .A3(new_n740), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n912), .A2(new_n919), .A3(new_n922), .ZN(G367));
  OAI21_X1  g0723(.A(new_n516), .B1(new_n511), .B2(new_n673), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n509), .A2(new_n483), .A3(new_n672), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n688), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT42), .ZN(new_n928));
  INV_X1    g0728(.A(new_n926), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n510), .B1(new_n929), .B2(new_n546), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n928), .B1(new_n673), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n673), .B1(new_n628), .B2(new_n629), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n726), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n645), .B2(new_n932), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT108), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n931), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT109), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n931), .A2(new_n938), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n941), .B2(KEYINPUT109), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n943), .A2(new_n945), .B1(new_n685), .B2(new_n929), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n941), .A2(KEYINPUT109), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n685), .A2(new_n929), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(new_n942), .A4(new_n944), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n695), .B(KEYINPUT41), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n689), .A2(new_n926), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT45), .ZN(new_n952));
  OR3_X1    g0752(.A1(new_n689), .A2(KEYINPUT44), .A3(new_n926), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT44), .B1(new_n689), .B2(new_n926), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n684), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n951), .B(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n958), .A2(new_n685), .A3(new_n954), .A4(new_n953), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n688), .B(KEYINPUT110), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n679), .A2(KEYINPUT111), .B1(new_n683), .B2(new_n687), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n679), .A2(KEYINPUT111), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n956), .A2(new_n959), .A3(new_n738), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n950), .B1(new_n965), .B2(new_n738), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n946), .B(new_n949), .C1(new_n966), .C2(new_n743), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n752), .B1(new_n208), .B2(new_n372), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n757), .A2(new_n239), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n744), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT112), .B1(new_n824), .B2(G116), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT46), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n769), .A2(new_n227), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n773), .A2(new_n594), .B1(new_n766), .B2(new_n793), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(G317), .C2(new_n782), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n755), .B1(G107), .B2(new_n836), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n786), .A2(G294), .B1(new_n788), .B2(G311), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n972), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT113), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n770), .A2(G77), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n360), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT114), .Z(new_n982));
  NOR2_X1   g0782(.A1(new_n776), .A2(new_n203), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n787), .A2(new_n275), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(G143), .C2(new_n788), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G58), .A2(new_n824), .B1(new_n782), .B2(G137), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G150), .A2(new_n828), .B1(new_n767), .B2(G50), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n979), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n970), .B1(new_n990), .B2(new_n750), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n807), .B2(new_n934), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n967), .A2(new_n992), .ZN(G387));
  NAND2_X1  g0793(.A1(new_n683), .A2(new_n749), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n756), .B1(new_n236), .B2(new_n324), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n693), .A2(new_n208), .A3(new_n360), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n256), .A2(G50), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT50), .ZN(new_n998));
  AOI211_X1 g0798(.A(G45), .B(new_n693), .C1(G68), .C2(G77), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n995), .A2(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n208), .A2(G107), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n752), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n744), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n778), .A2(new_n219), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n973), .B(new_n1004), .C1(G150), .C2(new_n782), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n755), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT115), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n773), .A2(new_n201), .B1(new_n766), .B2(new_n203), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G159), .B2(new_n788), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n776), .A2(new_n372), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n786), .B2(new_n370), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1007), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G116), .A2(new_n770), .B1(new_n782), .B2(G326), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n778), .A2(new_n800), .B1(new_n776), .B2(new_n793), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G317), .A2(new_n828), .B1(new_n767), .B2(G303), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n789), .B2(new_n797), .C1(new_n794), .C2(new_n787), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n835), .B(new_n1013), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1012), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1003), .B1(new_n750), .B2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n964), .A2(new_n743), .B1(new_n994), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n964), .A2(new_n738), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n695), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n964), .A2(new_n738), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(G393));
  INV_X1    g0829(.A(KEYINPUT117), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n956), .A2(new_n959), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n1026), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n695), .A3(new_n965), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n956), .A2(new_n959), .A3(new_n743), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n245), .A2(new_n757), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n752), .B1(new_n227), .B2(new_n208), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n744), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n778), .A2(new_n203), .B1(new_n766), .B2(new_n256), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n826), .B(new_n1038), .C1(G143), .C2(new_n782), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n776), .A2(new_n219), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1040), .B(new_n835), .C1(G50), .C2(new_n786), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n789), .A2(new_n840), .B1(new_n773), .B2(new_n275), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT51), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n828), .A2(G311), .B1(G317), .B2(new_n788), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n297), .B1(new_n769), .B2(new_n473), .C1(new_n787), .C2(new_n594), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G116), .B2(new_n836), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n766), .A2(new_n800), .B1(new_n781), .B2(new_n797), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G283), .B2(new_n824), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1044), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT116), .Z(new_n1053));
  AOI21_X1  g0853(.A(new_n1037), .B1(new_n1053), .B2(new_n750), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n926), .B2(new_n807), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1034), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1030), .B1(new_n1033), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1033), .A2(new_n1030), .A3(new_n1056), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(G390));
  NAND2_X1  g0860(.A1(new_n464), .A2(new_n718), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n908), .A2(new_n664), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n858), .B1(new_n718), .B2(new_n813), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n818), .A2(new_n859), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n897), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n818), .A2(new_n859), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n858), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n818), .B2(new_n814), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n896), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n733), .B2(new_n813), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1062), .B1(new_n1065), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1066), .A2(KEYINPUT119), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n903), .A2(new_n905), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n898), .A2(new_n902), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT118), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n722), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n721), .B1(new_n642), .B2(new_n640), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n723), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n647), .A2(new_n638), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n673), .B(new_n813), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1067), .B1(new_n1082), .B2(new_n896), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n883), .A2(new_n872), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n885), .A2(new_n884), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT38), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n902), .B1(new_n1086), .B2(new_n877), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1077), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n902), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT38), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n655), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n870), .B1(new_n312), .B2(new_n670), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n344), .A2(KEYINPUT105), .A3(new_n868), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n866), .A2(new_n882), .B1(new_n1094), .B2(new_n867), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n885), .A2(new_n884), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1090), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1089), .B1(new_n1097), .B2(new_n881), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1098), .B(KEYINPUT118), .C1(new_n1067), .C2(new_n1070), .ZN(new_n1099));
  AOI221_X4 g0899(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .C1(new_n1088), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1074), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1088), .A2(new_n1099), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1073), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1083), .A2(new_n1087), .A3(new_n1077), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n672), .B(new_n814), .C1(new_n725), .C2(new_n732), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n858), .B1(new_n1107), .B2(new_n1069), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT118), .B1(new_n1108), .B2(new_n1098), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1103), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1074), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1102), .A2(new_n1103), .A3(new_n1101), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n1072), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1105), .A2(new_n1113), .A3(new_n695), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT120), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT120), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1105), .A2(new_n1113), .A3(new_n1116), .A4(new_n695), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n778), .A2(new_n840), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT53), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n767), .A2(new_n1121), .B1(new_n770), .B2(G50), .ZN(new_n1122));
  INV_X1    g0922(.A(G125), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1119), .B(new_n1122), .C1(new_n1123), .C2(new_n781), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n297), .B1(new_n828), .B2(G132), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n786), .A2(G137), .B1(new_n788), .B2(G128), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(new_n275), .C2(new_n776), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n779), .A2(new_n1040), .A3(new_n360), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n473), .B2(new_n787), .C1(new_n793), .C2(new_n789), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G116), .A2(new_n828), .B1(new_n782), .B2(G294), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n203), .B2(new_n769), .C1(new_n227), .C2(new_n766), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1124), .A2(new_n1127), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1132), .A2(new_n750), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n744), .B1(new_n370), .B2(new_n822), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(new_n1075), .C2(new_n747), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n743), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1115), .A2(new_n1117), .A3(new_n1137), .ZN(G378));
  XNOR2_X1  g0938(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n463), .B(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n460), .A2(new_n868), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n463), .A2(new_n1139), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n463), .A2(new_n1139), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1143), .A2(new_n460), .A3(new_n868), .A4(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n747), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n822), .A2(G50), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n773), .A2(new_n473), .B1(new_n766), .B2(new_n372), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n835), .A2(new_n323), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(G283), .C2(new_n782), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n769), .A2(new_n202), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1004), .A2(new_n1152), .A3(new_n983), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n786), .A2(G97), .B1(new_n788), .B2(G116), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT58), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G50), .B1(new_n266), .B2(new_n323), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1155), .A2(new_n1156), .B1(new_n1150), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G33), .B(G41), .C1(new_n782), .C2(G124), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G128), .A2(new_n828), .B1(new_n824), .B2(new_n1121), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT121), .Z(new_n1161));
  OAI22_X1  g0961(.A1(new_n766), .A2(new_n839), .B1(new_n776), .B2(new_n840), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n787), .A2(new_n832), .B1(new_n789), .B2(new_n1123), .ZN(new_n1163));
  OR3_X1    g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT59), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1159), .B1(new_n275), .B2(new_n769), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1158), .B1(new_n1156), .B2(new_n1155), .C1(new_n1167), .C2(new_n1169), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n745), .B(new_n1148), .C1(new_n1170), .C2(new_n750), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1147), .A2(new_n1171), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n900), .A2(new_n906), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n879), .A2(new_n880), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n887), .A2(new_n888), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(G330), .A3(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(new_n1146), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n889), .B2(G330), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1173), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1176), .A2(new_n1146), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n889), .A2(G330), .A3(new_n1178), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n907), .A3(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(KEYINPUT122), .B(new_n1172), .C1(new_n1184), .C2(new_n742), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n742), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1172), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1065), .A2(new_n1071), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1062), .B1(new_n1136), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT123), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1180), .A2(new_n1193), .A3(new_n1183), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1181), .A2(new_n907), .A3(new_n1182), .A4(KEYINPUT123), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(KEYINPUT57), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n695), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1062), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1113), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1190), .B1(new_n1197), .B2(new_n1201), .ZN(G375));
  NAND2_X1  g1002(.A1(new_n1067), .A2(new_n747), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n744), .B1(G68), .B2(new_n822), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n836), .A2(G50), .B1(G132), .B2(new_n788), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n787), .B2(new_n1120), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n778), .A2(new_n275), .B1(new_n766), .B2(new_n840), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G137), .B2(new_n828), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1152), .B1(G128), .B2(new_n782), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(new_n755), .A3(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G97), .A2(new_n824), .B1(new_n782), .B2(G303), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n473), .B2(new_n766), .C1(new_n793), .C2(new_n773), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1010), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n786), .A2(G116), .B1(new_n788), .B2(G294), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1213), .A2(new_n980), .A3(new_n1214), .A4(new_n297), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1206), .A2(new_n1210), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1204), .B1(new_n1216), .B2(new_n750), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1191), .A2(new_n743), .B1(new_n1203), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n950), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1073), .A2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1191), .A2(new_n1198), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1218), .B1(new_n1220), .B2(new_n1221), .ZN(G381));
  NAND4_X1  g1022(.A1(new_n1058), .A2(new_n967), .A3(new_n992), .A4(new_n1059), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n852), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(G381), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT124), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1114), .A2(new_n1137), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1114), .A2(new_n1137), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT124), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G375), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1226), .A2(new_n1231), .ZN(G407));
  OAI21_X1  g1032(.A(new_n1231), .B1(new_n1226), .B2(new_n671), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(G213), .ZN(G409));
  NOR3_X1   g1034(.A1(new_n1100), .A2(new_n1104), .A3(new_n1073), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1219), .B(new_n1200), .C1(new_n1235), .C2(new_n1062), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1194), .A2(new_n743), .A3(new_n1195), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1172), .A3(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1114), .A2(new_n1137), .A3(new_n1227), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1227), .B1(new_n1114), .B2(new_n1137), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G378), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1241), .B1(new_n1242), .B2(G375), .ZN(new_n1243));
  INV_X1    g1043(.A(G213), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(G343), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT60), .B1(new_n1221), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n695), .A3(new_n1073), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1221), .A2(new_n1247), .A3(KEYINPUT60), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1218), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(G384), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n852), .B(new_n1218), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1243), .A2(new_n1246), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT62), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1245), .A2(G2897), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1252), .A2(new_n1253), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n695), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1194), .A2(KEYINPUT57), .A3(new_n1195), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1199), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT57), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1192), .B2(new_n1184), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1264), .A2(new_n1266), .B1(new_n1189), .B2(new_n1185), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1230), .A2(new_n1228), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1267), .A2(G378), .B1(new_n1268), .B2(new_n1238), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1261), .B1(new_n1269), .B2(new_n1245), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT62), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1243), .A2(new_n1271), .A3(new_n1246), .A4(new_n1254), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1256), .A2(new_n1257), .A3(new_n1270), .A4(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1059), .ZN(new_n1274));
  OAI21_X1  g1074(.A(G387), .B1(new_n1274), .B2(new_n1057), .ZN(new_n1275));
  AND2_X1   g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  OAI21_X1  g1076(.A(KEYINPUT126), .B1(new_n1276), .B2(new_n1224), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1275), .A2(new_n1223), .A3(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1276), .A2(new_n1224), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1275), .A2(new_n1223), .B1(new_n1281), .B2(new_n1277), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1273), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1275), .A2(new_n1223), .A3(new_n1277), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1275), .A2(new_n1223), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1281), .A2(new_n1277), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1289), .B2(new_n1261), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1255), .A2(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1243), .A2(KEYINPUT63), .A3(new_n1246), .A4(new_n1254), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1288), .A2(new_n1290), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1284), .A2(new_n1294), .ZN(G405));
  NAND2_X1  g1095(.A1(new_n1267), .A2(G378), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1268), .A2(G375), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(KEYINPUT127), .A3(new_n1254), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1254), .A2(KEYINPUT127), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1296), .A2(new_n1297), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1283), .ZN(G402));
endmodule


