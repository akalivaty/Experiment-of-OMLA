//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT64), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n458), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n458), .A2(new_n460), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n458), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G124), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n460), .A2(G112), .ZN(new_n473));
  OAI21_X1  g048(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n474));
  OAI22_X1  g049(.A1(new_n471), .A2(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n465), .B(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n475), .B1(new_n477), .B2(G136), .ZN(G162));
  NAND2_X1  g053(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n479), .A2(new_n481), .A3(G126), .A4(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n479), .A2(new_n481), .A3(G138), .A4(new_n460), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n458), .A2(new_n489), .A3(G138), .A4(new_n460), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(G164));
  NAND2_X1  g066(.A1(G75), .A2(G543), .ZN(new_n492));
  INV_X1    g067(.A(G543), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT5), .B1(new_n493), .B2(KEYINPUT67), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G62), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT66), .A3(G50), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n494), .A2(new_n497), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n511), .A2(new_n504), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT68), .B(G88), .Z(new_n513));
  AOI22_X1  g088(.A1(new_n507), .A2(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n503), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(new_n504), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT70), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n506), .A2(G51), .B1(new_n511), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT71), .B(G52), .Z(new_n528));
  OAI22_X1  g103(.A1(new_n519), .A2(new_n527), .B1(new_n505), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n511), .A2(G64), .ZN(new_n531));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n529), .A2(new_n533), .ZN(G171));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n498), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT72), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(KEYINPUT72), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n512), .A2(G81), .B1(G43), .B2(new_n506), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(G188));
  NAND2_X1  g123(.A1(new_n512), .A2(G91), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT73), .ZN(new_n550));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  OR3_X1    g126(.A1(new_n505), .A2(KEYINPUT9), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n505), .B2(new_n551), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n498), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n552), .A2(new_n553), .B1(G651), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n550), .A2(new_n557), .ZN(G299));
  XNOR2_X1  g133(.A(G171), .B(KEYINPUT74), .ZN(G301));
  OAI211_X1 g134(.A(KEYINPUT76), .B(G651), .C1(new_n511), .C2(G74), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  AOI21_X1  g136(.A(G74), .B1(new_n494), .B2(new_n497), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n562), .B2(new_n530), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n511), .A2(new_n565), .A3(G87), .A4(new_n504), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n504), .A2(G87), .A3(new_n494), .A4(new_n497), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT75), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n506), .A2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n564), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND4_X1  g146(.A1(new_n511), .A2(KEYINPUT77), .A3(G86), .A4(new_n504), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n504), .A2(G86), .A3(new_n494), .A4(new_n497), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n530), .A2(KEYINPUT6), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT6), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  AND4_X1   g154(.A1(G48), .A2(new_n577), .A3(new_n579), .A4(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n494), .A2(new_n497), .A3(G61), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n580), .B1(new_n583), .B2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n576), .A2(new_n584), .ZN(G305));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n519), .A2(new_n586), .B1(new_n587), .B2(new_n505), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n511), .A2(G60), .ZN(new_n589));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n530), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n512), .A2(G92), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT10), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(G54), .B2(new_n506), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n498), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n530), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n601), .B2(new_n600), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n594), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n594), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NOR2_X1   g188(.A1(new_n542), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n605), .A2(new_n612), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g193(.A(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n460), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI22_X1  g196(.A1(new_n471), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n477), .B2(G135), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n458), .A2(new_n463), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT80), .B(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n626), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n624), .A2(new_n629), .ZN(G156));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2435), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT16), .B(G1341), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(G14), .B1(new_n636), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n636), .B2(new_n642), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2067), .B(G2678), .Z(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT18), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n646), .A2(new_n647), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n652), .A2(KEYINPUT17), .A3(new_n649), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n652), .B2(KEYINPUT17), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n653), .A2(new_n654), .A3(new_n648), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2096), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT81), .ZN(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  AOI22_X1  g242(.A1(new_n665), .A2(KEYINPUT20), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n662), .A3(new_n664), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n668), .B(new_n670), .C1(KEYINPUT20), .C2(new_n665), .ZN(new_n671));
  XOR2_X1   g246(.A(G1991), .B(G1996), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1981), .B(G1986), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n605), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G4), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G1348), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(G19), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n542), .B2(new_n679), .ZN(new_n684));
  AOI22_X1  g259(.A1(new_n681), .A2(new_n682), .B1(G1341), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G2090), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G35), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G162), .B2(new_n687), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT29), .Z(new_n690));
  OAI221_X1 g265(.A(new_n685), .B1(G1341), .B2(new_n684), .C1(new_n686), .C2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT23), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n679), .A2(G20), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n692), .B(new_n693), .C1(G299), .C2(G16), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n692), .B2(new_n693), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT89), .B(G1956), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n690), .A2(new_n686), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n687), .A2(G26), .ZN(new_n699));
  OR2_X1    g274(.A1(G104), .A2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n700), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n701));
  INV_X1    g276(.A(G128), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n471), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n477), .B2(G140), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n699), .B1(new_n704), .B2(new_n687), .ZN(new_n705));
  MUX2_X1   g280(.A(new_n699), .B(new_n705), .S(KEYINPUT28), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G2067), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n697), .A2(new_n698), .A3(new_n707), .ZN(new_n708));
  OAI22_X1  g283(.A1(new_n681), .A2(new_n682), .B1(G2067), .B2(new_n706), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n691), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n477), .A2(G139), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n463), .A2(G103), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT25), .Z(new_n713));
  AOI22_X1  g288(.A1(new_n458), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n711), .B(new_n713), .C1(new_n460), .C2(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G33), .B(new_n715), .S(G29), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2072), .ZN(new_n717));
  NOR2_X1   g292(.A1(G5), .A2(G16), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G171), .B2(G16), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1961), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n679), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n679), .ZN(new_n723));
  INV_X1    g298(.A(G1966), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G29), .A2(G32), .ZN(new_n726));
  INV_X1    g301(.A(new_n471), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G129), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT86), .B(KEYINPUT26), .Z(new_n729));
  AND3_X1   g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n463), .A2(G105), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n728), .A2(new_n731), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G141), .B2(new_n477), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n726), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  INV_X1    g314(.A(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G160), .B2(new_n687), .ZN(new_n743));
  INV_X1    g318(.A(G2084), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G27), .A2(G29), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G164), .B2(G29), .ZN(new_n747));
  INV_X1    g322(.A(G2078), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G11), .ZN(new_n750));
  INV_X1    g325(.A(G28), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT87), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT30), .B2(new_n751), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n752), .A2(KEYINPUT87), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n623), .B2(G29), .ZN(new_n757));
  AND3_X1   g332(.A1(new_n745), .A2(new_n749), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n721), .A2(new_n725), .A3(new_n738), .A4(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n710), .B1(KEYINPUT88), .B2(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G6), .B(G305), .S(G16), .Z(new_n761));
  XOR2_X1   g336(.A(KEYINPUT32), .B(G1981), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n679), .A2(G22), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G166), .B2(new_n679), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G1971), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G16), .A2(G23), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT84), .ZN(new_n769));
  NAND2_X1  g344(.A1(G288), .A2(new_n769), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n566), .A2(new_n568), .B1(G49), .B2(new_n506), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n771), .A2(KEYINPUT84), .A3(new_n564), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(G16), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT33), .B(G1976), .Z(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n765), .A2(G1971), .ZN(new_n778));
  NOR4_X1   g353(.A1(new_n767), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT83), .B(KEYINPUT34), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n687), .A2(G25), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n477), .A2(G131), .ZN(new_n784));
  INV_X1    g359(.A(G119), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n460), .A2(G107), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n787));
  OAI22_X1  g362(.A1(new_n471), .A2(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n783), .B1(new_n789), .B2(new_n687), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT35), .B(G1991), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n790), .B(new_n791), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n679), .A2(G24), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n592), .B2(new_n679), .ZN(new_n794));
  INV_X1    g369(.A(G1986), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n781), .A2(new_n782), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(KEYINPUT85), .A2(KEYINPUT36), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n759), .A2(KEYINPUT88), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n760), .A2(new_n799), .A3(new_n800), .ZN(G311));
  INV_X1    g376(.A(G311), .ZN(G150));
  INV_X1    g377(.A(G93), .ZN(new_n803));
  INV_X1    g378(.A(G55), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n519), .A2(new_n803), .B1(new_n804), .B2(new_n505), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n511), .A2(G67), .ZN(new_n806));
  NAND2_X1  g381(.A1(G80), .A2(G543), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n530), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G860), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT91), .B(KEYINPUT37), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n605), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT39), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT90), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT38), .ZN(new_n817));
  INV_X1    g392(.A(new_n809), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n542), .B(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n810), .B1(new_n817), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n813), .B1(new_n820), .B2(new_n821), .ZN(G145));
  XNOR2_X1  g397(.A(new_n626), .B(KEYINPUT94), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(new_n735), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n789), .B(new_n715), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(G162), .B(new_n469), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT93), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n623), .B(KEYINPUT92), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G164), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n727), .A2(G130), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n460), .A2(G118), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G142), .B2(new_n477), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n704), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n831), .B(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n829), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G37), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n829), .B2(new_n838), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT40), .Z(G395));
  NAND2_X1  g418(.A1(new_n818), .A2(new_n608), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n773), .B(G305), .Z(new_n846));
  XNOR2_X1  g421(.A(G303), .B(G290), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n850), .B(KEYINPUT42), .C1(new_n845), .C2(new_n848), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(KEYINPUT42), .B2(new_n850), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n615), .B(new_n819), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n604), .B(G299), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(KEYINPUT41), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(KEYINPUT41), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n854), .B2(new_n853), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n852), .B(new_n858), .Z(new_n859));
  OAI21_X1  g434(.A(new_n844), .B1(new_n859), .B2(new_n608), .ZN(G295));
  OAI21_X1  g435(.A(new_n844), .B1(new_n859), .B2(new_n608), .ZN(G331));
  NAND2_X1  g436(.A1(G286), .A2(G171), .ZN(new_n862));
  INV_X1    g437(.A(G301), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(G286), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n819), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n855), .B2(new_n856), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n865), .A2(new_n854), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n848), .ZN(new_n872));
  INV_X1    g447(.A(new_n848), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n868), .B2(new_n870), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n874), .A3(new_n840), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n866), .A2(new_n869), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(KEYINPUT98), .A3(new_n873), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT98), .B1(new_n878), .B2(new_n873), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(G37), .ZN(new_n881));
  AND4_X1   g456(.A1(KEYINPUT43), .A2(new_n872), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT44), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n875), .A2(KEYINPUT43), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n872), .A2(new_n881), .A3(new_n876), .A4(new_n879), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n888), .ZN(G397));
  INV_X1    g464(.A(KEYINPUT111), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n459), .A2(new_n460), .ZN(new_n891));
  XNOR2_X1  g466(.A(KEYINPUT99), .B(G40), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n891), .A2(new_n467), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G1384), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n488), .A2(new_n490), .ZN(new_n895));
  INV_X1    g470(.A(new_n486), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(KEYINPUT105), .B(G8), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n902));
  INV_X1    g477(.A(G1981), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n584), .A2(new_n903), .A3(new_n572), .A4(new_n575), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n576), .A2(KEYINPUT108), .A3(new_n903), .A4(new_n584), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n580), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n573), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT109), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n912), .A3(new_n573), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n583), .A2(G651), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(G1981), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n902), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT49), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n901), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n906), .A2(new_n907), .B1(new_n915), .B2(G1981), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n920), .A2(new_n902), .A3(KEYINPUT49), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n890), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n918), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT49), .B1(new_n920), .B2(new_n902), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(KEYINPUT111), .A3(new_n924), .A4(new_n901), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  AND4_X1   g501(.A1(KEYINPUT84), .A2(new_n564), .A3(new_n570), .A4(new_n569), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT84), .B1(new_n771), .B2(new_n564), .ZN(new_n928));
  OAI21_X1  g503(.A(G1976), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n773), .A2(new_n931), .A3(G1976), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(G1976), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT52), .B1(G288), .B2(new_n933), .ZN(new_n934));
  AND4_X1   g509(.A1(new_n901), .A2(new_n930), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT52), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n900), .B1(new_n929), .B2(KEYINPUT106), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(new_n932), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n926), .A2(KEYINPUT112), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT112), .B1(new_n926), .B2(new_n939), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(G164), .B2(G1384), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n897), .A2(KEYINPUT45), .A3(new_n894), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n893), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT102), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n943), .A2(new_n944), .A3(new_n947), .A4(new_n893), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1971), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n892), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n461), .A2(new_n468), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n897), .A2(new_n894), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(KEYINPUT50), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT50), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n897), .A2(new_n956), .A3(new_n894), .ZN(new_n957));
  XNOR2_X1  g532(.A(KEYINPUT103), .B(G2090), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n951), .A2(KEYINPUT104), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n961));
  AOI21_X1  g536(.A(G1971), .B1(new_n946), .B2(new_n948), .ZN(new_n962));
  INV_X1    g537(.A(new_n959), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G303), .A2(G8), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n960), .A2(new_n964), .A3(G8), .A4(new_n967), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n940), .A2(new_n941), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1976), .ZN(new_n970));
  INV_X1    g545(.A(G288), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n926), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n900), .B1(new_n972), .B2(new_n908), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT113), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n908), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n901), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n970), .B1(new_n770), .B2(new_n772), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n901), .B1(new_n978), .B2(new_n931), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT52), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n937), .A2(new_n932), .A3(new_n934), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n922), .B2(new_n925), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT112), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n926), .A2(new_n939), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n976), .B(new_n977), .C1(new_n989), .C2(new_n968), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n974), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n899), .B1(new_n962), .B2(new_n963), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n965), .B(KEYINPUT55), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n926), .A2(new_n968), .A3(new_n939), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n945), .A2(new_n724), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n998), .A2(new_n744), .A3(new_n957), .A4(new_n893), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(G168), .A3(new_n899), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n992), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n968), .A2(new_n995), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1001), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1003), .A2(KEYINPUT114), .A3(new_n984), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n960), .A2(G8), .A3(new_n964), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n994), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n968), .A2(KEYINPUT63), .A3(new_n1004), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n985), .A2(new_n988), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT126), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n946), .A2(new_n748), .A3(new_n948), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n943), .A2(new_n944), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT123), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n748), .A4(new_n893), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT123), .B1(new_n945), .B2(G2078), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(KEYINPUT53), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1961), .B1(new_n955), .B2(new_n957), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1017), .A2(new_n1022), .A3(G301), .A4(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n748), .A2(KEYINPUT124), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n748), .A2(KEYINPUT124), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT53), .B(G40), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n469), .A2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1018), .A2(new_n1029), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1023), .B(new_n1030), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1031));
  INV_X1    g606(.A(G171), .ZN(new_n1032));
  OAI211_X1 g607(.A(KEYINPUT54), .B(new_n1025), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(KEYINPUT125), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT125), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1030), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1017), .A2(new_n1024), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n1038), .B2(G171), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1039), .B2(new_n1025), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1041));
  AND4_X1   g616(.A1(G301), .A2(new_n1017), .A3(new_n1024), .A4(new_n1037), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1023), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1043));
  AOI21_X1  g618(.A(G301), .B1(new_n1043), .B2(new_n1022), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1036), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G286), .A2(new_n899), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1000), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(KEYINPUT122), .A3(new_n1000), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1000), .A2(new_n899), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1046), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n997), .B2(new_n999), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT51), .B1(new_n1047), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1052), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1003), .A2(new_n984), .A3(new_n1045), .A4(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1014), .B1(new_n1041), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1348), .B1(new_n955), .B2(new_n957), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n898), .A2(G2067), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n998), .A2(new_n957), .A3(new_n893), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n682), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1065), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT118), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT60), .B(new_n604), .C1(new_n1066), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT121), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT60), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n605), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1064), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1068), .A2(new_n1069), .A3(KEYINPUT118), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(KEYINPUT60), .A4(new_n604), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1072), .A2(new_n1074), .A3(new_n1079), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1077), .A2(KEYINPUT60), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n953), .A2(new_n954), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT58), .B(G1341), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n945), .A2(G1996), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n542), .ZN(new_n1086));
  XOR2_X1   g661(.A(new_n1086), .B(KEYINPUT59), .Z(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(KEYINPUT116), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1018), .A2(new_n893), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1090), .A2(KEYINPUT117), .B1(new_n1091), .B2(new_n1067), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G299), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n550), .A2(KEYINPUT57), .A3(new_n557), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1018), .A2(new_n1097), .A3(new_n893), .A4(new_n1089), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1092), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1099), .A2(KEYINPUT61), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1096), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1090), .A2(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1067), .A2(new_n1091), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1098), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1092), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1087), .B1(new_n1104), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1082), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n605), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1111), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1116), .B2(new_n1111), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1045), .A2(new_n1060), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1033), .A2(KEYINPUT125), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1039), .A2(new_n1035), .A3(new_n1025), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n996), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1122), .A2(new_n1125), .A3(KEYINPUT126), .A4(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1062), .A2(new_n1121), .A3(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1060), .A2(KEYINPUT62), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1060), .A2(KEYINPUT62), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1129), .A2(new_n1126), .A3(new_n1044), .A4(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n991), .A2(new_n1013), .A3(new_n1128), .A4(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n704), .B(G2067), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT101), .Z(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n735), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n954), .A2(new_n893), .A3(new_n942), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1136), .B(new_n1138), .C1(G1996), .C2(new_n1134), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1137), .A2(G1996), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT100), .Z(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n735), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n789), .B(new_n791), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1137), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n592), .B(new_n795), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n1138), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1132), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1141), .B(KEYINPUT46), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT47), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1137), .A2(G290), .A3(G1986), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT48), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n784), .A2(new_n791), .A3(new_n788), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1144), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(G2067), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n704), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1137), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1156), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1149), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1149), .A2(KEYINPUT127), .A3(new_n1162), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g742(.A(new_n842), .ZN(new_n1169));
  INV_X1    g743(.A(G319), .ZN(new_n1170));
  NOR4_X1   g744(.A1(G229), .A2(new_n1170), .A3(G401), .A4(G227), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n886), .A2(new_n1169), .A3(new_n1171), .ZN(G225));
  INV_X1    g746(.A(G225), .ZN(G308));
endmodule


