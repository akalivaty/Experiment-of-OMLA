//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1234, new_n1235, new_n1236, new_n1237;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT68), .B(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n464), .A2(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n473), .A2(new_n474), .B1(G101), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT69), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n459), .A2(new_n460), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(new_n474), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G138), .B1(new_n459), .B2(new_n460), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n468), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n471), .A2(new_n472), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n493), .A2(new_n474), .A3(G138), .A4(new_n489), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n498), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT70), .B1(new_n498), .B2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n505), .B1(new_n464), .B2(G114), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n498), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n496), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(G126), .A2(G2105), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n471), .B2(new_n472), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n495), .A2(new_n503), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  AND2_X1   g088(.A1(KEYINPUT73), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT73), .A2(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT6), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT75), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(G88), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G50), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(KEYINPUT74), .B1(new_n519), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  AOI211_X1 g104(.A(new_n529), .B(new_n526), .C1(new_n516), .C2(new_n518), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n525), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT76), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n533), .B(new_n525), .C1(new_n528), .C2(new_n530), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n524), .A2(G62), .ZN(new_n535));
  AND2_X1   g110(.A1(G75), .A2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT73), .B(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n532), .A2(new_n534), .B1(new_n537), .B2(new_n538), .ZN(G166));
  INV_X1    g114(.A(new_n523), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT5), .B1(KEYINPUT75), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n518), .B2(new_n516), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G89), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n545), .B1(new_n540), .B2(new_n541), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n522), .A2(KEYINPUT77), .A3(new_n523), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n548), .A2(G63), .A3(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  INV_X1    g126(.A(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n516), .B2(new_n518), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G51), .ZN(new_n554));
  AND4_X1   g129(.A1(new_n544), .A2(new_n549), .A3(new_n551), .A4(new_n554), .ZN(G168));
  INV_X1    g130(.A(new_n538), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n548), .A2(G64), .ZN(new_n557));
  NAND2_X1  g132(.A1(G77), .A2(G543), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n553), .A2(G52), .ZN(new_n560));
  INV_X1    g135(.A(new_n543), .ZN(new_n561));
  INV_X1    g136(.A(G90), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n559), .A2(new_n563), .ZN(G171));
  XNOR2_X1  g139(.A(KEYINPUT80), .B(G43), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n543), .A2(G81), .B1(new_n553), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n546), .A2(G56), .A3(new_n547), .ZN(new_n568));
  NAND2_X1  g143(.A1(G68), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT78), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n568), .A2(new_n572), .A3(new_n569), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n538), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n567), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n571), .A2(KEYINPUT79), .A3(new_n573), .A4(new_n538), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G860), .ZN(G153));
  NAND4_X1  g154(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g155(.A1(G1), .A2(G3), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT8), .ZN(new_n582));
  NAND4_X1  g157(.A1(G319), .A2(G483), .A3(G661), .A4(new_n582), .ZN(G188));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n584));
  OR2_X1    g159(.A1(KEYINPUT73), .A2(G651), .ZN(new_n585));
  NAND2_X1  g160(.A1(KEYINPUT73), .A2(G651), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(G91), .B(new_n524), .C1(new_n587), .C2(new_n517), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n524), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G651), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT9), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n553), .B2(G53), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g170(.A(G53), .B(G543), .C1(new_n587), .C2(new_n517), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT81), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n553), .A2(new_n593), .A3(G53), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT9), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G299));
  OR2_X1    g175(.A1(new_n559), .A2(new_n563), .ZN(G301));
  INV_X1    g176(.A(G168), .ZN(G286));
  INV_X1    g177(.A(G166), .ZN(G303));
  NAND2_X1  g178(.A1(new_n553), .A2(G49), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n519), .A2(G87), .A3(new_n524), .ZN(new_n605));
  AOI21_X1  g180(.A(G74), .B1(new_n546), .B2(new_n547), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n590), .ZN(G288));
  NAND3_X1  g182(.A1(new_n519), .A2(G86), .A3(new_n524), .ZN(new_n608));
  OAI211_X1 g183(.A(G48), .B(G543), .C1(new_n587), .C2(new_n517), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G61), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n522), .B2(new_n523), .ZN(new_n612));
  AND2_X1   g187(.A1(G73), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n538), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(G305));
  AOI22_X1  g190(.A1(new_n543), .A2(G85), .B1(new_n553), .B2(G47), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n548), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n556), .ZN(G290));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G301), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n553), .A2(G54), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT82), .B(G66), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n542), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G651), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n543), .A2(KEYINPUT10), .A3(G92), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(KEYINPUT10), .B1(new_n543), .B2(G92), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n621), .B(new_n625), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT83), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n620), .B1(new_n630), .B2(new_n619), .ZN(G284));
  XNOR2_X1  g206(.A(G284), .B(KEYINPUT84), .ZN(G321));
  NAND2_X1  g207(.A1(G299), .A2(new_n619), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n619), .B2(G168), .ZN(G297));
  OAI21_X1  g209(.A(new_n633), .B1(new_n619), .B2(G168), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n630), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n578), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(KEYINPUT85), .A2(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n493), .A2(new_n475), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  NOR2_X1   g220(.A1(KEYINPUT85), .A2(G2100), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n485), .A2(G123), .ZN(new_n648));
  OAI221_X1 g223(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n474), .C2(G111), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n483), .A2(G135), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT86), .B(G2096), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n647), .B(new_n653), .C1(new_n645), .C2(new_n642), .ZN(G156));
  XNOR2_X1  g229(.A(G2427), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT15), .B(G2435), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT87), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n661), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n661), .B(new_n665), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n668), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n672), .A3(G14), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT88), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT18), .Z(new_n683));
  INV_X1    g258(.A(new_n680), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n681), .B1(new_n684), .B2(new_n678), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n678), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n685), .B1(new_n688), .B2(new_n684), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n684), .A3(new_n681), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G2096), .B(G2100), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G227));
  XOR2_X1   g268(.A(G1971), .B(G1976), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n696), .A2(new_n697), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n695), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n695), .A2(new_n698), .A3(new_n702), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT92), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT91), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n706), .B(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G21), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G168), .B2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT99), .B(G1966), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(KEYINPUT31), .A2(G11), .ZN(new_n720));
  NAND2_X1  g295(.A1(KEYINPUT31), .A2(G11), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n651), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT30), .B(G28), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n722), .B(new_n724), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n719), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G171), .A2(new_n714), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n714), .A2(G5), .ZN(new_n729));
  OAI21_X1  g304(.A(G1961), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n716), .A2(new_n718), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n727), .A2(new_n730), .A3(KEYINPUT100), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n723), .A2(G26), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  AOI22_X1  g310(.A1(G128), .A2(new_n485), .B1(new_n483), .B2(G140), .ZN(new_n736));
  OAI221_X1 g311(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n474), .C2(G116), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n735), .B1(new_n738), .B2(G29), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n739), .A2(G2067), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(G2067), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n481), .A2(G29), .A3(new_n484), .A4(new_n486), .ZN(new_n742));
  OR2_X1    g317(.A1(G29), .A2(G35), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT29), .B(G2090), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n740), .A2(new_n741), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n723), .A2(G33), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  AOI22_X1  g326(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(new_n474), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n483), .A2(G139), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n749), .B1(new_n756), .B2(new_n723), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n748), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n723), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n723), .ZN(new_n763));
  INV_X1    g338(.A(G2078), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT24), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(G34), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(G34), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n477), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT97), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G2084), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n723), .A2(G32), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n485), .A2(G129), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT26), .Z(new_n778));
  NAND3_X1  g353(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(G29), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT98), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n765), .A2(new_n772), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G1348), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n714), .A2(G4), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n787), .B(new_n788), .C1(new_n630), .C2(new_n714), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n732), .A2(new_n761), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n731), .A2(new_n730), .A3(new_n719), .A4(new_n726), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT100), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n714), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT23), .Z(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n782), .A2(new_n784), .ZN(new_n799));
  INV_X1    g374(.A(new_n783), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n729), .B1(G301), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1961), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n771), .A2(G2084), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n801), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT101), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n788), .B1(new_n630), .B2(new_n714), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G1348), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT101), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n801), .A2(new_n804), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  AND4_X1   g386(.A1(new_n798), .A2(new_n807), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n578), .A2(G16), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G16), .B2(G19), .ZN(new_n814));
  INV_X1    g389(.A(G1341), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n794), .A2(new_n812), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n714), .A2(G22), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n714), .ZN(new_n821));
  INV_X1    g396(.A(G1971), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g398(.A(G1971), .B(new_n820), .C1(G166), .C2(new_n714), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT33), .B(G1976), .Z(new_n826));
  INV_X1    g401(.A(KEYINPUT95), .ZN(new_n827));
  NOR2_X1   g402(.A1(G16), .A2(G23), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT94), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n827), .B(new_n829), .C1(G288), .C2(new_n714), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(G651), .B1(new_n548), .B2(G74), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n832), .A2(G16), .A3(new_n605), .A4(new_n604), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n827), .B1(new_n833), .B2(new_n829), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n826), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n608), .A2(new_n609), .A3(new_n614), .A4(G16), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT32), .ZN(new_n837));
  OR2_X1    g412(.A1(G6), .A2(G16), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  OAI21_X1  g415(.A(G1981), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n836), .A2(new_n838), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT32), .ZN(new_n843));
  INV_X1    g418(.A(G1981), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n829), .B1(G288), .B2(new_n714), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT95), .ZN(new_n849));
  INV_X1    g424(.A(new_n826), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n849), .A2(new_n830), .A3(new_n850), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n835), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n825), .A2(new_n852), .A3(KEYINPUT96), .ZN(new_n853));
  AOI21_X1  g428(.A(KEYINPUT96), .B1(new_n825), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n819), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n825), .A2(new_n852), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n825), .A2(new_n852), .A3(KEYINPUT96), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(KEYINPUT34), .A3(new_n859), .ZN(new_n860));
  MUX2_X1   g435(.A(G24), .B(G290), .S(G16), .Z(new_n861));
  AND2_X1   g436(.A1(new_n861), .A2(G1986), .ZN(new_n862));
  AOI22_X1  g437(.A1(G119), .A2(new_n485), .B1(new_n483), .B2(G131), .ZN(new_n863));
  OAI221_X1 g438(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n474), .C2(G107), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  MUX2_X1   g440(.A(G25), .B(new_n865), .S(G29), .Z(new_n866));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G1991), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT93), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n866), .B(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n861), .A2(G1986), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n862), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n855), .A2(new_n860), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT36), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT36), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n855), .A2(new_n860), .A3(new_n874), .A4(new_n871), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n818), .B1(new_n873), .B2(new_n875), .ZN(G311));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n875), .ZN(new_n878));
  INV_X1    g453(.A(new_n818), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI211_X1 g455(.A(KEYINPUT102), .B(new_n818), .C1(new_n873), .C2(new_n875), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(G150));
  NAND2_X1  g457(.A1(new_n630), .A2(G559), .ZN(new_n883));
  XNOR2_X1  g458(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n548), .A2(G67), .ZN(new_n886));
  NAND2_X1  g461(.A1(G80), .A2(G543), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n556), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n553), .A2(G55), .ZN(new_n889));
  INV_X1    g464(.A(G93), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n561), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n576), .A2(new_n577), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n576), .B2(new_n577), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n885), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n898));
  AOI21_X1  g473(.A(G860), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  INV_X1    g475(.A(new_n892), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G860), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT37), .Z(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(G145));
  NOR2_X1   g479(.A1(new_n508), .A2(new_n510), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n495), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n865), .B(new_n644), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n738), .A2(new_n779), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n738), .A2(new_n779), .ZN(new_n910));
  INV_X1    g485(.A(G118), .ZN(new_n911));
  OAI21_X1  g486(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n468), .A2(new_n911), .B1(KEYINPUT104), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(KEYINPUT104), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n483), .A2(G142), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n485), .A2(G130), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n909), .A2(new_n910), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n909), .B2(new_n910), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n908), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n907), .A3(new_n918), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n906), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n923), .A3(new_n906), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n756), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n755), .B1(new_n928), .B2(new_n924), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n651), .B(new_n477), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(new_n487), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(new_n929), .ZN(new_n935));
  INV_X1    g510(.A(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g514(.A(G166), .B(G290), .ZN(new_n940));
  XNOR2_X1  g515(.A(G305), .B(G288), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n942), .B(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n896), .B(new_n638), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n625), .A2(new_n621), .ZN(new_n946));
  INV_X1    g521(.A(new_n628), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(new_n626), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n594), .A2(new_n592), .ZN(new_n949));
  NAND2_X1  g524(.A1(G78), .A2(G543), .ZN(new_n950));
  INV_X1    g525(.A(G65), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n542), .B2(new_n951), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n543), .A2(G91), .B1(new_n952), .B2(G651), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n599), .A2(new_n949), .A3(new_n953), .A4(KEYINPUT105), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT105), .B1(new_n595), .B2(new_n599), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n956), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(KEYINPUT41), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n955), .A2(new_n956), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n957), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT106), .B1(new_n945), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n962), .A2(new_n957), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n945), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n945), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n967), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n944), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n944), .B(new_n973), .C1(new_n969), .C2(new_n966), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(G868), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n901), .A2(new_n619), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(G295));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n978), .ZN(G331));
  OAI21_X1  g555(.A(G171), .B1(new_n894), .B2(new_n895), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n576), .A2(new_n577), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n901), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(G301), .A3(new_n893), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n981), .A2(G168), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(G168), .B1(new_n981), .B2(new_n984), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n985), .A2(new_n986), .A3(new_n964), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n894), .A2(new_n895), .A3(G171), .ZN(new_n988));
  AOI21_X1  g563(.A(G301), .B1(new_n983), .B2(new_n893), .ZN(new_n989));
  OAI21_X1  g564(.A(G286), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n981), .A2(new_n984), .A3(G168), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n968), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n942), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n967), .B1(new_n985), .B2(new_n986), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n965), .A2(new_n990), .A3(new_n991), .ZN(new_n995));
  INV_X1    g570(.A(new_n942), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n933), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n993), .A2(new_n933), .A3(new_n999), .A4(new_n997), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(KEYINPUT44), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n998), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n993), .A2(KEYINPUT43), .A3(new_n933), .A4(new_n997), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1003), .A2(new_n1008), .ZN(G397));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n906), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n469), .A2(new_n476), .A3(G40), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1014), .B(KEYINPUT110), .Z(new_n1015));
  OR2_X1    g590(.A1(new_n738), .A2(G2067), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n738), .A2(G2067), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1996), .ZN(new_n1019));
  INV_X1    g594(.A(new_n779), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1014), .A2(G1996), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1015), .A2(new_n1021), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1015), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n865), .B(new_n868), .Z(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OR3_X1    g601(.A1(new_n1014), .A2(G290), .A3(G1986), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G290), .A2(G1986), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1014), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT109), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n501), .A2(new_n502), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1033), .A2(new_n504), .B1(new_n492), .B2(new_n494), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n1034), .B2(new_n503), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT111), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n512), .B2(new_n1010), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n469), .A2(new_n476), .A3(G40), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1384), .B1(new_n495), .B2(new_n905), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(new_n1036), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1037), .A2(new_n1040), .A3(new_n1041), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1012), .A2(G1384), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1042), .B1(new_n512), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n717), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1032), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT51), .B1(new_n1051), .B2(KEYINPUT125), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1045), .A2(G168), .A3(new_n1050), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1053), .A2(G8), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G286), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1052), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT62), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(G166), .B2(new_n1032), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n512), .A2(new_n1010), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1012), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1042), .B1(new_n906), .B2(new_n1047), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n822), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT112), .B(G2090), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1042), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n512), .A2(new_n1036), .A3(new_n1010), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1064), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1037), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1069), .B1(new_n1077), .B2(new_n1070), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT113), .B(new_n1069), .C1(new_n1077), .C2(new_n1070), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1063), .A3(G8), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1043), .A2(new_n1013), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n1032), .ZN(new_n1085));
  INV_X1    g660(.A(G1976), .ZN(new_n1086));
  OR2_X1    g661(.A1(G288), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(KEYINPUT114), .A3(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1083), .A2(G8), .A3(new_n1086), .A4(G288), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G305), .A2(G1981), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n610), .A2(new_n844), .A3(new_n614), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT49), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(KEYINPUT49), .A3(new_n1094), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1085), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1044), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1103));
  AOI211_X1 g678(.A(KEYINPUT111), .B(new_n1036), .C1(new_n512), .C2(new_n1010), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n803), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1046), .A2(new_n1048), .A3(KEYINPUT53), .A4(new_n764), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1066), .A2(new_n764), .A3(new_n1067), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1105), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G171), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AND4_X1   g687(.A1(new_n1076), .A2(new_n1082), .A3(new_n1102), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1055), .A2(G8), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1056), .A2(G8), .A3(new_n1053), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1059), .A2(new_n1113), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1094), .ZN(new_n1124));
  NOR2_X1   g699(.A1(G288), .A2(G1976), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n1099), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1085), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1127), .B2(new_n1126), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1082), .A2(new_n1101), .A3(new_n1100), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G1956), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1072), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1013), .B1(new_n1043), .B2(new_n1036), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(G2072), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1066), .A2(new_n1067), .A3(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1139));
  NAND2_X1  g714(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT117), .Z(new_n1141));
  NAND4_X1  g716(.A1(new_n595), .A2(new_n599), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n599), .A2(new_n949), .A3(new_n953), .A4(new_n1139), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1141), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1135), .A2(new_n1138), .A3(new_n1142), .A4(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n787), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1083), .A2(G2067), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n629), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1135), .A2(new_n1138), .B1(new_n1145), .B2(new_n1142), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT119), .B(new_n1146), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1145), .A2(new_n1142), .ZN(new_n1154));
  AOI21_X1  g729(.A(G1956), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT45), .B1(new_n512), .B2(new_n1010), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1033), .B1(new_n492), .B2(new_n494), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1047), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1013), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1137), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1156), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1154), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1148), .B1(new_n1077), .B2(new_n787), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(new_n629), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT119), .B1(new_n1164), .B2(new_n1146), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1146), .B1(new_n1151), .B2(KEYINPUT122), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1154), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1168), .A2(new_n1169), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1167), .A2(KEYINPUT123), .A3(KEYINPUT61), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1162), .A2(new_n1146), .ZN(new_n1172));
  XNOR2_X1  g747(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(KEYINPUT120), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT58), .B(G1341), .Z(new_n1177));
  AOI22_X1  g752(.A1(new_n1176), .A2(new_n1019), .B1(new_n1083), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1175), .B1(new_n1178), .B2(new_n982), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1083), .A2(new_n1177), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1180), .B1(new_n1068), .B2(G1996), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1175), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n578), .A3(new_n1182), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1172), .A2(new_n1173), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n948), .A2(KEYINPUT124), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1147), .A2(KEYINPUT60), .A3(new_n1149), .A4(new_n1185), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n948), .A2(KEYINPUT124), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1186), .B(new_n1187), .C1(KEYINPUT60), .C2(new_n1163), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1189));
  AND4_X1   g764(.A1(new_n1171), .A2(new_n1184), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1167), .A2(KEYINPUT61), .A3(new_n1170), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1166), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1046), .A2(new_n1067), .A3(KEYINPUT53), .A4(new_n764), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1105), .A2(G301), .A3(new_n1109), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT54), .B1(new_n1111), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1105), .A2(new_n1109), .A3(new_n1195), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(G171), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1105), .A2(G301), .A3(new_n1109), .A4(new_n1106), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1200), .A2(KEYINPUT54), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1202), .A2(KEYINPUT126), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1200), .A2(new_n1204), .A3(KEYINPUT54), .A4(new_n1201), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1082), .A2(new_n1102), .A3(new_n1076), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1198), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1123), .B(new_n1131), .C1(new_n1194), .C2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1207), .A2(G168), .A3(new_n1051), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT63), .ZN(new_n1211));
  AND2_X1   g786(.A1(new_n1082), .A2(new_n1102), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1051), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1080), .A2(G8), .A3(new_n1081), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1213), .B1(new_n1214), .B2(new_n1064), .ZN(new_n1215));
  AOI22_X1  g790(.A1(new_n1210), .A2(new_n1211), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1031), .B1(new_n1209), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1018), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1015), .B1(new_n779), .B2(new_n1218), .ZN(new_n1219));
  XOR2_X1   g794(.A(new_n1022), .B(KEYINPUT46), .Z(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n1221), .B(KEYINPUT47), .ZN(new_n1222));
  XOR2_X1   g797(.A(new_n1027), .B(KEYINPUT48), .Z(new_n1223));
  OAI21_X1  g798(.A(new_n1222), .B1(new_n1026), .B2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n865), .A2(new_n868), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1023), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1024), .B1(new_n1226), .B2(new_n1016), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1228));
  AND2_X1   g803(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g804(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1230));
  NOR3_X1   g805(.A1(new_n1224), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1217), .A2(new_n1231), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g807(.A(new_n457), .ZN(new_n1234));
  NOR3_X1   g808(.A1(G229), .A2(new_n1234), .A3(G227), .ZN(new_n1235));
  OAI21_X1  g809(.A(new_n1235), .B1(new_n675), .B2(new_n676), .ZN(new_n1236));
  AOI21_X1  g810(.A(new_n1236), .B1(new_n937), .B2(new_n934), .ZN(new_n1237));
  AND3_X1   g811(.A1(new_n1237), .A2(new_n1005), .A3(new_n1006), .ZN(G308));
  NAND3_X1  g812(.A1(new_n1237), .A2(new_n1005), .A3(new_n1006), .ZN(G225));
endmodule


