//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AND2_X1   g0017(.A1(KEYINPUT65), .A2(G68), .ZN(new_n218));
  NOR2_X1   g0018(.A1(KEYINPUT65), .A2(G68), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G58), .A2(G232), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  INV_X1    g0039(.A(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT66), .B(G50), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G97), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT75), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT65), .B(G68), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OR2_X1    g0052(.A1(KEYINPUT12), .A2(G68), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n251), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n213), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n206), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G68), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n250), .A2(new_n207), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n207), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G77), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n263), .A2(new_n202), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n257), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT11), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n254), .B(new_n260), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n267), .A2(new_n268), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT67), .B1(new_n272), .B2(new_n213), .ZN(new_n273));
  AND2_X1   g0073(.A1(G1), .A2(G13), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT3), .ZN(new_n281));
  OR2_X1    g0081(.A1(G226), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G232), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n281), .A2(new_n282), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G97), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n279), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n206), .A2(new_n294), .B1(new_n274), .B2(new_n276), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n274), .B2(new_n276), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n295), .A2(G238), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n290), .A2(new_n291), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n278), .B1(new_n288), .B2(new_n287), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n274), .A2(new_n276), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n298), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n221), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT13), .ZN(new_n308));
  OAI211_X1 g0108(.A(G179), .B(new_n301), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n291), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n302), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n291), .B1(new_n290), .B2(new_n300), .ZN(new_n312));
  OAI21_X1  g0112(.A(G169), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT74), .B(KEYINPUT14), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n309), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT72), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n310), .B1(new_n302), .B2(new_n306), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n301), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n318), .A2(new_n322), .A3(KEYINPUT14), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(new_n323), .B2(KEYINPUT73), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n318), .A2(new_n322), .A3(new_n325), .A4(KEYINPUT14), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n271), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(G200), .B1(new_n311), .B2(new_n312), .ZN(new_n328));
  OAI211_X1 g0128(.A(G190), .B(new_n301), .C1(new_n307), .C2(new_n308), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n271), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n248), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n303), .B1(new_n285), .B2(new_n305), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G87), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT76), .B1(new_n280), .B2(KEYINPUT3), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT76), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(new_n283), .A3(G33), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n338), .A3(new_n281), .ZN(new_n339));
  INV_X1    g0139(.A(G226), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G1698), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G223), .B2(G1698), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n335), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n278), .B1(new_n343), .B2(KEYINPUT78), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT78), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n335), .C1(new_n339), .C2(new_n342), .ZN(new_n346));
  AOI211_X1 g0146(.A(new_n333), .B(new_n334), .C1(new_n344), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n343), .A2(KEYINPUT78), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(new_n346), .A3(new_n279), .ZN(new_n349));
  INV_X1    g0149(.A(new_n334), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n319), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT79), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n216), .B1(new_n220), .B2(new_n240), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(G20), .B1(G159), .B2(new_n262), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT7), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n339), .A2(new_n355), .A3(new_n207), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G68), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n355), .B1(new_n339), .B2(new_n207), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n354), .B(KEYINPUT16), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n201), .B1(new_n250), .B2(G58), .ZN(new_n361));
  INV_X1    g0161(.A(G159), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n361), .A2(new_n207), .B1(new_n362), .B2(new_n263), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT77), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT7), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT3), .B(G33), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(G20), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n281), .A2(new_n284), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n207), .A3(new_n366), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n220), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n360), .B1(new_n363), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n359), .A2(new_n373), .A3(new_n257), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT8), .B(G58), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n206), .B2(G20), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(new_n258), .B1(new_n255), .B2(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n349), .A2(G179), .A3(new_n350), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT79), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n334), .B1(new_n344), .B2(new_n346), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n379), .B(new_n380), .C1(new_n319), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n352), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT18), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n352), .A2(KEYINPUT18), .A3(new_n382), .A4(new_n378), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT80), .ZN(new_n388));
  INV_X1    g0188(.A(new_n378), .ZN(new_n389));
  INV_X1    g0189(.A(G190), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n349), .A2(new_n390), .A3(new_n350), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(G200), .B2(new_n381), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT17), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  AOI211_X1 g0193(.A(G190), .B(new_n334), .C1(new_n344), .C2(new_n346), .ZN(new_n394));
  AOI21_X1  g0194(.A(G200), .B1(new_n349), .B2(new_n350), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n396), .A2(new_n378), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n388), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(new_n396), .B2(new_n378), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n374), .A4(new_n377), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(KEYINPUT80), .A3(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n387), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G150), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n375), .A2(new_n264), .B1(new_n404), .B2(new_n263), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(G20), .B2(new_n203), .ZN(new_n406));
  INV_X1    g0206(.A(new_n257), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n258), .A2(G50), .A3(new_n259), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(G50), .B2(new_n251), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT9), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n409), .B1(G50), .B2(new_n251), .C1(new_n406), .C2(new_n407), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT9), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G223), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(G222), .B2(G1698), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n368), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n279), .B(new_n419), .C1(G77), .C2(new_n368), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n295), .A2(G226), .B1(new_n297), .B2(new_n299), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G200), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n420), .A2(new_n421), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G190), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n412), .A2(new_n415), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT10), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n411), .B1(new_n319), .B2(new_n422), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(G179), .B2(new_n422), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n258), .A2(G77), .A3(new_n259), .ZN(new_n430));
  XOR2_X1   g0230(.A(new_n430), .B(KEYINPUT69), .Z(new_n431));
  INV_X1    g0231(.A(new_n375), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n264), .B2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(new_n257), .B1(new_n265), .B2(new_n255), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G244), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n303), .B1(new_n438), .B2(new_n305), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT68), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n221), .A2(G1698), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(G232), .B2(G1698), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n368), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n279), .B(new_n444), .C1(G107), .C2(new_n368), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n439), .A2(new_n440), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n441), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G200), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n437), .B(new_n448), .C1(new_n390), .C2(new_n447), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n319), .A2(new_n447), .B1(new_n431), .B2(new_n436), .ZN(new_n450));
  INV_X1    g0250(.A(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n333), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n427), .A2(new_n429), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT14), .B1(new_n321), .B2(KEYINPUT72), .ZN(new_n456));
  AOI211_X1 g0256(.A(new_n317), .B(new_n319), .C1(new_n320), .C2(new_n301), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT73), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n316), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n326), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n271), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(KEYINPUT75), .A3(new_n330), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n332), .A2(new_n403), .A3(new_n455), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n427), .A2(new_n429), .A3(new_n454), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n330), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(new_n248), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n403), .A4(new_n463), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G264), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G1698), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(G257), .B2(G1698), .ZN(new_n474));
  INV_X1    g0274(.A(G303), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n339), .A2(new_n474), .B1(new_n475), .B2(new_n368), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n279), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n293), .A2(G1), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(G270), .A3(new_n304), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n297), .A2(new_n483), .A3(new_n478), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT85), .B(G116), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n251), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n206), .A2(G33), .ZN(new_n489));
  AND4_X1   g0289(.A1(new_n213), .A2(new_n251), .A3(new_n256), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n490), .B2(G116), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(G33), .B2(G283), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n280), .A2(G97), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n492), .A2(new_n493), .B1(new_n256), .B2(new_n213), .ZN(new_n494));
  OR2_X1    g0294(.A1(KEYINPUT85), .A2(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(KEYINPUT85), .A2(G116), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(G20), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT20), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n494), .A2(KEYINPUT20), .A3(new_n497), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n491), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n486), .A2(new_n500), .A3(KEYINPUT21), .A4(G169), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n500), .A2(G179), .A3(new_n477), .A4(new_n485), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n500), .B1(new_n486), .B2(G200), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n390), .B2(new_n486), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n486), .A2(new_n500), .A3(G169), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT21), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n506), .A2(KEYINPUT87), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT87), .B1(new_n506), .B2(new_n507), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n503), .B(new_n505), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT88), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(new_n507), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT87), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n506), .A2(KEYINPUT87), .A3(new_n507), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n517), .A2(KEYINPUT88), .A3(new_n503), .A4(new_n505), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G107), .ZN(new_n520));
  INV_X1    g0320(.A(new_n490), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT25), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n251), .A2(new_n522), .A3(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT25), .B1(new_n255), .B2(new_n520), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n520), .A2(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(new_n520), .A3(G20), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n280), .B1(new_n495), .B2(new_n496), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(new_n207), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n207), .A2(G87), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n370), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n336), .A2(new_n338), .A3(new_n207), .A4(new_n281), .ZN(new_n536));
  NAND2_X1  g0336(.A1(KEYINPUT22), .A2(G87), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT24), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n538), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n540), .A2(new_n531), .A3(new_n541), .A4(new_n534), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n525), .B1(new_n543), .B2(new_n257), .ZN(new_n544));
  INV_X1    g0344(.A(G257), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G1698), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G250), .B2(G1698), .ZN(new_n547));
  INV_X1    g0347(.A(G294), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n339), .A2(new_n547), .B1(new_n280), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n483), .A2(new_n478), .B1(new_n274), .B2(new_n276), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n549), .A2(new_n279), .B1(G264), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n390), .A3(new_n484), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n279), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(G264), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n553), .A2(new_n484), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n552), .B1(new_n555), .B2(G200), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n544), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n333), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n551), .A2(new_n484), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n319), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n407), .B1(new_n539), .B2(new_n542), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n558), .B(new_n560), .C1(new_n561), .C2(new_n525), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT89), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT89), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n557), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT84), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n438), .A2(G1698), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n336), .A2(new_n338), .A3(new_n281), .A4(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G250), .A2(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(KEYINPUT4), .A2(G244), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(G1698), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n368), .A2(new_n575), .B1(G33), .B2(G283), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n279), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n481), .A2(G257), .A3(new_n304), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n484), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT82), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n484), .A3(KEYINPUT82), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n578), .A2(new_n582), .A3(new_n333), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n278), .B1(new_n572), .B2(new_n576), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n319), .B1(new_n585), .B2(new_n580), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g0387(.A(G97), .B(G107), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT6), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G97), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n589), .A2(new_n591), .A3(G107), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n369), .A2(new_n371), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G107), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n407), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n251), .A2(G97), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n490), .B2(G97), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT83), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n592), .B1(new_n589), .B2(new_n588), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n603), .A2(new_n207), .B1(new_n265), .B2(new_n263), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n520), .B1(new_n369), .B2(new_n371), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n257), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT83), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n600), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n587), .B1(new_n602), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(G200), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n579), .A2(new_n484), .A3(KEYINPUT82), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT82), .B1(new_n579), .B2(new_n484), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n613), .B2(new_n578), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n606), .A2(new_n600), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n585), .A2(new_n390), .A3(new_n580), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n568), .B1(new_n609), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n615), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G200), .ZN(new_n621));
  INV_X1    g0421(.A(new_n616), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n606), .A2(new_n607), .A3(new_n600), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n607), .B1(new_n606), .B2(new_n600), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(KEYINPUT84), .B(new_n623), .C1(new_n626), .C2(new_n587), .ZN(new_n627));
  OR2_X1    g0427(.A1(KEYINPUT86), .A2(G87), .ZN(new_n628));
  NOR2_X1   g0428(.A1(G97), .A2(G107), .ZN(new_n629));
  NAND2_X1  g0429(.A1(KEYINPUT86), .A2(G87), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT19), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n288), .B2(new_n207), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n264), .B2(new_n591), .ZN(new_n635));
  INV_X1    g0435(.A(G68), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n634), .B(new_n635), .C1(new_n536), .C2(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n257), .B1(new_n255), .B2(new_n434), .ZN(new_n638));
  INV_X1    g0438(.A(new_n434), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n490), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n304), .A2(G274), .A3(new_n478), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n206), .A2(G45), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n304), .A2(G250), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n438), .A2(G1698), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(G238), .B2(G1698), .ZN(new_n647));
  INV_X1    g0447(.A(new_n496), .ZN(new_n648));
  NOR2_X1   g0448(.A1(KEYINPUT85), .A2(G116), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI22_X1  g0450(.A1(new_n339), .A2(new_n647), .B1(new_n650), .B2(new_n280), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n645), .B1(new_n651), .B2(new_n279), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n333), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n641), .B(new_n653), .C1(G169), .C2(new_n652), .ZN(new_n654));
  INV_X1    g0454(.A(new_n652), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G200), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n490), .A2(G87), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(G190), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n656), .A2(new_n638), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n618), .A2(new_n627), .A3(new_n660), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n471), .A2(new_n519), .A3(new_n567), .A4(new_n661), .ZN(G372));
  OAI21_X1  g0462(.A(new_n379), .B1(new_n319), .B2(new_n381), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n378), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g0464(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n378), .A2(new_n663), .A3(new_n665), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n331), .B1(new_n462), .B2(new_n453), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n400), .A2(KEYINPUT80), .A3(new_n401), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT80), .B1(new_n400), .B2(new_n401), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n669), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n427), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n429), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n471), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n654), .A2(new_n659), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n544), .B2(new_n556), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n609), .A2(new_n617), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n562), .B(new_n503), .C1(new_n508), .C2(new_n509), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  INV_X1    g0484(.A(new_n587), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n660), .A2(new_n684), .A3(new_n685), .A4(new_n615), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n625), .B2(new_n624), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT26), .B1(new_n687), .B2(new_n679), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n688), .A3(new_n654), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n677), .B1(new_n678), .B2(new_n690), .ZN(G369));
  NAND3_X1  g0491(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n567), .B1(new_n544), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n562), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n697), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n500), .A2(new_n697), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n517), .B2(new_n503), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n519), .B2(new_n704), .ZN(new_n706));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n517), .A2(new_n503), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n698), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n566), .B2(new_n564), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n697), .B(KEYINPUT91), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n700), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n709), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n210), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G1), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n631), .A2(G116), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n719), .A2(new_n720), .B1(new_n217), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n660), .A2(new_n684), .A3(new_n609), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n685), .A2(new_n615), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT26), .B1(new_n679), .B2(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n723), .A2(new_n725), .A3(new_n654), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n687), .A2(new_n727), .A3(new_n623), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT93), .B1(new_n609), .B2(new_n617), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n680), .A2(new_n728), .A3(new_n729), .A4(new_n682), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n697), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n713), .B1(new_n683), .B2(new_n689), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n477), .A2(new_n485), .A3(G179), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n585), .A2(new_n580), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n551), .A3(new_n739), .A4(new_n652), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n551), .A2(new_n652), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n477), .A2(new_n485), .A3(G179), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(new_n739), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n655), .A2(new_n486), .A3(new_n333), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n620), .A2(new_n559), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n741), .A2(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n749), .A2(new_n750), .A3(new_n713), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(new_n747), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n745), .B1(new_n744), .B2(new_n739), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT92), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n757), .A2(new_n758), .A3(new_n697), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n751), .B1(new_n759), .B2(new_n750), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n661), .A2(new_n519), .A3(new_n567), .A4(new_n713), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n707), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n737), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n722), .B1(new_n763), .B2(G1), .ZN(G364));
  AND2_X1   g0564(.A1(new_n207), .A2(G13), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n206), .B1(new_n765), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n717), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n213), .B1(G20), .B2(new_n319), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n333), .A2(new_n610), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT100), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n207), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G97), .ZN(new_n777));
  NAND3_X1  g0577(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n777), .B1(new_n636), .B2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT102), .Z(new_n782));
  NOR2_X1   g0582(.A1(new_n778), .A2(new_n390), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n202), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n207), .A2(new_n390), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n610), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n628), .B2(new_n630), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n207), .A2(G190), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n333), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n789), .B1(G77), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n790), .A2(new_n787), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n794), .B(new_n368), .C1(new_n520), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n786), .A2(new_n791), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT99), .Z(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n785), .B(new_n796), .C1(G58), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n773), .A2(new_n790), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT101), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT101), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OR3_X1    g0604(.A1(new_n804), .A2(KEYINPUT32), .A3(new_n362), .ZN(new_n805));
  OAI21_X1  g0605(.A(KEYINPUT32), .B1(new_n804), .B2(new_n362), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n782), .A2(new_n800), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n783), .A2(G326), .ZN(new_n808));
  INV_X1    g0608(.A(G322), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n808), .B(new_n370), .C1(new_n809), .C2(new_n797), .ZN(new_n810));
  INV_X1    g0610(.A(new_n788), .ZN(new_n811));
  INV_X1    g0611(.A(new_n795), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G303), .A2(new_n811), .B1(new_n812), .B2(G283), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n792), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n810), .B(new_n815), .C1(new_n779), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n804), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G329), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n817), .B(new_n819), .C1(new_n548), .C2(new_n775), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n771), .B1(new_n807), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G13), .A2(G33), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT95), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n207), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT96), .Z(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n770), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT97), .Z(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT98), .Z(new_n829));
  NOR2_X1   g0629(.A1(new_n716), .A2(new_n370), .ZN(new_n830));
  OR2_X1    g0630(.A1(G355), .A2(KEYINPUT94), .ZN(new_n831));
  NAND2_X1  g0631(.A1(G355), .A2(KEYINPUT94), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n243), .A2(G45), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n336), .A2(new_n338), .A3(new_n281), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n716), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(G45), .B2(new_n217), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n833), .B1(G116), .B2(new_n210), .C1(new_n834), .C2(new_n837), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n769), .B(new_n821), .C1(new_n829), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n706), .A2(new_n826), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n708), .A2(new_n768), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n706), .A2(new_n707), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G396));
  NOR2_X1   g0646(.A1(new_n770), .A2(new_n822), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n768), .B1(G77), .B2(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n793), .A2(G159), .B1(G137), .B2(new_n783), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n404), .B2(new_n780), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n799), .B2(G143), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n852), .A2(KEYINPUT34), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(KEYINPUT34), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n818), .A2(G132), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n835), .B1(new_n202), .B2(new_n788), .C1(new_n636), .C2(new_n795), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n776), .B2(G58), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n804), .A2(new_n814), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n520), .A2(new_n788), .B1(new_n797), .B2(new_n548), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n487), .B2(new_n793), .ZN(new_n861));
  INV_X1    g0661(.A(G87), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n370), .B1(new_n795), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(KEYINPUT103), .B(G283), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n780), .A2(new_n864), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n863), .B(new_n865), .C1(G303), .C2(new_n783), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n777), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n858), .B1(new_n859), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(new_n770), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n449), .B1(new_n437), .B2(new_n698), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n453), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n453), .A2(new_n697), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n849), .B(new_n869), .C1(new_n823), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n870), .B2(new_n453), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n733), .B(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n762), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n768), .B1(new_n878), .B2(new_n879), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n875), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(G384));
  NOR2_X1   g0684(.A1(new_n765), .A2(new_n206), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n759), .A2(new_n750), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n757), .A2(new_n758), .A3(KEYINPUT31), .A4(new_n697), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n761), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n471), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT104), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n359), .A2(new_n257), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT7), .B1(new_n835), .B2(G20), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(G68), .A3(new_n356), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT16), .B1(new_n894), .B2(new_n354), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n377), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n695), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n673), .B2(new_n387), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n663), .A2(KEYINPUT79), .B1(new_n374), .B2(new_n377), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT37), .B1(new_n900), .B2(new_n382), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n392), .A2(new_n374), .A3(new_n377), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n378), .A2(new_n897), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n896), .A2(new_n663), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n902), .A2(new_n898), .A3(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n901), .A2(new_n904), .B1(new_n906), .B2(KEYINPUT37), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n891), .B1(new_n899), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n387), .A2(new_n399), .A3(new_n402), .ZN(new_n909));
  INV_X1    g0709(.A(new_n898), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n461), .A2(new_n697), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n462), .A2(new_n330), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n461), .B(new_n697), .C1(new_n460), .C2(new_n331), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n874), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n888), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT40), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n667), .A2(new_n400), .A3(new_n401), .A4(new_n668), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(new_n378), .A3(new_n897), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n902), .A2(new_n903), .ZN(new_n922));
  INV_X1    g0722(.A(new_n664), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT37), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT37), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n383), .A2(new_n925), .A3(new_n902), .A4(new_n903), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n921), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n912), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n888), .A2(KEYINPUT40), .A3(new_n917), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n919), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n707), .B1(new_n890), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n890), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n891), .B(new_n907), .C1(new_n909), .C2(new_n910), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n936), .B2(new_n928), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n908), .A2(new_n912), .A3(KEYINPUT39), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n462), .A2(new_n697), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n897), .B1(new_n667), .B2(new_n668), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n915), .A2(new_n916), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n713), .B(new_n876), .C1(new_n683), .C2(new_n689), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(new_n873), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n941), .B1(new_n913), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n676), .B1(new_n471), .B2(new_n737), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n885), .B1(new_n934), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n934), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n594), .A2(KEYINPUT35), .ZN(new_n952));
  INV_X1    g0752(.A(G116), .ZN(new_n953));
  NOR4_X1   g0753(.A1(new_n951), .A2(new_n952), .A3(new_n215), .A4(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT36), .ZN(new_n955));
  INV_X1    g0755(.A(new_n217), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n956), .B(G77), .C1(new_n240), .C2(new_n220), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n202), .A2(G68), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n206), .B(G13), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n950), .A2(new_n960), .ZN(G367));
  NAND2_X1  g0761(.A1(new_n728), .A2(new_n729), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n619), .B2(new_n713), .ZN(new_n963));
  INV_X1    g0763(.A(new_n713), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n587), .A3(new_n615), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n709), .A2(KEYINPUT105), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT105), .B1(new_n709), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n638), .A2(new_n657), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n697), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n660), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n654), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n970), .B1(KEYINPUT43), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n968), .A2(new_n976), .A3(new_n969), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n966), .A2(new_n712), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT42), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n609), .B1(new_n966), .B2(new_n700), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n964), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n978), .A2(new_n984), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n717), .B(KEYINPUT41), .Z(new_n987));
  AOI21_X1  g0787(.A(new_n712), .B1(new_n702), .B2(new_n711), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(new_n708), .Z(new_n989));
  AND2_X1   g0789(.A1(new_n989), .A2(new_n763), .ZN(new_n990));
  INV_X1    g0790(.A(new_n709), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n714), .A2(new_n966), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT45), .ZN(new_n993));
  XOR2_X1   g0793(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OR3_X1    g0795(.A1(new_n714), .A2(new_n966), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n714), .B2(new_n966), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n991), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n992), .B(new_n1000), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n1001), .A2(new_n709), .A3(new_n996), .A4(new_n997), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n990), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n987), .B1(new_n1003), .B2(new_n763), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n985), .B(new_n986), .C1(new_n1004), .C2(new_n767), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n836), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n1006), .A2(new_n237), .B1(new_n210), .B2(new_n434), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n828), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT107), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n768), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n1009), .B2(new_n1008), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n370), .B1(new_n812), .B2(G77), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n362), .B2(new_n780), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G58), .A2(new_n811), .B1(new_n793), .B2(G50), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n404), .B2(new_n797), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G143), .C2(new_n783), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n776), .A2(G68), .ZN(new_n1017));
  INV_X1    g0817(.A(G137), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1017), .C1(new_n1018), .C2(new_n804), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT108), .Z(new_n1020));
  NOR2_X1   g0820(.A1(new_n795), .A2(new_n591), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n811), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n792), .B2(new_n864), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(new_n799), .C2(G303), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n339), .B1(new_n780), .B2(new_n548), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT46), .B1(new_n811), .B2(new_n487), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(G311), .C2(new_n783), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(G317), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1028), .B1(new_n520), .B2(new_n775), .C1(new_n1029), .C2(new_n804), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1020), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT47), .Z(new_n1032));
  OAI221_X1 g0832(.A(new_n1011), .B1(new_n825), .B2(new_n974), .C1(new_n1032), .C2(new_n771), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1005), .A2(new_n1033), .ZN(G387));
  NOR2_X1   g0834(.A1(new_n990), .A2(new_n718), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n763), .B2(new_n989), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n989), .A2(new_n767), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n818), .A2(G150), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n776), .A2(new_n639), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n788), .A2(new_n265), .B1(new_n792), .B2(new_n636), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n797), .A2(new_n202), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n1040), .A2(new_n1021), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n835), .B1(new_n780), .B2(new_n375), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G159), .B2(new_n783), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1038), .A2(new_n1039), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n793), .A2(G303), .B1(G311), .B2(new_n779), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n809), .B2(new_n784), .C1(new_n798), .C2(new_n1029), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n775), .A2(new_n864), .B1(new_n548), .B2(new_n788), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT109), .Z(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n339), .B1(new_n650), .B2(new_n795), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n818), .B2(G326), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1045), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n770), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n830), .A2(new_n720), .B1(new_n520), .B2(new_n716), .ZN(new_n1061));
  AOI211_X1 g0861(.A(G45), .B(new_n720), .C1(G68), .C2(G77), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT50), .B1(new_n432), .B2(new_n202), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n432), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n836), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n234), .A2(new_n293), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1061), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n769), .B1(new_n829), .B2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1060), .B(new_n1069), .C1(new_n703), .C2(new_n825), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1036), .A2(new_n1037), .A3(new_n1070), .ZN(G393));
  INV_X1    g0871(.A(KEYINPUT110), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n999), .A2(new_n1002), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n999), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n717), .B(new_n1003), .C1(new_n1074), .C2(new_n990), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n818), .A2(G143), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n776), .A2(G77), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n375), .A2(new_n792), .B1(new_n795), .B2(new_n862), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n835), .B1(new_n780), .B2(new_n202), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n250), .C2(new_n811), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n784), .A2(new_n404), .B1(new_n797), .B2(new_n362), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1076), .A2(new_n1077), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n818), .A2(G322), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n784), .A2(new_n1029), .B1(new_n797), .B2(new_n814), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n776), .A2(new_n487), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n370), .B1(new_n795), .B2(new_n520), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n788), .A2(new_n864), .B1(new_n792), .B2(new_n548), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G303), .C2(new_n779), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .A4(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1083), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n836), .A2(new_n246), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n591), .B2(new_n210), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n768), .B1(new_n1093), .B2(new_n771), .C1(new_n828), .C2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n967), .B2(new_n826), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1074), .B2(new_n767), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1075), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT112), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT112), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1075), .A2(new_n1101), .A3(new_n1098), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(G390));
  NAND2_X1  g0903(.A1(new_n762), .A2(new_n917), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT113), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT113), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n762), .A2(new_n1106), .A3(new_n917), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n939), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n872), .B1(new_n731), .B2(new_n871), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n930), .B(new_n1109), .C1(new_n942), .C2(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n937), .A2(new_n938), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n943), .A2(new_n873), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n915), .A2(new_n916), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n939), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1108), .B(new_n1111), .C1(new_n1112), .C2(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n888), .A2(G330), .A3(new_n917), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1115), .B1(new_n937), .B2(new_n938), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1109), .B1(new_n1110), .B2(new_n942), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n928), .B1(new_n911), .B2(KEYINPUT38), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1117), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1116), .A2(new_n767), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1112), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n823), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n370), .B1(new_n795), .B2(new_n636), .C1(new_n780), .C2(new_n520), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n793), .A2(G97), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n862), .B2(new_n788), .C1(new_n953), .C2(new_n797), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(G283), .C2(new_n783), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1129), .B(new_n1077), .C1(new_n548), .C2(new_n804), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n818), .A2(G125), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n811), .A2(G150), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n780), .A2(new_n1018), .B1(new_n784), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n368), .B1(new_n792), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(G132), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n797), .A2(new_n1138), .B1(new_n795), .B2(new_n202), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n1133), .A2(new_n1135), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1131), .B(new_n1140), .C1(new_n362), .C2(new_n775), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n771), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n769), .B(new_n1142), .C1(new_n375), .C2(new_n847), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1125), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1123), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n888), .A2(G330), .A3(new_n876), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n942), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n762), .A2(new_n1106), .A3(new_n917), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1106), .B1(new_n762), .B2(new_n917), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1110), .B(new_n1148), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1114), .B1(new_n762), .B2(new_n876), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1113), .B1(new_n1152), .B2(new_n1117), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n736), .B1(new_n465), .B2(new_n470), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n888), .A2(G330), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n465), .B2(new_n470), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1155), .A2(new_n1157), .A3(new_n676), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1116), .A2(new_n1122), .A3(new_n1154), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT114), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n717), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1160), .B1(new_n1159), .B2(new_n717), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1146), .B1(new_n1165), .B2(new_n1166), .ZN(G378));
  NOR4_X1   g0967(.A1(new_n1155), .A2(new_n1157), .A3(KEYINPUT118), .A4(new_n676), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT118), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1157), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n947), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1159), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n940), .A2(new_n945), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n427), .A2(new_n429), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n411), .A2(new_n695), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1175), .B(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1177), .B(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT40), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n909), .A2(new_n910), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n907), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT38), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n936), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n888), .A2(new_n917), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1181), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n707), .B1(new_n931), .B2(new_n930), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1180), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n888), .A2(KEYINPUT40), .A3(new_n917), .ZN(new_n1190));
  OAI21_X1  g0990(.A(G330), .B1(new_n1190), .B2(new_n1120), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1177), .B(new_n1178), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n919), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1174), .B1(new_n1189), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n919), .B2(new_n1191), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1187), .A2(new_n1188), .A3(new_n1180), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n946), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1173), .A2(new_n1198), .A3(KEYINPUT57), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1159), .A2(new_n1172), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n717), .C1(KEYINPUT57), .C2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n766), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1192), .A2(new_n823), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n768), .B1(G50), .B2(new_n848), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n339), .A2(new_n292), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n280), .A2(new_n292), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT115), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1207), .A3(new_n202), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT116), .Z(new_n1209));
  OAI22_X1  g1009(.A1(new_n780), .A2(new_n591), .B1(new_n784), .B2(new_n953), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n788), .A2(new_n265), .B1(new_n792), .B2(new_n434), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n797), .A2(new_n520), .B1(new_n795), .B2(new_n240), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1205), .ZN(new_n1213));
  INV_X1    g1013(.A(G283), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1017), .B(new_n1213), .C1(new_n1214), .C2(new_n804), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1209), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1134), .A2(new_n797), .B1(new_n788), .B2(new_n1136), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G137), .B2(new_n793), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n779), .A2(G132), .B1(new_n783), .B2(G125), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n775), .C2(new_n404), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n818), .A2(G124), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1207), .B1(G159), .B2(new_n812), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1217), .B1(new_n1216), .B2(new_n1215), .C1(new_n1222), .C2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1204), .B1(new_n1227), .B2(new_n770), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1203), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT117), .B1(new_n1202), .B2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n946), .A2(new_n1196), .A3(new_n1195), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1195), .A2(new_n1196), .B1(new_n940), .B2(new_n945), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n767), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT117), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1229), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1231), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1201), .A2(new_n1237), .ZN(G375));
  AOI21_X1  g1038(.A(new_n769), .B1(new_n636), .B2(new_n847), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n804), .A2(new_n475), .B1(new_n591), .B2(new_n788), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT120), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n370), .B1(new_n795), .B2(new_n265), .C1(new_n1214), .C2(new_n797), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G294), .B2(new_n783), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n780), .A2(new_n650), .B1(new_n792), .B2(new_n520), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT119), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1039), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n775), .A2(new_n202), .B1(new_n404), .B2(new_n792), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT121), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n835), .B1(new_n240), .B2(new_n795), .C1(new_n362), .C2(new_n788), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n1138), .A2(new_n784), .B1(new_n780), .B2(new_n1136), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n799), .C2(G137), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1134), .B2(new_n804), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1241), .A2(new_n1246), .B1(new_n1248), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT122), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n770), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n822), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1239), .B1(new_n1255), .B2(new_n1257), .C1(new_n1114), .C2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1154), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1259), .B1(new_n1260), .B2(new_n766), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1163), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(new_n987), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1262), .B1(new_n1264), .B2(new_n1265), .ZN(G381));
  OR4_X1    g1066(.A1(G396), .A2(G387), .A3(G384), .A4(G393), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1173), .A2(new_n1198), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT57), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1269), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n718), .B1(new_n1271), .B2(new_n1173), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1270), .A2(new_n1272), .B1(new_n1231), .B2(new_n1236), .ZN(new_n1273));
  INV_X1    g1073(.A(G378), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G390), .A2(new_n1267), .A3(G381), .A4(new_n1275), .ZN(G407));
  NAND2_X1  g1076(.A1(new_n696), .A2(G213), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT123), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G407), .B(G213), .C1(new_n1275), .C2(new_n1279), .ZN(G409));
  AOI21_X1  g1080(.A(new_n1230), .B1(new_n1198), .B2(new_n767), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1281), .A2(KEYINPUT125), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(KEYINPUT125), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1268), .A2(new_n987), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1274), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT124), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1273), .B2(G378), .ZN(new_n1288));
  AND4_X1   g1088(.A1(new_n1287), .A2(new_n1201), .A3(new_n1237), .A4(G378), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1286), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1163), .A2(KEYINPUT60), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1265), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n717), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1262), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n883), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(G384), .A3(new_n1262), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1290), .A2(new_n1279), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT62), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1290), .A2(new_n1303), .A3(new_n1279), .A4(new_n1300), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1278), .A2(G2897), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1299), .A2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1297), .A2(G2897), .A3(new_n1278), .A4(new_n1298), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT124), .B1(G375), .B2(new_n1274), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1273), .A2(new_n1287), .A3(G378), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1309), .A2(new_n1310), .B1(new_n1274), .B2(new_n1285), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1308), .B1(new_n1311), .B2(new_n1278), .ZN(new_n1312));
  XOR2_X1   g1112(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1313));
  NAND4_X1  g1113(.A1(new_n1302), .A2(new_n1304), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(G393), .B(new_n845), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  AND3_X1   g1116(.A1(G387), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G387), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1316), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(G387), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G390), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(G387), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(new_n1315), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1314), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT61), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1319), .A2(new_n1326), .A3(new_n1323), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1327), .B1(new_n1328), .B2(new_n1301), .ZN(new_n1329));
  OAI21_X1  g1129(.A(KEYINPUT126), .B1(new_n1311), .B2(new_n1278), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1290), .A2(new_n1331), .A3(new_n1279), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1330), .A2(new_n1308), .A3(new_n1332), .ZN(new_n1333));
  OR2_X1    g1133(.A1(new_n1301), .A2(new_n1328), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1329), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1325), .A2(new_n1335), .ZN(G405));
  NOR2_X1   g1136(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1273), .A2(G378), .ZN(new_n1338));
  OR3_X1    g1138(.A1(new_n1337), .A2(new_n1300), .A3(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1300), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1341), .B(new_n1324), .ZN(G402));
endmodule


