//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1161, new_n1162, new_n1163, new_n1165,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NAND2_X1  g0003(.A1(G68), .A2(G238), .ZN(new_n204));
  INV_X1    g0004(.A(G50), .ZN(new_n205));
  INV_X1    g0005(.A(G226), .ZN(new_n206));
  OAI21_X1  g0006(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  AOI211_X1 g0009(.A(new_n207), .B(new_n209), .C1(G77), .C2(G244), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G116), .A2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n203), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n203), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  NOR2_X1   g0023(.A1(G58), .A2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR4_X1   g0029(.A1(new_n219), .A2(new_n220), .A3(new_n223), .A4(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n216), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n206), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n213), .A2(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G97), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n252), .A2(new_n256), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n228), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT67), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(new_n259), .B2(new_n228), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(KEYINPUT67), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n262), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n264), .A2(new_n267), .ZN(new_n273));
  INV_X1    g0073(.A(new_n271), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(G238), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n261), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n261), .A2(new_n272), .A3(new_n278), .A4(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G200), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT73), .B1(new_n283), .B2(new_n205), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n227), .A2(G33), .A3(G77), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT73), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n282), .A2(new_n286), .A3(G50), .ZN(new_n287));
  INV_X1    g0087(.A(G68), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G20), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n284), .A2(new_n285), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n228), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT68), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(KEYINPUT68), .A3(new_n228), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n290), .A2(KEYINPUT11), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n227), .A2(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G13), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G68), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT12), .ZN(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT11), .B1(new_n290), .B2(new_n296), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n296), .A2(new_n288), .A3(new_n298), .ZN(new_n303));
  NOR4_X1   g0103(.A1(new_n297), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n277), .A2(G190), .A3(new_n279), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n281), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT74), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT75), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT14), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n280), .B2(G169), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  AOI211_X1 g0113(.A(new_n313), .B(new_n310), .C1(new_n277), .C2(new_n279), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n280), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G179), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n304), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT17), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n259), .A2(new_n263), .A3(new_n228), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT67), .B1(new_n265), .B2(new_n266), .ZN(new_n322));
  OAI211_X1 g0122(.A(G232), .B(new_n274), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT78), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT78), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n273), .A2(new_n325), .A3(G232), .A4(new_n274), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n324), .A2(new_n272), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n260), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT76), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n248), .B2(G33), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n250), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n206), .A2(G1698), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n334), .C1(G223), .C2(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G87), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n328), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(G200), .B1(new_n327), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n324), .A2(new_n272), .A3(new_n326), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT79), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n324), .A2(KEYINPUT79), .A3(new_n326), .A4(new_n272), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n337), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT16), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n252), .A2(new_n227), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n288), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(G58), .B(G68), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(G20), .B1(G159), .B2(new_n282), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n347), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n333), .B2(G20), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n331), .A2(new_n332), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n249), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n227), .ZN(new_n361));
  OR2_X1    g0161(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n358), .B(G68), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n354), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n296), .B(new_n356), .C1(new_n364), .C2(new_n347), .ZN(new_n365));
  INV_X1    g0165(.A(new_n296), .ZN(new_n366));
  INV_X1    g0166(.A(new_n298), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT69), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G58), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT8), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n370), .B(new_n371), .ZN(new_n372));
  MUX2_X1   g0172(.A(new_n368), .B(new_n299), .S(new_n372), .Z(new_n373));
  NAND2_X1  g0173(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n320), .B1(new_n346), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n374), .ZN(new_n376));
  AOI211_X1 g0176(.A(G190), .B(new_n337), .C1(new_n342), .C2(new_n343), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n376), .B(KEYINPUT17), .C1(new_n377), .C2(new_n339), .ZN(new_n378));
  INV_X1    g0178(.A(G179), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n344), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(G169), .B1(new_n327), .B2(new_n338), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AND4_X1   g0182(.A1(KEYINPUT18), .A2(new_n380), .A3(new_n374), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n381), .B1(new_n344), .B2(new_n379), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT18), .B1(new_n384), .B2(new_n374), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n375), .B(new_n378), .C1(new_n383), .C2(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n319), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n225), .B2(G50), .ZN(new_n388));
  INV_X1    g0188(.A(G150), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n227), .A2(G33), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n388), .B1(new_n389), .B2(new_n283), .C1(new_n372), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n299), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n391), .A2(new_n296), .B1(new_n205), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n367), .A2(G50), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT70), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(new_n366), .A3(new_n299), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT9), .ZN(new_n398));
  INV_X1    g0198(.A(new_n252), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n253), .A2(G222), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G223), .A2(G1698), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n260), .C1(G77), .C2(new_n399), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n273), .A2(G226), .A3(new_n274), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n272), .A3(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n397), .A2(new_n398), .B1(G200), .B2(new_n405), .ZN(new_n406));
  OAI221_X1 g0206(.A(new_n406), .B1(new_n398), .B2(new_n397), .C1(new_n345), .C2(new_n405), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT10), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n405), .A2(G179), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n313), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n397), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n273), .A2(G244), .A3(new_n274), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n253), .A2(G232), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G238), .A2(G1698), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n249), .A2(new_n251), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n260), .C1(new_n399), .C2(G107), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n272), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT71), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT71), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n272), .A2(new_n413), .A3(new_n417), .A4(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(G200), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n366), .A2(G77), .A3(new_n367), .ZN(new_n423));
  INV_X1    g0223(.A(G77), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n392), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT8), .B(G58), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n426), .A2(new_n283), .B1(new_n227), .B2(new_n424), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT15), .B(G87), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n390), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n296), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n423), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n422), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT72), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n419), .A2(new_n421), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G190), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n422), .A2(KEYINPUT72), .A3(new_n432), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n379), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n419), .A2(new_n313), .A3(new_n421), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n431), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n387), .A2(new_n412), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G250), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n253), .ZN(new_n446));
  INV_X1    g0246(.A(G257), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G1698), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n359), .A2(new_n249), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G294), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT86), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT86), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(new_n453), .A3(new_n450), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n260), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G41), .ZN(new_n458));
  INV_X1    g0258(.A(G1), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(KEYINPUT82), .A3(new_n459), .A4(G45), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT82), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(G45), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n268), .A2(new_n456), .A3(new_n460), .A4(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n456), .A3(new_n460), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G264), .A3(new_n273), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n455), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G200), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n359), .A2(KEYINPUT22), .A3(G87), .A4(new_n249), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G116), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n227), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT85), .B1(new_n215), .B2(G20), .ZN(new_n474));
  XOR2_X1   g0274(.A(new_n474), .B(KEYINPUT23), .Z(new_n475));
  INV_X1    g0275(.A(G87), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n252), .A2(G20), .A3(new_n476), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n477), .A2(KEYINPUT22), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT24), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n473), .A2(KEYINPUT24), .A3(new_n475), .A4(new_n478), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n296), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n459), .A2(KEYINPUT80), .A3(G33), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n294), .A2(new_n299), .A3(new_n295), .A4(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT80), .B1(new_n459), .B2(G33), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n487), .A2(new_n215), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n299), .A2(G107), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT25), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n483), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n468), .A2(new_n345), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n455), .A2(new_n465), .A3(new_n467), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT87), .B1(new_n494), .B2(new_n313), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(G179), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT87), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n468), .A2(new_n497), .A3(G169), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n469), .A2(new_n493), .B1(new_n499), .B2(new_n491), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n227), .C1(G33), .C2(new_n257), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n502), .B(new_n292), .C1(new_n227), .C2(G116), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT20), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G116), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n392), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n505), .B(new_n507), .C1(new_n487), .C2(new_n506), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n447), .A2(new_n253), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n216), .A2(G1698), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n359), .A2(new_n249), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n252), .A2(G303), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n260), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n466), .A2(G270), .A3(new_n273), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n465), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n508), .A2(G169), .A3(new_n516), .ZN(new_n517));
  XOR2_X1   g0317(.A(KEYINPUT84), .B(KEYINPUT21), .Z(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT21), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT84), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n508), .A2(G169), .A3(new_n521), .A4(new_n516), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n516), .A2(new_n379), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n508), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n519), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n516), .A2(G200), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n345), .B2(new_n516), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n527), .A2(new_n508), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n333), .A2(G244), .A3(new_n253), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n253), .A2(KEYINPUT4), .A3(G244), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n445), .B2(new_n253), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n399), .A2(new_n534), .B1(G33), .B2(G283), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n328), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n466), .A2(G257), .A3(new_n273), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n465), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n313), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n532), .A2(new_n535), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n260), .ZN(new_n541));
  INV_X1    g0341(.A(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n539), .B1(new_n543), .B2(G179), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n350), .A2(new_n351), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G107), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n215), .A2(KEYINPUT6), .A3(G97), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n257), .A2(new_n215), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n550), .B2(KEYINPUT6), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(G20), .B1(G77), .B2(new_n282), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n366), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(G97), .B1(new_n485), .B2(new_n486), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n299), .A2(new_n257), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT81), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(KEYINPUT81), .A3(new_n555), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n544), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n543), .A2(G200), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n560), .B(new_n562), .C1(new_n345), .C2(new_n543), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  MUX2_X1   g0364(.A(G238), .B(G244), .S(G1698), .Z(new_n565));
  AOI22_X1  g0365(.A1(new_n333), .A2(new_n565), .B1(G33), .B2(G116), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n566), .A2(new_n328), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n463), .A2(new_n445), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n273), .B(new_n568), .C1(G274), .C2(new_n463), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n379), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n566), .B2(new_n328), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n313), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n333), .A2(new_n227), .A3(G68), .ZN(new_n573));
  NAND3_X1  g0373(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n574), .A2(new_n227), .ZN(new_n575));
  NOR3_X1   g0375(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT83), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n390), .B2(new_n257), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n227), .A2(new_n574), .B1(new_n549), .B2(new_n476), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT83), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n573), .A2(new_n577), .A3(new_n579), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n296), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n392), .A2(new_n428), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n487), .A2(new_n428), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n570), .B(new_n572), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n487), .A2(new_n476), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n567), .A2(G190), .A3(new_n569), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n571), .A2(G200), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n583), .A2(new_n296), .B1(new_n392), .B2(new_n428), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n564), .A2(new_n594), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n444), .A2(new_n500), .A3(new_n529), .A4(new_n595), .ZN(G372));
  NAND2_X1  g0396(.A1(new_n499), .A2(new_n491), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n525), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n493), .A2(new_n469), .ZN(new_n599));
  INV_X1    g0399(.A(new_n564), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n593), .A4(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n594), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n544), .A2(new_n560), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT26), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT26), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(KEYINPUT88), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT88), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n602), .A2(new_n603), .A3(new_n607), .A4(KEYINPUT26), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n601), .A2(new_n609), .A3(new_n588), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n444), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n411), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n378), .A2(new_n375), .ZN(new_n613));
  INV_X1    g0413(.A(new_n306), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n442), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n318), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT89), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n383), .B2(new_n385), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n380), .A2(new_n374), .A3(new_n382), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT18), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n384), .A2(KEYINPUT18), .A3(new_n374), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(KEYINPUT89), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n612), .B1(new_n625), .B2(new_n408), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n611), .A2(new_n626), .ZN(G369));
  INV_X1    g0427(.A(G13), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n628), .A2(G20), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n459), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(G213), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G343), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n508), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n636), .B(KEYINPUT90), .Z(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n525), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n529), .B2(new_n637), .ZN(new_n639));
  INV_X1    g0439(.A(G330), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n599), .A2(new_n597), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n491), .A2(new_n635), .ZN(new_n643));
  INV_X1    g0443(.A(new_n635), .ZN(new_n644));
  OAI22_X1  g0444(.A1(new_n642), .A2(new_n643), .B1(new_n597), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT91), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n525), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n644), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n642), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n635), .B(KEYINPUT92), .Z(new_n652));
  NOR2_X1   g0452(.A1(new_n597), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n648), .A2(new_n654), .ZN(G399));
  INV_X1    g0455(.A(new_n221), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G41), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G1), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n576), .A2(new_n506), .ZN(new_n660));
  OAI22_X1  g0460(.A1(new_n659), .A2(new_n660), .B1(new_n226), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT28), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT31), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n514), .A2(new_n465), .A3(new_n515), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n664), .A2(G179), .A3(new_n467), .A4(new_n455), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n541), .A2(new_n542), .A3(new_n567), .A4(new_n569), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT30), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n455), .A2(new_n467), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n536), .A2(new_n571), .A3(new_n538), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT30), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n668), .A2(new_n669), .A3(new_n523), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n516), .B(new_n379), .C1(new_n536), .C2(new_n538), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n494), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n571), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT93), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n667), .A2(new_n671), .B1(new_n674), .B2(new_n571), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n635), .B1(new_n679), .B2(KEYINPUT93), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n663), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n652), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n500), .A2(new_n595), .A3(new_n529), .A4(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n676), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n610), .A2(new_n682), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n604), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n601), .B(new_n588), .C1(new_n690), .C2(new_n605), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(KEYINPUT29), .A3(new_n644), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n686), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n662), .B1(new_n693), .B2(G1), .ZN(G364));
  NOR2_X1   g0494(.A1(new_n227), .A2(G190), .ZN(new_n695));
  INV_X1    g0495(.A(G200), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(new_n379), .A3(new_n696), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT95), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT95), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G159), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT32), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n227), .A2(new_n345), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n696), .A2(G179), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G87), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n695), .A2(G179), .A3(new_n696), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G77), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(G179), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G200), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n695), .A2(G179), .A3(G200), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n714), .A2(new_n212), .B1(new_n288), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n712), .A2(new_n696), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n399), .B1(new_n718), .B2(new_n205), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n345), .A2(G179), .A3(G200), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n227), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n257), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n705), .A2(new_n695), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n215), .ZN(new_n724));
  NOR4_X1   g0524(.A1(new_n716), .A2(new_n719), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n703), .A2(new_n708), .A3(new_n711), .A4(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n700), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n727), .A2(KEYINPUT98), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(KEYINPUT98), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n723), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n731), .A2(G329), .B1(G283), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT99), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n717), .B(KEYINPUT96), .Z(new_n735));
  INV_X1    g0535(.A(new_n721), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n735), .A2(G326), .B1(G294), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT97), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  XOR2_X1   g0539(.A(KEYINPUT33), .B(G317), .Z(new_n740));
  OAI221_X1 g0540(.A(new_n252), .B1(new_n709), .B2(new_n739), .C1(new_n715), .C2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n734), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G322), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n743), .B2(new_n714), .ZN(new_n744));
  INV_X1    g0544(.A(G303), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n706), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n726), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n228), .B1(G20), .B2(new_n313), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(G355), .B(KEYINPUT94), .Z(new_n750));
  NOR2_X1   g0550(.A1(new_n656), .A2(new_n252), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n243), .A2(new_n270), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n333), .A2(new_n656), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G45), .B2(new_n226), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n752), .B1(G116), .B2(new_n221), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n748), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n659), .B1(G45), .B2(new_n629), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n639), .A2(new_n759), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n749), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n641), .ZN(new_n765));
  INV_X1    g0565(.A(new_n762), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n639), .A2(new_n640), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n764), .A2(new_n768), .ZN(G396));
  AND2_X1   g0569(.A1(new_n440), .A2(new_n441), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n431), .A3(new_n635), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT101), .Z(new_n772));
  NAND2_X1  g0572(.A1(new_n431), .A2(new_n635), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n439), .A2(new_n442), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT100), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT100), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n439), .A2(new_n776), .A3(new_n442), .A4(new_n773), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n687), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n610), .A2(new_n682), .A3(new_n779), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(new_n686), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n766), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n757), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n748), .A2(new_n757), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n424), .ZN(new_n788));
  INV_X1    g0588(.A(new_n715), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n713), .A2(G143), .B1(new_n789), .B2(G150), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n717), .A2(G137), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n790), .B(new_n791), .C1(new_n701), .C2(new_n709), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT34), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n360), .B1(new_n731), .B2(G132), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n723), .A2(new_n288), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(new_n792), .B2(new_n793), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n795), .B(new_n797), .C1(new_n212), .C2(new_n721), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n794), .B(new_n798), .C1(G50), .C2(new_n707), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n718), .A2(new_n745), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n722), .B1(new_n731), .B2(G311), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n252), .B1(new_n706), .B2(new_n215), .C1(new_n506), .C2(new_n709), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G87), .B2(new_n732), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n801), .B(new_n803), .C1(new_n804), .C2(new_n715), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n800), .B(new_n805), .C1(G294), .C2(new_n713), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n748), .B1(new_n799), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n786), .A2(new_n762), .A3(new_n788), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n785), .A2(new_n808), .ZN(G384));
  INV_X1    g0609(.A(KEYINPUT38), .ZN(new_n810));
  INV_X1    g0610(.A(new_n633), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n374), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n624), .B2(new_n613), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n376), .B1(new_n339), .B2(new_n377), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n814), .A2(new_n812), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n815), .A2(new_n617), .A3(KEYINPUT37), .A4(new_n619), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n812), .B(KEYINPUT89), .C1(new_n346), .C2(new_n374), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT37), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n814), .A2(new_n619), .A3(new_n812), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n810), .B1(new_n813), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n364), .A2(KEYINPUT103), .A3(new_n347), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n347), .A2(KEYINPUT103), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n363), .A2(new_n354), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n823), .A2(new_n296), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n373), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n384), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n814), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n633), .B1(new_n826), .B2(new_n373), .ZN(new_n830));
  OAI21_X1  g0630(.A(KEYINPUT37), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(KEYINPUT37), .B2(new_n819), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n386), .A2(KEYINPUT104), .A3(new_n830), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT104), .B1(new_n386), .B2(new_n830), .ZN(new_n834));
  OAI211_X1 g0634(.A(KEYINPUT38), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n822), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n644), .B1(new_n676), .B2(new_n677), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n679), .A2(KEYINPUT93), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n837), .A2(KEYINPUT31), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n681), .A2(new_n839), .A3(new_n683), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n304), .A2(new_n644), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n307), .B2(new_n318), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n614), .A2(new_n841), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n315), .A2(new_n317), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(new_n304), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n772), .A2(new_n778), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n836), .A2(KEYINPUT40), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n810), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n850), .A2(KEYINPUT105), .A3(new_n835), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT105), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n849), .A2(new_n852), .A3(new_n810), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n848), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n444), .A2(new_n840), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n856), .B(new_n857), .Z(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(G330), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n318), .A2(new_n644), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n851), .A2(KEYINPUT39), .A3(new_n853), .ZN(new_n861));
  XNOR2_X1  g0661(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n822), .A2(new_n835), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n860), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n851), .A2(new_n853), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n770), .A2(new_n431), .A3(new_n644), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n782), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n842), .A2(new_n845), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n865), .A2(new_n869), .B1(new_n624), .B2(new_n811), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n689), .A2(new_n444), .A3(new_n692), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n626), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n871), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n859), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n459), .B2(new_n629), .ZN(new_n876));
  OAI211_X1 g0676(.A(G20), .B(new_n265), .C1(new_n551), .C2(KEYINPUT35), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n506), .B(new_n877), .C1(KEYINPUT35), .C2(new_n551), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT36), .Z(new_n879));
  OAI21_X1  g0679(.A(G77), .B1(new_n212), .B2(new_n288), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n226), .A2(new_n880), .B1(G50), .B2(new_n288), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G1), .A3(new_n628), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT102), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n876), .A2(new_n879), .A3(new_n883), .ZN(G367));
  NAND2_X1  g0684(.A1(new_n589), .A2(new_n592), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n635), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n602), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n588), .B2(new_n886), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT43), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n600), .B1(new_n560), .B2(new_n682), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n561), .B2(new_n682), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n651), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT42), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n561), .B1(new_n890), .B2(new_n597), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(new_n682), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n889), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n647), .A2(new_n891), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n888), .A2(KEYINPUT43), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  XNOR2_X1  g0701(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n657), .B(new_n902), .Z(new_n903));
  MUX2_X1   g0703(.A(new_n642), .B(new_n645), .S(new_n650), .Z(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(new_n765), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n693), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n648), .A2(KEYINPUT110), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n654), .A2(new_n891), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT45), .Z(new_n910));
  NOR2_X1   g0710(.A1(new_n654), .A2(new_n891), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT44), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n912), .A2(KEYINPUT109), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(KEYINPUT109), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n647), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n907), .B1(new_n908), .B2(new_n917), .C1(new_n918), .C2(KEYINPUT110), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n903), .B1(new_n919), .B2(new_n693), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n459), .B1(new_n629), .B2(G45), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n900), .B(new_n901), .C1(new_n920), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n735), .A2(G143), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n727), .A2(G137), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n723), .A2(new_n424), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n252), .B(new_n926), .C1(G159), .C2(new_n789), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n714), .A2(new_n389), .B1(new_n212), .B2(new_n706), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n721), .A2(new_n288), .B1(new_n709), .B2(new_n205), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n924), .A2(new_n925), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n360), .B1(new_n714), .B2(new_n745), .ZN(new_n932));
  INV_X1    g0732(.A(G317), .ZN(new_n933));
  INV_X1    g0733(.A(G294), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n700), .A2(new_n933), .B1(new_n934), .B2(new_n715), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n932), .B(new_n935), .C1(G283), .C2(new_n710), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n732), .A2(G97), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT46), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n706), .B2(new_n506), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n707), .A2(KEYINPUT46), .A3(G116), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT111), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(G107), .B2(new_n736), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n936), .A2(new_n937), .A3(new_n939), .A4(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n735), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n739), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n931), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT47), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n748), .ZN(new_n948));
  INV_X1    g0748(.A(new_n759), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n888), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n754), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n760), .B1(new_n221), .B2(new_n428), .C1(new_n239), .C2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n948), .A2(new_n762), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n923), .A2(KEYINPUT112), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT112), .B1(new_n923), .B2(new_n953), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n955), .ZN(G387));
  NAND2_X1  g0756(.A1(new_n905), .A2(new_n922), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n707), .A2(G77), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n372), .B2(new_n715), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n360), .B(new_n959), .C1(G159), .C2(new_n717), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n727), .A2(G150), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n721), .A2(new_n428), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n288), .B2(new_n709), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G50), .B2(new_n713), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n960), .A2(new_n937), .A3(new_n961), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n713), .A2(G317), .B1(new_n789), .B2(G311), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n745), .B2(new_n709), .C1(new_n944), .C2(new_n743), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT48), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n804), .B2(new_n721), .C1(new_n934), .C2(new_n706), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT49), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n727), .A2(G326), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n732), .A2(G116), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n971), .A2(new_n360), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n969), .A2(new_n970), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n965), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n951), .B1(new_n236), .B2(G45), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n660), .B2(new_n751), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n426), .A2(G50), .ZN(new_n979));
  XOR2_X1   g0779(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n288), .A2(new_n424), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n981), .A2(G45), .A3(new_n982), .A4(new_n660), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n978), .A2(new_n983), .B1(G107), .B2(new_n221), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n976), .A2(new_n748), .B1(new_n760), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n762), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n645), .A2(new_n949), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n657), .B(KEYINPUT114), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n906), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n905), .A2(new_n693), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n957), .B1(new_n986), .B2(new_n987), .C1(new_n989), .C2(new_n990), .ZN(G393));
  NAND4_X1  g0791(.A1(new_n648), .A2(new_n910), .A3(new_n914), .A4(new_n916), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n918), .A2(KEYINPUT115), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT115), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n917), .A2(new_n994), .A3(new_n647), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n919), .B(new_n988), .C1(new_n996), .C2(new_n907), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n891), .A2(new_n949), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G311), .A2(new_n713), .B1(new_n717), .B2(G317), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT52), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n399), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n804), .B2(new_n706), .C1(new_n743), .C2(new_n700), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n715), .A2(new_n745), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n709), .A2(new_n934), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n721), .A2(new_n506), .B1(new_n215), .B2(new_n723), .ZN(new_n1005));
  NOR4_X1   g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G150), .A2(new_n717), .B1(new_n713), .B2(G159), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT116), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT51), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n709), .A2(new_n426), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n360), .B1(new_n727), .B2(G143), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n288), .B2(new_n706), .C1(new_n424), .C2(new_n721), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n715), .A2(new_n205), .B1(new_n723), .B2(new_n476), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n748), .B1(new_n1006), .B2(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n760), .B1(new_n257), .B2(new_n221), .C1(new_n246), .C2(new_n951), .ZN(new_n1016));
  AND4_X1   g0816(.A1(new_n762), .A2(new_n998), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n996), .B2(new_n922), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n997), .A2(new_n1018), .ZN(G390));
  NAND2_X1  g0819(.A1(new_n857), .A2(G330), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1020), .A2(new_n626), .A3(new_n872), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n847), .A2(G330), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n685), .A2(G330), .A3(new_n779), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n868), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n867), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n691), .A2(new_n644), .A3(new_n779), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1029), .A2(new_n866), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n686), .A2(new_n779), .A3(new_n868), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n840), .A2(G330), .A3(new_n779), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1030), .B(new_n1031), .C1(new_n868), .C2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1022), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n869), .A2(new_n860), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n861), .A2(new_n1036), .A3(new_n863), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n836), .B(new_n860), .C1(new_n1030), .C2(new_n1025), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n1031), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1023), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1023), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1037), .A2(new_n1038), .A3(new_n1031), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1021), .B1(new_n1033), .B2(new_n1028), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1041), .A2(new_n1047), .A3(new_n988), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n861), .A2(new_n757), .A3(new_n863), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n372), .A2(new_n787), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n731), .A2(G294), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n789), .A2(G107), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n252), .B1(new_n714), .B2(new_n506), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n718), .A2(new_n804), .B1(new_n424), .B2(new_n721), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(G97), .C2(new_n710), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1051), .A2(new_n708), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n731), .A2(G125), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n789), .A2(G137), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT54), .B(G143), .Z(new_n1059));
  AOI22_X1  g0859(.A1(new_n710), .A2(new_n1059), .B1(new_n732), .B2(G50), .ZN(new_n1060));
  INV_X1    g0860(.A(G132), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n399), .B1(new_n701), .B2(new_n721), .C1(new_n714), .C2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G128), .B2(new_n717), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .A4(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n706), .A2(new_n389), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1066));
  XNOR2_X1  g0866(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n796), .A2(new_n1056), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n748), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1049), .A2(new_n762), .A3(new_n1050), .A4(new_n1069), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT118), .Z(new_n1071));
  NAND3_X1  g0871(.A1(new_n1044), .A2(new_n922), .A3(new_n1045), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1048), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(G378));
  NAND2_X1  g0874(.A1(new_n1047), .A2(new_n1022), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n864), .A2(new_n870), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n854), .A2(new_n855), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n848), .ZN(new_n1078));
  XOR2_X1   g0878(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1079));
  XOR2_X1   g0879(.A(new_n412), .B(new_n1079), .Z(new_n1080));
  AOI21_X1  g0880(.A(new_n633), .B1(new_n393), .B2(new_n396), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  AND4_X1   g0882(.A1(G330), .A2(new_n1077), .A3(new_n1078), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1082), .B1(new_n856), .B2(G330), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1076), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1077), .A2(G330), .A3(new_n1078), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1082), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n856), .A2(G330), .A3(new_n1082), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n871), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1075), .A2(KEYINPUT57), .A3(new_n1085), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT123), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1088), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n871), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1076), .A2(new_n1088), .A3(new_n1092), .A4(new_n1089), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1094), .A2(new_n1095), .B1(new_n1022), .B2(new_n1047), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n988), .B(new_n1091), .C1(new_n1096), .C2(KEYINPUT57), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1087), .A2(new_n758), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G68), .A2(new_n736), .B1(new_n717), .B2(G116), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT119), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n958), .C1(new_n257), .C2(new_n715), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(G41), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n732), .A2(G58), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n428), .B2(new_n709), .C1(new_n714), .C2(new_n215), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n731), .B2(G283), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(new_n1105), .A3(new_n360), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT120), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT58), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G150), .A2(new_n736), .B1(new_n717), .B2(G125), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(KEYINPUT121), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1110), .A2(new_n1111), .B1(G128), .B2(new_n713), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n789), .A2(G132), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n710), .A2(G137), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n707), .A2(new_n1059), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1117));
  OR2_X1    g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n732), .A2(G159), .ZN(new_n1119));
  AOI21_X1  g0919(.A(G41), .B1(new_n727), .B2(G124), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1118), .A2(new_n250), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1122));
  AOI21_X1  g0922(.A(G41), .B1(new_n333), .B2(G33), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1121), .A2(new_n1122), .B1(G50), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n748), .B1(new_n1108), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n787), .A2(new_n205), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n762), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1098), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n922), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1097), .A2(new_n1130), .ZN(G375));
  AND2_X1   g0931(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1021), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT124), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(KEYINPUT124), .A3(new_n1021), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n903), .B(new_n1046), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT125), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1103), .B1(new_n701), .B2(new_n706), .C1(new_n718), .C2(new_n1061), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n731), .B2(G128), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n713), .A2(G137), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n789), .A2(new_n1059), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n333), .B1(new_n721), .B2(new_n205), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G150), .B2(new_n710), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n730), .A2(new_n745), .B1(new_n257), .B2(new_n706), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT126), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n962), .B1(new_n215), .B2(new_n709), .C1(new_n718), .C2(new_n934), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n713), .A2(G283), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n789), .A2(G116), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1149), .A2(new_n252), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1145), .B1(new_n1152), .B2(new_n926), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n748), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n787), .A2(new_n288), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1025), .A2(new_n757), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1154), .A2(new_n762), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1132), .B2(new_n921), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1138), .A2(new_n1159), .ZN(G381));
  NOR3_X1   g0960(.A1(G387), .A2(G381), .A3(G384), .ZN(new_n1161));
  INV_X1    g0961(.A(G375), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1161), .A2(new_n1073), .A3(new_n1162), .A4(new_n1163), .ZN(G407));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1073), .ZN(new_n1165));
  OAI211_X1 g0965(.A(G407), .B(G213), .C1(G343), .C2(new_n1165), .ZN(G409));
  XOR2_X1   g0966(.A(G393), .B(G396), .Z(new_n1167));
  AOI21_X1  g0967(.A(G390), .B1(new_n923), .B2(new_n953), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n923), .A2(new_n953), .A3(G390), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(KEYINPUT127), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT127), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(G390), .C1(new_n923), .C2(new_n953), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1167), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1169), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(new_n1167), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n954), .A2(new_n955), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(G390), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1173), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1073), .B1(new_n1097), .B2(new_n1130), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n903), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1076), .B1(new_n1182), .B2(new_n1092), .ZN(new_n1183));
  AND4_X1   g0983(.A1(new_n1092), .A2(new_n1076), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1181), .B(new_n1075), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1128), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1085), .A2(new_n1090), .A3(new_n922), .ZN(new_n1187));
  AND4_X1   g0987(.A1(new_n1073), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1135), .A2(new_n1136), .B1(KEYINPUT60), .B2(new_n1035), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT60), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n988), .B1(new_n1133), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1159), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n785), .A3(new_n808), .ZN(new_n1193));
  OAI211_X1 g0993(.A(G384), .B(new_n1159), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(G213), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(G343), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1180), .A2(new_n1188), .A3(new_n1195), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT62), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1180), .A2(new_n1188), .A3(new_n1197), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(G2897), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1193), .A2(new_n1194), .A3(new_n1201), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1198), .A2(new_n1199), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1197), .B1(G375), .B2(G378), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1195), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1188), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1207), .A2(new_n1199), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT61), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1179), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT61), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1198), .A2(KEYINPUT63), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT63), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(G375), .A2(G378), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1197), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1209), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1204), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(new_n1202), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1216), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1214), .B(new_n1215), .C1(new_n1222), .C2(new_n1198), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1213), .A2(new_n1223), .ZN(G405));
  NAND2_X1  g1024(.A1(new_n1165), .A2(new_n1217), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1208), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1165), .A2(new_n1195), .A3(new_n1217), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1178), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1179), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(G402));
endmodule


