//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT28), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  AND2_X1   g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT0), .B(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT11), .A2(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT65), .A2(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT11), .A2(G134), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT11), .A2(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G137), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n208), .B2(new_n212), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n202), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n208), .A2(new_n212), .A3(new_n209), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n205), .A2(new_n217), .A3(new_n207), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n209), .B1(G134), .B2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n194), .B(new_n196), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT1), .B1(new_n195), .B2(G146), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n195), .A2(G146), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n193), .A2(G143), .ZN(new_n225));
  OAI211_X1 g039(.A(G128), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n216), .A2(new_n220), .A3(new_n222), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n215), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G116), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT2), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(G113), .ZN(new_n236));
  INV_X1    g050(.A(G113), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT2), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n232), .B(new_n234), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(new_n234), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n230), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n228), .A2(new_n229), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n192), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n228), .A2(new_n243), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n244), .B1(new_n215), .B2(new_n227), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n191), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT30), .B1(new_n228), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  AOI211_X1 g069(.A(KEYINPUT64), .B(new_n255), .C1(new_n215), .C2(new_n227), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n243), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n249), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n191), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT31), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n208), .A2(new_n212), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G131), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n201), .B1(new_n263), .B2(new_n216), .ZN(new_n264));
  AND4_X1   g078(.A1(new_n216), .A2(new_n222), .A3(new_n220), .A4(new_n226), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n253), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n255), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n228), .A2(new_n253), .A3(KEYINPUT30), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n249), .B1(new_n269), .B2(new_n243), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT31), .A3(new_n191), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n252), .B1(new_n261), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G472), .A2(G902), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT32), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n247), .A2(new_n251), .ZN(new_n276));
  INV_X1    g090(.A(new_n191), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT31), .B1(new_n270), .B2(new_n191), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n244), .B1(new_n267), .B2(new_n268), .ZN(new_n280));
  NOR4_X1   g094(.A1(new_n280), .A2(new_n260), .A3(new_n277), .A4(new_n249), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n273), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT68), .B(G902), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT28), .B1(new_n249), .B2(new_n250), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n247), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n277), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n276), .A2(new_n277), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n289), .B1(new_n270), .B2(new_n191), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n275), .A2(new_n284), .B1(new_n294), .B2(G472), .ZN(new_n295));
  INV_X1    g109(.A(G140), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G125), .ZN(new_n297));
  INV_X1    g111(.A(G125), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G140), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n297), .A2(new_n299), .A3(KEYINPUT70), .A4(KEYINPUT16), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n297), .A2(new_n299), .A3(KEYINPUT16), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n297), .B2(KEYINPUT16), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G146), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n193), .B(new_n300), .C1(new_n301), .C2(new_n303), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT24), .B(G110), .Z(new_n308));
  XNOR2_X1  g122(.A(G119), .B(G128), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G110), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n231), .A2(G128), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n312), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n221), .A2(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n231), .A2(G128), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n307), .B(new_n310), .C1(new_n311), .C2(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT71), .B(G110), .Z(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(KEYINPUT72), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n308), .A2(new_n309), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n324), .B1(new_n321), .B2(new_n317), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(KEYINPUT72), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT73), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n322), .A2(new_n325), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT72), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n328), .A4(new_n326), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G125), .B(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n193), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n305), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT74), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n344));
  AOI211_X1 g158(.A(new_n344), .B(new_n341), .C1(new_n332), .C2(new_n337), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n323), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G953), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G221), .A3(G234), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT75), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n323), .B(new_n351), .C1(new_n343), .C2(new_n345), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G217), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n285), .B2(G234), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n355), .A2(G902), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n357), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n285), .A3(new_n354), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n353), .A2(KEYINPUT25), .A3(new_n285), .A4(new_n354), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n295), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT9), .B(G234), .ZN(new_n366));
  OAI21_X1  g180(.A(G221), .B1(new_n366), .B2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT78), .B(G469), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n213), .A2(new_n214), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(G104), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(G104), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT76), .A3(G107), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G101), .ZN(new_n379));
  INV_X1    g193(.A(G101), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(G107), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n373), .A2(KEYINPUT3), .A3(G104), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n373), .B2(G104), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n379), .A2(new_n384), .A3(new_n222), .A4(new_n226), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n379), .A2(new_n384), .B1(new_n226), .B2(new_n222), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n371), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT12), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n389), .A2(KEYINPUT77), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(KEYINPUT77), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n379), .A2(new_n384), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n226), .A2(new_n222), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n370), .B1(new_n395), .B2(new_n385), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT77), .A3(new_n389), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n385), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n226), .A2(new_n222), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n400), .A2(KEYINPUT10), .A3(new_n384), .A4(new_n379), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G101), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n373), .A2(G104), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n376), .B2(G107), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n373), .A2(KEYINPUT3), .A3(G104), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT4), .B1(new_n409), .B2(new_n380), .ZN(new_n410));
  AOI211_X1 g224(.A(G101), .B(new_n405), .C1(new_n407), .C2(new_n408), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n404), .B(new_n202), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n399), .A2(new_n401), .A3(new_n412), .A4(new_n370), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n347), .A2(G227), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n392), .A2(new_n397), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n399), .A2(new_n401), .A3(new_n412), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n371), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n420), .B2(new_n413), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n418), .B1(new_n421), .B2(KEYINPUT79), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n423), .B(new_n417), .C1(new_n420), .C2(new_n413), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n285), .B(new_n369), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n392), .A2(new_n413), .A3(new_n397), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n413), .A2(new_n417), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n426), .A2(new_n416), .B1(new_n427), .B2(new_n420), .ZN(new_n428));
  OAI21_X1  g242(.A(G469), .B1(new_n428), .B2(G902), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n368), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n433));
  AOI21_X1  g247(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n434));
  OAI21_X1  g248(.A(G131), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT17), .ZN(new_n436));
  INV_X1    g250(.A(G237), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n347), .A3(G214), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n195), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n209), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n435), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT17), .B(G131), .C1(new_n433), .C2(new_n434), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n305), .A2(new_n442), .A3(new_n306), .A4(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G113), .B(G122), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(new_n376), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n439), .A2(new_n447), .A3(new_n440), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT18), .A2(G131), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n297), .A2(new_n299), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G146), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n448), .A2(new_n450), .B1(new_n452), .B2(new_n340), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n450), .B2(new_n448), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n444), .A2(new_n446), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n435), .A2(new_n441), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n451), .B1(new_n457), .B2(KEYINPUT19), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n458), .B1(new_n451), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n305), .B(new_n456), .C1(G146), .C2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n446), .B1(new_n461), .B2(new_n454), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n464));
  NOR2_X1   g278(.A1(G475), .A2(G902), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n465), .B1(new_n455), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT20), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G475), .ZN(new_n470));
  INV_X1    g284(.A(G902), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n446), .B1(new_n444), .B2(new_n454), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n455), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n473), .B2(KEYINPUT86), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(new_n471), .C1(new_n455), .C2(new_n472), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n366), .A2(new_n356), .A3(G953), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n233), .A2(G122), .ZN(new_n482));
  INV_X1    g296(.A(G122), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G116), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n484), .A3(new_n373), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n195), .A2(G128), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n221), .A2(G143), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n217), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n217), .B1(new_n486), .B2(new_n487), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT87), .B1(new_n482), .B2(KEYINPUT14), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT87), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT14), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n233), .A4(G122), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n482), .A2(KEYINPUT14), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n484), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n491), .B1(G107), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n482), .A2(new_n484), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G107), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n485), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT13), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n221), .B2(G143), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n487), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n486), .A2(new_n502), .ZN(new_n505));
  OAI21_X1  g319(.A(G134), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n501), .A2(new_n506), .A3(new_n488), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n481), .B1(new_n498), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n497), .A2(G107), .ZN(new_n509));
  INV_X1    g323(.A(new_n485), .ZN(new_n510));
  INV_X1    g324(.A(new_n490), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n488), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n489), .B1(new_n500), .B2(new_n485), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n506), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT88), .A4(new_n480), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n512), .A2(new_n509), .B1(new_n514), .B2(new_n506), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT88), .B1(new_n518), .B2(new_n480), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n285), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT89), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G478), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT89), .B(new_n285), .C1(new_n517), .C2(new_n519), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n520), .A2(new_n524), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI211_X1 g342(.A(new_n347), .B(new_n285), .C1(G234), .C2(G237), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT21), .B(G898), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G952), .ZN(new_n532));
  AOI211_X1 g346(.A(G953), .B(new_n532), .C1(G234), .C2(G237), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n479), .A2(new_n528), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G214), .B1(G237), .B2(G902), .ZN(new_n537));
  OAI21_X1  g351(.A(G210), .B1(G237), .B2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n404), .B(new_n243), .C1(new_n410), .C2(new_n411), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n232), .A2(new_n234), .A3(KEYINPUT5), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n541), .B(G113), .C1(KEYINPUT5), .C2(new_n232), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n542), .A2(new_n379), .A3(new_n239), .A4(new_n384), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(G110), .B(G122), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n540), .A2(new_n543), .A3(new_n545), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(KEYINPUT6), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT6), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(new_n550), .A3(new_n546), .ZN(new_n551));
  AOI21_X1  g365(.A(G125), .B1(new_n226), .B2(new_n222), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(G125), .B2(new_n201), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n347), .A2(G224), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n549), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n545), .B(KEYINPUT8), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n542), .A2(new_n239), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n393), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT81), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT81), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n393), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n558), .B1(new_n564), .B2(new_n543), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n554), .A2(KEYINPUT7), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT82), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n552), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n201), .A2(G125), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n552), .B2(new_n567), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n553), .A2(KEYINPUT7), .A3(new_n554), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n548), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n471), .B1(new_n565), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n539), .B1(new_n556), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n571), .A2(new_n572), .A3(new_n548), .ZN(new_n576));
  INV_X1    g390(.A(new_n563), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n562), .B1(new_n559), .B2(new_n393), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n543), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n557), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n549), .A2(new_n551), .A3(new_n555), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n538), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n575), .A2(KEYINPUT83), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT83), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(new_n539), .C1(new_n556), .C2(new_n574), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n536), .A2(new_n537), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n365), .A2(new_n432), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  NAND2_X1  g404(.A1(new_n282), .A2(new_n285), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n282), .A2(new_n273), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n362), .A2(new_n363), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n358), .B1(new_n596), .B2(new_n357), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n595), .A2(new_n432), .A3(new_n597), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n517), .A2(new_n519), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n518), .A2(new_n480), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n508), .A2(KEYINPUT33), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n599), .A2(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(G478), .A3(new_n285), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n537), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n575), .B2(new_n583), .ZN(new_n608));
  AND4_X1   g422(.A1(new_n478), .A2(new_n606), .A3(new_n535), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n598), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  NAND2_X1  g426(.A1(new_n526), .A2(new_n527), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n466), .A2(new_n468), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT90), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n477), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n474), .A2(KEYINPUT90), .A3(new_n476), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n613), .A2(new_n618), .A3(new_n535), .A4(new_n608), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n598), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n620), .B(KEYINPUT91), .Z(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT35), .B(G107), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  NAND2_X1  g437(.A1(new_n596), .A2(new_n357), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n346), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n357), .A2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n346), .A2(new_n625), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n588), .A2(new_n432), .A3(new_n595), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT37), .B(G110), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G12));
  NAND2_X1  g448(.A1(new_n294), .A2(G472), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n272), .A2(KEYINPUT32), .A3(new_n274), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n283), .B1(new_n282), .B2(new_n273), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n432), .A2(new_n638), .A3(new_n608), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT92), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n529), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n534), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n474), .A2(KEYINPUT90), .A3(new_n476), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT90), .B1(new_n474), .B2(new_n476), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n469), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n640), .B1(new_n646), .B2(new_n528), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n618), .A2(KEYINPUT92), .A3(new_n613), .A4(new_n643), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n647), .B(new_n648), .C1(new_n364), .C2(new_n629), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n639), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n221), .ZN(G30));
  NAND2_X1  g465(.A1(new_n275), .A2(new_n284), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n191), .B1(new_n280), .B2(new_n249), .ZN(new_n653));
  OR3_X1    g467(.A1(new_n249), .A2(new_n191), .A3(new_n250), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(KEYINPUT94), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n471), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT94), .B1(new_n653), .B2(new_n654), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT95), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(KEYINPUT95), .B(G472), .C1(new_n656), .C2(new_n657), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n652), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT96), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n587), .B(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n478), .A2(new_n613), .A3(new_n537), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n665), .A2(new_n631), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT97), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n663), .A2(KEYINPUT97), .A3(new_n667), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n643), .B(KEYINPUT39), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n432), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT40), .Z(new_n674));
  NAND3_X1  g488(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  INV_X1    g490(.A(new_n608), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n652), .B2(new_n635), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n606), .A2(new_n478), .A3(new_n643), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n631), .A3(new_n432), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  OAI21_X1  g495(.A(new_n285), .B1(new_n422), .B2(new_n424), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n367), .A3(new_n425), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n365), .A2(KEYINPUT98), .A3(new_n609), .A4(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n638), .A2(new_n597), .A3(new_n609), .A4(new_n685), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT98), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  NAND4_X1  g506(.A1(new_n619), .A2(new_n638), .A3(new_n597), .A4(new_n685), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  NAND3_X1  g508(.A1(new_n631), .A2(new_n638), .A3(new_n536), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n608), .A2(new_n683), .A3(new_n367), .A4(new_n425), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n696), .A2(KEYINPUT99), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(KEYINPUT99), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n231), .ZN(G21));
  NAND4_X1  g515(.A1(new_n608), .A2(new_n478), .A3(new_n613), .A4(new_n535), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n684), .ZN(new_n703));
  OAI22_X1  g517(.A1(new_n279), .A2(new_n281), .B1(new_n191), .B2(new_n288), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n273), .B(KEYINPUT100), .Z(new_n705));
  AOI22_X1  g519(.A1(new_n591), .A2(G472), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n597), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT101), .B(G122), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G24));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n629), .B1(new_n596), .B2(new_n357), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n704), .A2(new_n705), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n592), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n710), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n706), .B(KEYINPUT102), .C1(new_n364), .C2(new_n629), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n679), .ZN(new_n717));
  INV_X1    g531(.A(new_n698), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n696), .A2(KEYINPUT99), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n367), .A2(new_n537), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n584), .B2(new_n586), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n425), .A2(new_n429), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n425), .A2(KEYINPUT103), .A3(new_n429), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n725), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n638), .A3(new_n597), .A4(new_n679), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n723), .B1(new_n731), .B2(KEYINPUT104), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(KEYINPUT105), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n731), .B1(KEYINPUT104), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n209), .ZN(G33));
  NAND4_X1  g552(.A1(new_n365), .A2(new_n647), .A3(new_n648), .A4(new_n730), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  INV_X1    g555(.A(G469), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n426), .A2(new_n416), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n427), .A2(new_n420), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n742), .A2(new_n471), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n741), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n751), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n747), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n753), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n754), .A2(new_n759), .A3(new_n425), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n760), .A2(new_n367), .A3(new_n672), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n479), .A2(new_n606), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n594), .A3(new_n631), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n607), .B1(new_n584), .B2(new_n586), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n631), .A3(KEYINPUT44), .A4(new_n594), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n761), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT107), .B(G137), .Z(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G39));
  NAND2_X1  g586(.A1(new_n760), .A2(new_n367), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n768), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n638), .A2(new_n597), .A3(new_n717), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n687), .B(KEYINPUT98), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n693), .B(new_n707), .C1(new_n695), .C2(new_n699), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n782), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT110), .A3(new_n690), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n730), .A2(new_n679), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n613), .A2(KEYINPUT111), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n613), .A2(KEYINPUT111), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n646), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n432), .A2(new_n768), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n711), .A2(new_n295), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n716), .A2(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n734), .A2(new_n793), .A3(new_n736), .A4(new_n739), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n479), .B1(new_n788), .B2(new_n789), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n606), .A2(new_n478), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n587), .A2(new_n537), .A3(new_n535), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n598), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n589), .A3(new_n632), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n786), .A2(new_n794), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n679), .B1(new_n697), .B2(new_n698), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n714), .B2(new_n715), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n643), .A2(new_n367), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n677), .A2(new_n479), .A3(new_n528), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n728), .A2(new_n729), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n662), .A2(new_n711), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n680), .A2(new_n809), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n805), .A2(new_n810), .A3(new_n650), .A4(KEYINPUT52), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n430), .B(KEYINPUT80), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n295), .A3(new_n677), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n647), .A2(new_n648), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n711), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n716), .A2(new_n720), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT112), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n805), .B2(new_n650), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n817), .A2(new_n819), .A3(new_n680), .A4(new_n809), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n811), .B1(new_n820), .B2(KEYINPUT52), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n803), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n801), .B1(new_n783), .B2(new_n785), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  INV_X1    g638(.A(new_n810), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n824), .B1(new_n816), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n811), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n827), .A3(new_n794), .ZN(new_n828));
  XOR2_X1   g642(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n802), .A2(new_n784), .A3(KEYINPUT53), .A4(new_n690), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n734), .A2(new_n793), .A3(new_n736), .A4(new_n739), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n821), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n832), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n764), .A2(new_n533), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n713), .A2(new_n358), .A3(new_n364), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n683), .A2(new_n425), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n367), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n768), .B(new_n843), .C1(new_n775), .C2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT50), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n537), .B(new_n684), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n850), .A2(new_n665), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n843), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n843), .B(new_n851), .C1(new_n848), .C2(new_n849), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n776), .A2(new_n684), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n840), .A2(new_n716), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n663), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n855), .A2(new_n597), .A3(new_n533), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n606), .A2(new_n478), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n853), .A2(new_n854), .A3(new_n856), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n847), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n847), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n842), .A2(new_n699), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n532), .A3(G953), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n857), .A2(new_n478), .A3(new_n606), .A4(new_n858), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n866), .A2(KEYINPUT116), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT116), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n840), .A2(new_n365), .A3(new_n855), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT48), .Z(new_n871));
  NOR3_X1   g685(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n863), .A2(new_n864), .A3(new_n872), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n839), .A2(new_n873), .B1(G952), .B2(G953), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n762), .A2(new_n724), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n597), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n876), .A2(KEYINPUT108), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n844), .B(KEYINPUT49), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n665), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n876), .A2(KEYINPUT108), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n663), .A2(new_n877), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT109), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n874), .A2(new_n882), .ZN(G75));
  NOR2_X1   g697(.A1(new_n347), .A2(G952), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n285), .B1(new_n832), .B2(new_n836), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(new_n539), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n549), .A2(new_n551), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n555), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n885), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n886), .A2(new_n539), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n893), .A2(new_n896), .ZN(G51));
  XNOR2_X1  g711(.A(new_n753), .B(KEYINPUT118), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT57), .Z(new_n899));
  AND3_X1   g713(.A1(new_n832), .A2(new_n836), .A3(new_n837), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n837), .B1(new_n832), .B2(new_n836), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n422), .A2(new_n424), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n886), .A2(new_n752), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n884), .B1(new_n904), .B2(new_n905), .ZN(G54));
  NAND2_X1  g720(.A1(new_n832), .A2(new_n836), .ZN(new_n907));
  AND2_X1   g721(.A1(KEYINPUT58), .A2(G475), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n463), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n286), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n885), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n463), .B1(new_n886), .B2(new_n908), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT119), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n907), .A2(new_n286), .A3(new_n908), .ZN(new_n914));
  INV_X1    g728(.A(new_n463), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n884), .B1(new_n886), .B2(new_n909), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n913), .A2(new_n919), .ZN(G60));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT59), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n603), .B1(new_n839), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n603), .A2(new_n922), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n900), .B2(new_n901), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n885), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n923), .A2(new_n926), .ZN(G63));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n928));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n832), .B2(new_n836), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n626), .A2(new_n628), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n355), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n885), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n928), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n832), .A2(new_n836), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n355), .B1(new_n938), .B2(new_n930), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(KEYINPUT61), .A3(new_n885), .A4(new_n933), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(G66));
  INV_X1    g755(.A(G224), .ZN(new_n942));
  OAI21_X1  g756(.A(G953), .B1(new_n530), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n823), .B(KEYINPUT120), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n944), .A2(KEYINPUT121), .A3(new_n347), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT121), .B1(new_n944), .B2(new_n347), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n888), .B1(G898), .B2(new_n347), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n948), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n950), .B(new_n943), .C1(new_n945), .C2(new_n946), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(G69));
  AOI21_X1  g766(.A(new_n347), .B1(G227), .B2(G900), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n770), .A2(new_n817), .A3(new_n819), .A4(new_n680), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n955));
  INV_X1    g769(.A(new_n680), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n721), .B1(new_n639), .B2(new_n649), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n818), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n959), .A3(new_n770), .A4(new_n817), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n734), .A2(new_n736), .A3(new_n739), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n734), .A2(new_n964), .A3(new_n736), .A4(new_n739), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n677), .A2(new_n479), .A3(new_n528), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n761), .A2(new_n365), .A3(new_n966), .ZN(new_n967));
  AND4_X1   g781(.A1(new_n778), .A2(new_n963), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n961), .A2(new_n968), .A3(new_n347), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n269), .B(KEYINPUT122), .Z(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(new_n460), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(G900), .B2(G953), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n953), .B1(new_n973), .B2(KEYINPUT123), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n797), .A2(new_n776), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n975), .A2(new_n365), .A3(new_n432), .A4(new_n672), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n778), .A2(new_n770), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n817), .A2(new_n819), .A3(new_n680), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n958), .A2(new_n675), .A3(KEYINPUT62), .A4(new_n817), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n971), .B1(new_n983), .B2(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n973), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n974), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n984), .B(new_n973), .C1(KEYINPUT123), .C2(new_n953), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(G72));
  XNOR2_X1  g802(.A(new_n270), .B(new_n277), .ZN(new_n989));
  XNOR2_X1  g803(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n990));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n885), .ZN(new_n994));
  INV_X1    g808(.A(new_n653), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n983), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n961), .A2(new_n968), .A3(new_n277), .A4(new_n270), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n944), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n822), .A2(new_n830), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n989), .A2(new_n992), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n994), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(G57));
endmodule


