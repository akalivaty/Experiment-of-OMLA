

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590;

  XNOR2_X1 U321 ( .A(n321), .B(n320), .ZN(n325) );
  XNOR2_X1 U322 ( .A(n316), .B(n315), .ZN(n432) );
  XNOR2_X1 U323 ( .A(n453), .B(n452), .ZN(n527) );
  XNOR2_X1 U324 ( .A(n327), .B(n326), .ZN(n517) );
  NOR2_X1 U325 ( .A1(n488), .A2(n500), .ZN(n482) );
  OR2_X1 U326 ( .A1(n570), .A2(n467), .ZN(n289) );
  AND2_X1 U327 ( .A1(n464), .A2(n289), .ZN(n290) );
  INV_X1 U328 ( .A(KEYINPUT85), .ZN(n313) );
  XNOR2_X1 U329 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U330 ( .A(n369), .B(KEYINPUT76), .ZN(n370) );
  INV_X1 U331 ( .A(KEYINPUT92), .ZN(n318) );
  XNOR2_X1 U332 ( .A(n371), .B(n370), .ZN(n374) );
  XNOR2_X1 U333 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U334 ( .A(n376), .B(G155GAT), .ZN(n377) );
  NOR2_X1 U335 ( .A1(n486), .A2(n485), .ZN(n487) );
  NOR2_X1 U336 ( .A1(n419), .A2(n514), .ZN(n572) );
  XNOR2_X1 U337 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U338 ( .A(KEYINPUT110), .B(n583), .ZN(n568) );
  XNOR2_X1 U339 ( .A(KEYINPUT38), .B(n489), .ZN(n498) );
  XNOR2_X1 U340 ( .A(n456), .B(G190GAT), .ZN(n457) );
  XNOR2_X1 U341 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(G43GAT), .B(G50GAT), .Z(n292) );
  XNOR2_X1 U343 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n291) );
  XNOR2_X1 U344 ( .A(n292), .B(n291), .ZN(n328) );
  XOR2_X1 U345 ( .A(G36GAT), .B(G190GAT), .Z(n317) );
  XNOR2_X1 U346 ( .A(n328), .B(n317), .ZN(n293) );
  XOR2_X1 U347 ( .A(G29GAT), .B(G134GAT), .Z(n410) );
  XNOR2_X1 U348 ( .A(n293), .B(n410), .ZN(n299) );
  XOR2_X1 U349 ( .A(G85GAT), .B(KEYINPUT68), .Z(n295) );
  XNOR2_X1 U350 ( .A(G99GAT), .B(G106GAT), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n349) );
  XOR2_X1 U352 ( .A(n349), .B(G92GAT), .Z(n297) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U355 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U356 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n301) );
  XNOR2_X1 U357 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U359 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n303) );
  XNOR2_X1 U360 ( .A(G162GAT), .B(KEYINPUT9), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n558) );
  INV_X1 U364 ( .A(n558), .ZN(n455) );
  XNOR2_X1 U365 ( .A(G8GAT), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n308), .B(KEYINPUT74), .ZN(n372) );
  XOR2_X1 U367 ( .A(G64GAT), .B(G92GAT), .Z(n310) );
  XNOR2_X1 U368 ( .A(G176GAT), .B(G204GAT), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n358) );
  XNOR2_X1 U370 ( .A(n372), .B(n358), .ZN(n327) );
  XOR2_X1 U371 ( .A(KEYINPUT21), .B(KEYINPUT84), .Z(n312) );
  XNOR2_X1 U372 ( .A(G218GAT), .B(KEYINPUT83), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n316) );
  XNOR2_X1 U374 ( .A(G197GAT), .B(G211GAT), .ZN(n314) );
  XOR2_X1 U375 ( .A(n317), .B(n432), .Z(n321) );
  NAND2_X1 U376 ( .A1(G226GAT), .A2(G233GAT), .ZN(n319) );
  XOR2_X1 U377 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n323) );
  XNOR2_X1 U378 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n445) );
  XNOR2_X1 U380 ( .A(n445), .B(KEYINPUT91), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U382 ( .A(KEYINPUT120), .B(n517), .ZN(n394) );
  XNOR2_X1 U383 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n393) );
  XOR2_X1 U384 ( .A(G22GAT), .B(G15GAT), .Z(n375) );
  XOR2_X1 U385 ( .A(n328), .B(n375), .Z(n330) );
  NAND2_X1 U386 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U388 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n332) );
  XNOR2_X1 U389 ( .A(KEYINPUT67), .B(KEYINPUT66), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U391 ( .A(n334), .B(n333), .Z(n342) );
  XOR2_X1 U392 ( .A(G141GAT), .B(G197GAT), .Z(n336) );
  XNOR2_X1 U393 ( .A(G36GAT), .B(G29GAT), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U395 ( .A(G1GAT), .B(G8GAT), .Z(n338) );
  XNOR2_X1 U396 ( .A(G169GAT), .B(G113GAT), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n573) );
  INV_X1 U400 ( .A(n573), .ZN(n546) );
  XOR2_X1 U401 ( .A(G120GAT), .B(G148GAT), .Z(n405) );
  XOR2_X1 U402 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n344) );
  XNOR2_X1 U403 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U405 ( .A(n405), .B(n345), .Z(n347) );
  NAND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U408 ( .A(n348), .B(KEYINPUT33), .Z(n351) );
  XNOR2_X1 U409 ( .A(n349), .B(KEYINPUT32), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n360) );
  INV_X1 U411 ( .A(KEYINPUT13), .ZN(n352) );
  NAND2_X1 U412 ( .A1(n352), .A2(G57GAT), .ZN(n355) );
  INV_X1 U413 ( .A(G57GAT), .ZN(n353) );
  NAND2_X1 U414 ( .A1(n353), .A2(KEYINPUT13), .ZN(n354) );
  NAND2_X1 U415 ( .A1(n355), .A2(n354), .ZN(n357) );
  XNOR2_X1 U416 ( .A(G71GAT), .B(G78GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n365) );
  XOR2_X1 U418 ( .A(n365), .B(n358), .Z(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n388) );
  INV_X1 U420 ( .A(n388), .ZN(n579) );
  XNOR2_X1 U421 ( .A(n579), .B(KEYINPUT41), .ZN(n550) );
  NAND2_X1 U422 ( .A1(n546), .A2(n550), .ZN(n361) );
  XNOR2_X1 U423 ( .A(KEYINPUT46), .B(n361), .ZN(n381) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(G64GAT), .Z(n363) );
  XNOR2_X1 U425 ( .A(KEYINPUT14), .B(KEYINPUT75), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n380) );
  INV_X1 U427 ( .A(n365), .ZN(n364) );
  XOR2_X1 U428 ( .A(G1GAT), .B(G127GAT), .Z(n406) );
  NAND2_X1 U429 ( .A1(n364), .A2(n406), .ZN(n368) );
  INV_X1 U430 ( .A(n406), .ZN(n366) );
  NAND2_X1 U431 ( .A1(n366), .A2(n365), .ZN(n367) );
  NAND2_X1 U432 ( .A1(n368), .A2(n367), .ZN(n371) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XOR2_X1 U434 ( .A(n372), .B(KEYINPUT15), .Z(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U436 ( .A(n375), .B(G211GAT), .Z(n376) );
  XOR2_X1 U437 ( .A(n380), .B(n379), .Z(n555) );
  INV_X1 U438 ( .A(n555), .ZN(n583) );
  NAND2_X1 U439 ( .A1(n381), .A2(n568), .ZN(n382) );
  NOR2_X1 U440 ( .A1(n382), .A2(n558), .ZN(n383) );
  XNOR2_X1 U441 ( .A(KEYINPUT47), .B(n383), .ZN(n391) );
  XOR2_X1 U442 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n385) );
  XNOR2_X1 U443 ( .A(KEYINPUT36), .B(n558), .ZN(n586) );
  NAND2_X1 U444 ( .A1(n555), .A2(n586), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  NAND2_X1 U446 ( .A1(n573), .A2(n386), .ZN(n387) );
  NOR2_X1 U447 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U448 ( .A(KEYINPUT111), .B(n389), .ZN(n390) );
  NAND2_X1 U449 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X2 U450 ( .A(n393), .B(n392), .ZN(n543) );
  NAND2_X1 U451 ( .A1(n394), .A2(n543), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n395), .B(KEYINPUT54), .ZN(n396) );
  XOR2_X1 U453 ( .A(KEYINPUT121), .B(n396), .Z(n419) );
  XOR2_X1 U454 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n398) );
  XNOR2_X1 U455 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U457 ( .A(n399), .B(KEYINPUT3), .Z(n401) );
  XNOR2_X1 U458 ( .A(G141GAT), .B(G155GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n431) );
  XOR2_X1 U460 ( .A(KEYINPUT1), .B(KEYINPUT88), .Z(n403) );
  XNOR2_X1 U461 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n431), .B(n404), .ZN(n418) );
  XOR2_X1 U464 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n408) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n414) );
  XNOR2_X1 U467 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n409), .B(KEYINPUT77), .ZN(n443) );
  XOR2_X1 U469 ( .A(n410), .B(n443), .Z(n412) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U472 ( .A(n414), .B(n413), .Z(n416) );
  XNOR2_X1 U473 ( .A(G85GAT), .B(G57GAT), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n465) );
  XNOR2_X1 U476 ( .A(KEYINPUT90), .B(n465), .ZN(n514) );
  XOR2_X1 U477 ( .A(KEYINPUT81), .B(G78GAT), .Z(n421) );
  XNOR2_X1 U478 ( .A(G50GAT), .B(G106GAT), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U480 ( .A(KEYINPUT23), .B(G148GAT), .Z(n423) );
  XNOR2_X1 U481 ( .A(G22GAT), .B(G204GAT), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U483 ( .A(n425), .B(n424), .Z(n430) );
  XOR2_X1 U484 ( .A(KEYINPUT82), .B(KEYINPUT22), .Z(n427) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U487 ( .A(KEYINPUT24), .B(n428), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U489 ( .A(n432), .B(n431), .Z(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n469) );
  NAND2_X1 U491 ( .A1(n572), .A2(n469), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n435), .B(KEYINPUT55), .ZN(n454) );
  XOR2_X1 U493 ( .A(G176GAT), .B(KEYINPUT78), .Z(n437) );
  XNOR2_X1 U494 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n453) );
  XOR2_X1 U496 ( .A(G120GAT), .B(G127GAT), .Z(n439) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(G134GAT), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U499 ( .A(G190GAT), .B(G99GAT), .Z(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n449) );
  XNOR2_X1 U501 ( .A(G183GAT), .B(KEYINPUT20), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n442), .B(G71GAT), .ZN(n444) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n447) );
  XNOR2_X1 U504 ( .A(G15GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n451) );
  NAND2_X1 U507 ( .A1(G227GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n452) );
  NAND2_X1 U509 ( .A1(n454), .A2(n527), .ZN(n567) );
  NOR2_X1 U510 ( .A1(n455), .A2(n567), .ZN(n458) );
  INV_X1 U511 ( .A(KEYINPUT58), .ZN(n456) );
  NAND2_X1 U512 ( .A1(n579), .A2(n546), .ZN(n488) );
  NOR2_X1 U513 ( .A1(n558), .A2(n583), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n459), .B(KEYINPUT16), .ZN(n473) );
  NAND2_X1 U515 ( .A1(n527), .A2(n517), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n460), .A2(n469), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n461), .B(KEYINPUT25), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT93), .ZN(n464) );
  NOR2_X1 U519 ( .A1(n469), .A2(n527), .ZN(n463) );
  XOR2_X1 U520 ( .A(n463), .B(KEYINPUT26), .Z(n570) );
  XOR2_X1 U521 ( .A(n517), .B(KEYINPUT27), .Z(n467) );
  NOR2_X1 U522 ( .A1(n465), .A2(n290), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT94), .ZN(n471) );
  INV_X1 U524 ( .A(n514), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n544) );
  XNOR2_X1 U526 ( .A(KEYINPUT28), .B(n469), .ZN(n481) );
  NAND2_X1 U527 ( .A1(n544), .A2(n481), .ZN(n529) );
  NOR2_X1 U528 ( .A1(n527), .A2(n529), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n471), .A2(n470), .ZN(n486) );
  INV_X1 U530 ( .A(n486), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n500) );
  NAND2_X1 U532 ( .A1(n514), .A2(n482), .ZN(n477) );
  XOR2_X1 U533 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n475) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n482), .A2(n517), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U540 ( .A1(n482), .A2(n527), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  XOR2_X1 U542 ( .A(G22GAT), .B(KEYINPUT97), .Z(n484) );
  INV_X1 U543 ( .A(n481), .ZN(n521) );
  NAND2_X1 U544 ( .A1(n482), .A2(n521), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT39), .Z(n491) );
  NAND2_X1 U547 ( .A1(n586), .A2(n583), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT37), .ZN(n513) );
  NOR2_X1 U549 ( .A1(n513), .A2(n488), .ZN(n489) );
  NAND2_X1 U550 ( .A1(n498), .A2(n514), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n498), .A2(n517), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(KEYINPUT98), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n497) );
  XOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n495) );
  NAND2_X1 U557 ( .A1(n498), .A2(n527), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n521), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT101), .B(n550), .ZN(n562) );
  INV_X1 U564 ( .A(n562), .ZN(n532) );
  NAND2_X1 U565 ( .A1(n573), .A2(n532), .ZN(n512) );
  NOR2_X1 U566 ( .A1(n512), .A2(n500), .ZN(n508) );
  NAND2_X1 U567 ( .A1(n508), .A2(n514), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n503), .Z(G1332GAT) );
  XOR2_X1 U570 ( .A(G64GAT), .B(KEYINPUT103), .Z(n505) );
  NAND2_X1 U571 ( .A1(n508), .A2(n517), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n505), .B(n504), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n527), .A2(n508), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n506), .B(KEYINPUT104), .ZN(n507) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U577 ( .A1(n508), .A2(n521), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n511), .Z(G1335GAT) );
  NOR2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n514), .A2(n522), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(KEYINPUT106), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n522), .A2(n517), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U586 ( .A(G99GAT), .B(KEYINPUT107), .Z(n520) );
  NAND2_X1 U587 ( .A1(n522), .A2(n527), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n526) );
  XOR2_X1 U590 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n524) );
  NAND2_X1 U591 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT113), .Z(n531) );
  NAND2_X1 U595 ( .A1(n527), .A2(n543), .ZN(n528) );
  NOR2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n540), .A2(n546), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n534) );
  NAND2_X1 U600 ( .A1(n540), .A2(n532), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(n535), .ZN(G1341GAT) );
  INV_X1 U603 ( .A(n540), .ZN(n536) );
  NOR2_X1 U604 ( .A1(n568), .A2(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U609 ( .A1(n540), .A2(n558), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n548) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U613 ( .A1(n570), .A2(n545), .ZN(n559) );
  NAND2_X1 U614 ( .A1(n559), .A2(n546), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n554) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U619 ( .A1(n559), .A2(n550), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  XOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT119), .Z(n557) );
  NAND2_X1 U623 ( .A1(n559), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U627 ( .A1(n573), .A2(n567), .ZN(n561) );
  XOR2_X1 U628 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n567), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  INV_X1 U636 ( .A(n570), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n585) );
  NOR2_X1 U638 ( .A1(n573), .A2(n585), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(KEYINPUT123), .B(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n585), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n589) );
  INV_X1 U651 ( .A(n585), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(G218GAT), .B(n590), .Z(G1355GAT) );
endmodule

