//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n453), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  AND2_X1   g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(new_n463), .B2(new_n464), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  MUX2_X1   g053(.A(G100), .B(G112), .S(G2105), .Z(new_n479));
  AOI22_X1  g054(.A1(G136), .A2(new_n465), .B1(new_n479), .B2(G2104), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n478), .A2(new_n480), .ZN(G162));
  AND2_X1   g056(.A1(KEYINPUT70), .A2(G114), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT70), .A2(G114), .ZN(new_n483));
  OAI21_X1  g058(.A(G2105), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n475), .A2(G102), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n486), .A2(G2104), .B1(G126), .B2(new_n476), .ZN(new_n487));
  AND2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n475), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n463), .A2(new_n464), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n492), .A2(new_n493), .A3(G138), .A4(new_n475), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n487), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  OR2_X1    g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT71), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT71), .A2(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT6), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n500), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G88), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n508), .B1(new_n505), .B2(new_n502), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n500), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n503), .A2(new_n504), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n507), .A2(new_n510), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND2_X1  g093(.A1(new_n509), .A2(G51), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n498), .A2(new_n499), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT71), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT71), .A2(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g099(.A(G89), .B(new_n520), .C1(new_n524), .C2(new_n501), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n520), .B2(new_n529), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n519), .A2(new_n525), .A3(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n509), .A2(G52), .ZN(new_n532));
  OAI211_X1 g107(.A(G90), .B(new_n520), .C1(new_n524), .C2(new_n501), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n498), .B2(new_n499), .ZN(new_n535));
  AND2_X1   g110(.A1(G77), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n515), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(new_n506), .A2(G81), .ZN(new_n540));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n500), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(new_n515), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n509), .A2(G43), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  OAI21_X1  g127(.A(new_n520), .B1(new_n524), .B2(new_n501), .ZN(new_n553));
  INV_X1    g128(.A(G91), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G651), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n553), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(KEYINPUT72), .B2(KEYINPUT9), .ZN(new_n560));
  OAI211_X1 g135(.A(G543), .B(new_n560), .C1(new_n524), .C2(new_n501), .ZN(new_n561));
  NOR2_X1   g136(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n562), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n509), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n563), .A2(KEYINPUT73), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT73), .B1(new_n563), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n558), .B1(new_n566), .B2(new_n567), .ZN(G299));
  NAND3_X1  g143(.A1(new_n519), .A2(new_n525), .A3(new_n530), .ZN(G286));
  NAND2_X1  g144(.A1(new_n509), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n553), .ZN(G288));
  NAND2_X1  g148(.A1(new_n509), .A2(G48), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n498), .B2(new_n499), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n515), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n574), .B(new_n579), .C1(new_n580), .C2(new_n553), .ZN(G305));
  NAND2_X1  g156(.A1(new_n509), .A2(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n582), .B1(new_n514), .B2(new_n583), .C1(new_n584), .C2(new_n553), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n506), .A2(KEYINPUT10), .A3(G92), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n553), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(new_n509), .B2(G54), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT74), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n586), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n586), .B1(new_n596), .B2(G868), .ZN(G321));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(G286), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n599), .ZN(G297));
  XOR2_X1   g177(.A(G297), .B(KEYINPUT75), .Z(G280));
  XOR2_X1   g178(.A(KEYINPUT76), .B(G559), .Z(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(G860), .B2(new_n604), .ZN(G148));
  NAND3_X1  g180(.A1(new_n540), .A2(new_n545), .A3(new_n544), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n596), .A2(new_n604), .ZN(new_n607));
  MUX2_X1   g182(.A(new_n606), .B(new_n607), .S(G868), .Z(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n465), .A2(G2104), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT12), .Z(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT13), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n477), .A2(G123), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n465), .A2(G135), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT77), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n617), .A2(KEYINPUT78), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(KEYINPUT78), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n618), .B(new_n619), .C1(G111), .C2(new_n475), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n614), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n613), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2430), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(KEYINPUT14), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT80), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XOR2_X1   g214(.A(G2443), .B(G2446), .Z(new_n640));
  XOR2_X1   g215(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n635), .A2(new_n636), .A3(new_n641), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n643), .A2(KEYINPUT81), .A3(G14), .A4(new_n644), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  INV_X1    g230(.A(new_n651), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(new_n653), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n656), .B2(new_n657), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n651), .A2(new_n653), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n652), .B1(new_n661), .B2(KEYINPUT17), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n655), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n622), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(G2100), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(G2100), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT82), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT83), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT20), .Z(new_n676));
  OR2_X1    g251(.A1(new_n669), .A2(new_n671), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n674), .A3(new_n672), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n678), .C1(new_n674), .C2(new_n677), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  NOR2_X1   g261(.A1(G29), .A2(G33), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT92), .Z(new_n688));
  AND2_X1   g263(.A1(new_n467), .A2(G103), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(KEYINPUT25), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(KEYINPUT25), .ZN(new_n691));
  AOI22_X1  g266(.A1(new_n690), .A2(new_n691), .B1(G139), .B2(new_n465), .ZN(new_n692));
  AOI22_X1  g267(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n475), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n688), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G2072), .ZN(new_n697));
  AND2_X1   g272(.A1(KEYINPUT24), .A2(G34), .ZN(new_n698));
  NOR2_X1   g273(.A1(KEYINPUT24), .A2(G34), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n695), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n473), .B2(new_n695), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G2084), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT93), .B1(G29), .B2(G32), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n467), .A2(G105), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT26), .ZN(new_n706));
  AOI211_X1 g281(.A(new_n704), .B(new_n706), .C1(G141), .C2(new_n465), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n477), .A2(G129), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G29), .ZN(new_n710));
  MUX2_X1   g285(.A(KEYINPUT93), .B(new_n703), .S(new_n710), .Z(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n697), .B(new_n702), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NOR2_X1   g289(.A1(G27), .A2(G29), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G164), .B2(G29), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT97), .B(G2078), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT31), .B(G11), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT30), .B(G28), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n695), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n621), .B2(new_n695), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT95), .Z(new_n724));
  NOR2_X1   g299(.A1(G16), .A2(G19), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n546), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1341), .ZN(new_n727));
  OR4_X1    g302(.A1(new_n713), .A2(new_n719), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G29), .A2(G35), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G162), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G5), .A2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT96), .Z(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(G301), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NOR2_X1   g315(.A1(G168), .A2(new_n736), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n736), .B2(G21), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n739), .B(new_n740), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT94), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n695), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n477), .A2(G128), .ZN(new_n749));
  MUX2_X1   g324(.A(G104), .B(G116), .S(G2105), .Z(new_n750));
  AOI22_X1  g325(.A1(G140), .A2(new_n465), .B1(new_n750), .B2(G2104), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n752), .A2(KEYINPUT91), .A3(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(KEYINPUT91), .B1(new_n752), .B2(G29), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n748), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n733), .A2(new_n744), .A3(new_n746), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G4), .A2(G16), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n596), .B2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1348), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n736), .A2(G20), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT23), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n601), .B2(new_n736), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT98), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR4_X1   g342(.A1(new_n728), .A2(new_n758), .A3(new_n761), .A4(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(G16), .A2(G22), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G303), .B2(new_n736), .ZN(new_n771));
  INV_X1    g346(.A(G1971), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  OR2_X1    g349(.A1(G16), .A2(G23), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G288), .B2(new_n736), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT33), .B(G1976), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT88), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n776), .A2(new_n779), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n773), .B(new_n774), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(G6), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G305), .B2(new_n736), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT86), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n520), .A2(G61), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n514), .B1(new_n787), .B2(new_n577), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G48), .B2(new_n509), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n506), .A2(G86), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n789), .A2(G16), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(KEYINPUT86), .B1(new_n791), .B2(new_n783), .ZN(new_n792));
  OAI21_X1  g367(.A(KEYINPUT87), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n784), .A2(new_n785), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(KEYINPUT86), .A3(new_n783), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT87), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n782), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n799), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n793), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n800), .A2(KEYINPUT89), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(KEYINPUT89), .B1(new_n800), .B2(new_n802), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT34), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n798), .A2(new_n799), .ZN(new_n808));
  INV_X1    g383(.A(new_n782), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n808), .A2(new_n802), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n800), .A2(KEYINPUT89), .A3(new_n802), .ZN(new_n813));
  AOI21_X1  g388(.A(KEYINPUT34), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n477), .A2(G119), .ZN(new_n815));
  MUX2_X1   g390(.A(G95), .B(G107), .S(G2105), .Z(new_n816));
  AOI22_X1  g391(.A1(G131), .A2(new_n465), .B1(new_n816), .B2(G2104), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G29), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G25), .B2(G29), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n821), .A2(KEYINPUT84), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(KEYINPUT84), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT35), .B(G1991), .Z(new_n824));
  NOR3_X1   g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n824), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n821), .A2(KEYINPUT84), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n821), .A2(KEYINPUT84), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n736), .A2(G24), .ZN(new_n831));
  XOR2_X1   g406(.A(G290), .B(KEYINPUT85), .Z(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n736), .ZN(new_n833));
  INV_X1    g408(.A(G1986), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT90), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n814), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n805), .B1(new_n803), .B2(new_n804), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n830), .A2(new_n835), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT90), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n807), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n837), .B1(new_n814), .B2(new_n836), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT90), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT36), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n807), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n769), .B1(new_n843), .B2(new_n848), .ZN(G311));
  AOI21_X1  g424(.A(new_n847), .B1(new_n846), .B2(new_n807), .ZN(new_n850));
  AOI211_X1 g425(.A(KEYINPUT36), .B(new_n806), .C1(new_n844), .C2(new_n845), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n768), .B1(new_n850), .B2(new_n851), .ZN(G150));
  NAND2_X1  g427(.A1(new_n509), .A2(G55), .ZN(new_n853));
  OAI211_X1 g428(.A(G93), .B(new_n520), .C1(new_n524), .C2(new_n501), .ZN(new_n854));
  INV_X1    g429(.A(G67), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n498), .B2(new_n499), .ZN(new_n856));
  AND2_X1   g431(.A1(G80), .A2(G543), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n515), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT99), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n853), .A2(new_n861), .A3(new_n854), .A4(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n596), .A2(G559), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n860), .A2(new_n606), .A3(new_n862), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n546), .A2(new_n859), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n867), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(G860), .B1(new_n872), .B2(new_n873), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n874), .A2(KEYINPUT100), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT100), .B1(new_n874), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n865), .B1(new_n876), .B2(new_n877), .ZN(G145));
  NOR2_X1   g453(.A1(new_n819), .A2(new_n611), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n465), .A2(G142), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n882));
  OAI22_X1  g457(.A1(new_n881), .A2(KEYINPUT102), .B1(G118), .B2(new_n475), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n477), .B2(G130), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n611), .A2(new_n815), .A3(new_n817), .ZN(new_n886));
  OR3_X1    g461(.A1(new_n879), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n879), .B2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n490), .B(new_n493), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n476), .A2(G126), .ZN(new_n891));
  INV_X1    g466(.A(new_n485), .ZN(new_n892));
  XNOR2_X1  g467(.A(KEYINPUT70), .B(G114), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(G2105), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n894), .B2(new_n466), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT101), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n487), .A2(new_n897), .A3(new_n495), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n752), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n889), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n887), .A2(new_n888), .A3(new_n900), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n709), .B(new_n694), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G162), .B(new_n473), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n621), .ZN(new_n908));
  INV_X1    g483(.A(new_n905), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n902), .A2(new_n903), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n908), .B1(new_n906), .B2(new_n910), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g491(.A(G290), .B(G288), .ZN(new_n917));
  XNOR2_X1  g492(.A(G303), .B(G305), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n917), .B(new_n918), .Z(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n607), .A2(new_n871), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n596), .A2(new_n604), .A3(new_n870), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(G543), .B1(new_n524), .B2(new_n501), .ZN(new_n924));
  INV_X1    g499(.A(G54), .ZN(new_n925));
  OAI22_X1  g500(.A1(new_n924), .A2(new_n925), .B1(new_n592), .B2(new_n556), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n590), .B2(new_n587), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n927), .B(new_n558), .C1(new_n566), .C2(new_n567), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT73), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n561), .A2(new_n562), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n564), .B1(new_n509), .B2(new_n560), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT73), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n927), .B1(new_n935), .B2(new_n558), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n923), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT41), .B1(new_n929), .B2(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(G299), .A2(new_n595), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n928), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n921), .A3(new_n922), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n938), .A2(new_n939), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n939), .B1(new_n938), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n920), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n938), .A2(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n938), .A2(new_n939), .A3(new_n945), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n919), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G868), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n863), .A2(G868), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT103), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n599), .B1(new_n948), .B2(new_n952), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n958), .A2(new_n959), .A3(new_n955), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n957), .A2(new_n960), .ZN(G295));
  NOR2_X1   g536(.A1(new_n958), .A2(new_n955), .ZN(G331));
  NAND3_X1  g537(.A1(G286), .A2(G301), .A3(KEYINPUT104), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n532), .A2(new_n964), .A3(new_n533), .A4(new_n537), .ZN(new_n965));
  NAND2_X1  g540(.A1(G168), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n533), .A2(new_n537), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n967), .B2(new_n532), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n963), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(new_n869), .A3(new_n868), .ZN(new_n970));
  NAND2_X1  g545(.A1(G301), .A2(KEYINPUT104), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(G168), .A3(new_n965), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n870), .A2(new_n972), .A3(new_n963), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n937), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n970), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n941), .A2(new_n942), .A3(new_n928), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n942), .B1(new_n941), .B2(new_n928), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT105), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n944), .A2(new_n981), .A3(new_n976), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n975), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(G37), .B1(new_n983), .B2(new_n920), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT106), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n976), .B1(new_n940), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n974), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n919), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n983), .A2(new_n920), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(KEYINPUT43), .A3(new_n984), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT44), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n984), .B2(new_n989), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n979), .A2(KEYINPUT105), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n981), .B1(new_n944), .B2(new_n976), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n920), .B(new_n974), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  AND4_X1   g575(.A1(new_n996), .A2(new_n1000), .A3(new_n989), .A4(new_n912), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT43), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n993), .A2(new_n991), .A3(new_n984), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n995), .B1(new_n1004), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g580(.A(G1384), .B1(new_n487), .B2(new_n495), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT109), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n890), .B2(new_n895), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT108), .B(G40), .Z(new_n1014));
  AND3_X1   g589(.A1(new_n468), .A2(new_n472), .A3(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n896), .A2(KEYINPUT45), .A3(new_n1008), .A4(new_n898), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT56), .B(G2072), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n557), .A2(new_n1019), .ZN(new_n1020));
  OAI221_X1 g595(.A(KEYINPUT117), .B1(new_n555), .B2(new_n556), .C1(new_n553), .C2(new_n554), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT57), .ZN(new_n1023));
  AOI22_X1  g598(.A1(G299), .A2(KEYINPUT57), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT50), .B1(new_n496), .B2(new_n1008), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  AOI211_X1 g601(.A(new_n1026), .B(G1384), .C1(new_n487), .C2(new_n495), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1015), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n766), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1018), .A2(new_n1024), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1024), .B1(new_n1018), .B2(new_n1029), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n927), .B(KEYINPUT74), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1015), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(new_n1009), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n756), .ZN(new_n1035));
  INV_X1    g610(.A(G1348), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1032), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1030), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT60), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1009), .A2(new_n1026), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1006), .A2(KEYINPUT50), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1035), .B1(new_n1045), .B2(G1348), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n596), .B1(new_n1046), .B2(KEYINPUT60), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1047), .A2(new_n1038), .A3(new_n1048), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1028), .A2(new_n1036), .B1(new_n1034), .B2(new_n756), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1032), .B1(new_n1050), .B2(new_n1042), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n596), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT121), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1042), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1048), .B1(new_n1047), .B2(new_n1038), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(KEYINPUT121), .A3(new_n1052), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1030), .A2(KEYINPUT120), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1018), .A2(new_n1024), .A3(new_n1060), .A4(new_n1029), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT61), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1031), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1010), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1006), .A2(KEYINPUT109), .A3(KEYINPUT45), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1015), .B(new_n1016), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT58), .B(G1341), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1068), .A2(G1996), .B1(new_n1034), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n546), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n546), .A3(new_n1072), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1030), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1063), .B1(new_n1077), .B2(new_n1031), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1065), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1041), .B1(new_n1058), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G8), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1976), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G288), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT52), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n1084), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1087), .B(new_n1082), .C1(new_n1084), .C2(G288), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(G1981), .B1(new_n788), .B2(KEYINPUT112), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n789), .A2(new_n790), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1981), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n579), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G305), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT49), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(KEYINPUT113), .A3(new_n1097), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1091), .A2(new_n1095), .A3(KEYINPUT49), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1103), .A2(new_n1082), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1089), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(G303), .A2(G8), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT55), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1016), .A2(new_n1015), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n772), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n732), .B(new_n1015), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1081), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1105), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT110), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1117), .A2(KEYINPUT110), .A3(new_n732), .A4(new_n1015), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(KEYINPUT111), .A3(new_n1111), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G8), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT111), .B1(new_n1119), .B2(new_n1111), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1114), .B1(new_n1123), .B2(new_n1108), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  NOR2_X1   g700(.A1(G168), .A2(new_n1081), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1015), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1015), .B(KEYINPUT115), .C1(new_n1006), .C2(KEYINPUT45), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n743), .ZN(new_n1136));
  INV_X1    g711(.A(G2084), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1045), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(G8), .B(new_n1129), .C1(new_n1139), .C2(G286), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1126), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1135), .A2(new_n743), .B1(new_n1137), .B2(new_n1045), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1141), .B(new_n1128), .C1(new_n1142), .C2(new_n1081), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(G8), .A3(G286), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT53), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1068), .B2(G2078), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1028), .A2(new_n738), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1146), .A2(G2078), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(G301), .B(KEYINPUT54), .Z(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1011), .B1(new_n899), .B2(G1384), .ZN(new_n1154));
  AND3_X1   g729(.A1(G160), .A2(G40), .A3(new_n1149), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1016), .A3(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1156), .A2(new_n1148), .A3(new_n1152), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1151), .A2(new_n1153), .B1(new_n1147), .B2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1124), .A2(KEYINPUT123), .A3(new_n1145), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1145), .A2(new_n1158), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1119), .A2(new_n1111), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT111), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1164), .A2(G8), .A3(new_n1108), .A4(new_n1120), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT113), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1099), .B(KEYINPUT49), .C1(new_n1091), .C2(new_n1095), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1104), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(G8), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1170), .B1(new_n1172), .B2(new_n1107), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1165), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1160), .B1(new_n1161), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1080), .A2(new_n1159), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1168), .ZN(new_n1177));
  OR2_X1    g752(.A1(G288), .A2(G1976), .ZN(new_n1178));
  OAI22_X1  g753(.A1(new_n1177), .A2(new_n1178), .B1(G1981), .B2(G305), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1082), .B(KEYINPUT114), .Z(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n1183));
  AND4_X1   g758(.A1(new_n1183), .A2(new_n1140), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1151), .A2(G171), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1165), .A2(new_n1173), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1145), .A2(KEYINPUT62), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1182), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT116), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1116), .A2(new_n1118), .B1(new_n1068), .B2(new_n772), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1081), .B1(new_n1191), .B2(KEYINPUT111), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1108), .B1(new_n1192), .B2(new_n1164), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1190), .B1(new_n1193), .B2(new_n1170), .ZN(new_n1194));
  OAI211_X1 g769(.A(KEYINPUT116), .B(new_n1105), .C1(new_n1123), .C2(new_n1108), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1142), .A2(new_n1081), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1196), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n1123), .B2(new_n1108), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1194), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1196), .A2(G168), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1200), .B1(new_n1174), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1176), .A2(new_n1189), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(G1996), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n709), .B(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n752), .B(G2067), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n818), .B(new_n826), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(G290), .B(new_n834), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1154), .A2(new_n1033), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1204), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT48), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1213), .ZN(new_n1217));
  OR3_X1    g792(.A1(new_n1217), .A2(G1986), .A3(G290), .ZN(new_n1218));
  OAI22_X1  g793(.A1(new_n1216), .A2(new_n1218), .B1(new_n1210), .B2(new_n1217), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1219), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1220));
  INV_X1    g795(.A(new_n709), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1213), .B1(new_n1221), .B2(new_n1207), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n1223));
  OAI211_X1 g798(.A(new_n1213), .B(new_n1205), .C1(new_n1223), .C2(KEYINPUT46), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1223), .A2(KEYINPUT46), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1222), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1226), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1227), .B(KEYINPUT47), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n819), .A2(new_n824), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n1229), .B(KEYINPUT124), .ZN(new_n1230));
  OAI22_X1  g805(.A1(new_n1208), .A2(new_n1230), .B1(G2067), .B2(new_n752), .ZN(new_n1231));
  AOI211_X1 g806(.A(new_n1220), .B(new_n1228), .C1(new_n1213), .C2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1215), .A2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g808(.A(new_n685), .B1(new_n913), .B2(new_n914), .ZN(new_n1235));
  NOR2_X1   g809(.A1(G227), .A2(new_n461), .ZN(new_n1236));
  INV_X1    g810(.A(new_n1236), .ZN(new_n1237));
  OAI21_X1  g811(.A(KEYINPUT126), .B1(G401), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n1239));
  NAND3_X1  g813(.A1(new_n649), .A2(new_n1239), .A3(new_n1236), .ZN(new_n1240));
  AOI21_X1  g814(.A(new_n1235), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  AND2_X1   g815(.A1(new_n992), .A2(new_n994), .ZN(new_n1242));
  AND2_X1   g816(.A1(new_n1241), .A2(new_n1242), .ZN(G308));
  NAND2_X1  g817(.A1(new_n1241), .A2(new_n1242), .ZN(G225));
endmodule


