

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  XNOR2_X1 U323 ( .A(n368), .B(KEYINPUT96), .ZN(n370) );
  NOR2_X1 U324 ( .A1(n476), .A2(n521), .ZN(n578) );
  XNOR2_X1 U325 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U326 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U327 ( .A(n477), .B(KEYINPUT28), .Z(n537) );
  XOR2_X1 U328 ( .A(n308), .B(n307), .Z(n309) );
  XOR2_X1 U329 ( .A(G169GAT), .B(n347), .Z(n291) );
  XOR2_X1 U330 ( .A(G85GAT), .B(G92GAT), .Z(n292) );
  INV_X1 U331 ( .A(KEYINPUT46), .ZN(n457) );
  XNOR2_X1 U332 ( .A(n457), .B(KEYINPUT111), .ZN(n458) );
  XNOR2_X1 U333 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U334 ( .A(n464), .B(KEYINPUT66), .ZN(n465) );
  XNOR2_X1 U335 ( .A(n466), .B(n465), .ZN(n469) );
  INV_X1 U336 ( .A(n521), .ZN(n369) );
  NAND2_X1 U337 ( .A1(n578), .A2(n477), .ZN(n478) );
  AND2_X1 U338 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U339 ( .A(KEYINPUT26), .B(n364), .ZN(n577) );
  XNOR2_X1 U340 ( .A(n448), .B(n447), .ZN(n456) );
  XNOR2_X1 U341 ( .A(n393), .B(n392), .ZN(n560) );
  NOR2_X1 U342 ( .A1(n520), .A2(n489), .ZN(n450) );
  INV_X1 U343 ( .A(G43GAT), .ZN(n451) );
  XNOR2_X1 U344 ( .A(n450), .B(KEYINPUT38), .ZN(n504) );
  XNOR2_X1 U345 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U346 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U347 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(G183GAT), .B(KEYINPUT18), .Z(n294) );
  XNOR2_X1 U350 ( .A(KEYINPUT17), .B(KEYINPUT84), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n296) );
  XOR2_X1 U352 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n295) );
  XOR2_X1 U353 ( .A(n296), .B(n295), .Z(n335) );
  XOR2_X1 U354 ( .A(G176GAT), .B(KEYINPUT20), .Z(n298) );
  XNOR2_X1 U355 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n297) );
  XNOR2_X1 U356 ( .A(n298), .B(n297), .ZN(n308) );
  INV_X1 U357 ( .A(G190GAT), .ZN(n481) );
  XOR2_X1 U358 ( .A(G190GAT), .B(G134GAT), .Z(n300) );
  XOR2_X1 U359 ( .A(G120GAT), .B(G71GAT), .Z(n444) );
  XOR2_X1 U360 ( .A(G15GAT), .B(G127GAT), .Z(n399) );
  XNOR2_X1 U361 ( .A(n444), .B(n399), .ZN(n299) );
  XNOR2_X1 U362 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U363 ( .A(n301), .B(G99GAT), .Z(n306) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U365 ( .A(n302), .B(KEYINPUT82), .ZN(n347) );
  NAND2_X1 U366 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U367 ( .A(n291), .B(n303), .ZN(n304) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(n304), .ZN(n305) );
  XNOR2_X1 U369 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X2 U370 ( .A(n335), .B(n309), .Z(n535) );
  XOR2_X1 U371 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n311) );
  XNOR2_X1 U372 ( .A(G218GAT), .B(G106GAT), .ZN(n310) );
  XNOR2_X1 U373 ( .A(n311), .B(n310), .ZN(n326) );
  XOR2_X1 U374 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n313) );
  NAND2_X1 U375 ( .A1(G228GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U376 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U377 ( .A(n314), .B(KEYINPUT90), .Z(n320) );
  XOR2_X1 U378 ( .A(G211GAT), .B(KEYINPUT21), .Z(n316) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n315) );
  XNOR2_X1 U380 ( .A(n316), .B(n315), .ZN(n331) );
  XOR2_X1 U381 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n318) );
  XNOR2_X1 U382 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n318), .B(n317), .ZN(n350) );
  XNOR2_X1 U384 ( .A(n331), .B(n350), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n320), .B(n319), .ZN(n322) );
  XNOR2_X1 U386 ( .A(G78GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U387 ( .A(n321), .B(G148GAT), .ZN(n437) );
  XOR2_X1 U388 ( .A(n322), .B(n437), .Z(n324) );
  XOR2_X1 U389 ( .A(G50GAT), .B(G162GAT), .Z(n382) );
  XOR2_X1 U390 ( .A(G22GAT), .B(G155GAT), .Z(n400) );
  XNOR2_X1 U391 ( .A(n382), .B(n400), .ZN(n323) );
  XNOR2_X1 U392 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U393 ( .A(n326), .B(n325), .Z(n477) );
  XOR2_X1 U394 ( .A(KEYINPUT93), .B(G92GAT), .Z(n328) );
  NAND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U396 ( .A(n328), .B(n327), .ZN(n330) );
  XNOR2_X1 U397 ( .A(G36GAT), .B(G190GAT), .ZN(n329) );
  XNOR2_X1 U398 ( .A(n329), .B(G218GAT), .ZN(n374) );
  XOR2_X1 U399 ( .A(n330), .B(n374), .Z(n333) );
  XNOR2_X1 U400 ( .A(n331), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U401 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U402 ( .A(G176GAT), .B(G64GAT), .Z(n443) );
  XOR2_X1 U403 ( .A(n334), .B(n443), .Z(n338) );
  XOR2_X1 U404 ( .A(G169GAT), .B(G8GAT), .Z(n428) );
  INV_X1 U405 ( .A(n335), .ZN(n336) );
  XOR2_X1 U406 ( .A(n428), .B(n336), .Z(n337) );
  XOR2_X1 U407 ( .A(n338), .B(n337), .Z(n523) );
  XNOR2_X1 U408 ( .A(n523), .B(KEYINPUT27), .ZN(n365) );
  XOR2_X1 U409 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n340) );
  XNOR2_X1 U410 ( .A(KEYINPUT92), .B(KEYINPUT6), .ZN(n339) );
  XNOR2_X1 U411 ( .A(n340), .B(n339), .ZN(n358) );
  XOR2_X1 U412 ( .A(G155GAT), .B(G162GAT), .Z(n342) );
  XNOR2_X1 U413 ( .A(G120GAT), .B(G127GAT), .ZN(n341) );
  XNOR2_X1 U414 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U415 ( .A(KEYINPUT1), .B(G57GAT), .Z(n344) );
  XNOR2_X1 U416 ( .A(G1GAT), .B(G148GAT), .ZN(n343) );
  XNOR2_X1 U417 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U418 ( .A(n346), .B(n345), .Z(n356) );
  XOR2_X1 U419 ( .A(KEYINPUT5), .B(n347), .Z(n349) );
  NAND2_X1 U420 ( .A1(G225GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U421 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U422 ( .A(G134GAT), .B(KEYINPUT74), .Z(n373) );
  XOR2_X1 U423 ( .A(n373), .B(G85GAT), .Z(n352) );
  XNOR2_X1 U424 ( .A(G29GAT), .B(n350), .ZN(n351) );
  XNOR2_X1 U425 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U427 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n521) );
  NAND2_X1 U429 ( .A1(n365), .A2(n521), .ZN(n533) );
  NOR2_X1 U430 ( .A1(n537), .A2(n533), .ZN(n359) );
  XOR2_X1 U431 ( .A(KEYINPUT94), .B(n359), .Z(n360) );
  NOR2_X1 U432 ( .A1(n535), .A2(n360), .ZN(n372) );
  NAND2_X1 U433 ( .A1(n535), .A2(n523), .ZN(n361) );
  NAND2_X1 U434 ( .A1(n477), .A2(n361), .ZN(n362) );
  XOR2_X1 U435 ( .A(KEYINPUT25), .B(n362), .Z(n367) );
  NOR2_X1 U436 ( .A1(n535), .A2(n477), .ZN(n363) );
  XOR2_X1 U437 ( .A(KEYINPUT95), .B(n363), .Z(n364) );
  NAND2_X1 U438 ( .A1(n365), .A2(n577), .ZN(n366) );
  NAND2_X1 U439 ( .A1(n367), .A2(n366), .ZN(n368) );
  NOR2_X1 U440 ( .A1(n372), .A2(n371), .ZN(n488) );
  XNOR2_X1 U441 ( .A(n374), .B(n373), .ZN(n378) );
  INV_X1 U442 ( .A(n378), .ZN(n376) );
  AND2_X1 U443 ( .A1(G232GAT), .A2(G233GAT), .ZN(n377) );
  INV_X1 U444 ( .A(n377), .ZN(n375) );
  NAND2_X1 U445 ( .A1(n376), .A2(n375), .ZN(n380) );
  NAND2_X1 U446 ( .A1(n378), .A2(n377), .ZN(n379) );
  NAND2_X1 U447 ( .A1(n380), .A2(n379), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n381), .B(KEYINPUT73), .ZN(n384) );
  XOR2_X1 U449 ( .A(n382), .B(KEYINPUT9), .Z(n383) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n393) );
  XOR2_X1 U451 ( .A(G29GAT), .B(G43GAT), .Z(n386) );
  XNOR2_X1 U452 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n386), .B(n385), .ZN(n431) );
  XNOR2_X1 U454 ( .A(G99GAT), .B(G106GAT), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n292), .B(n387), .ZN(n438) );
  XOR2_X1 U456 ( .A(n431), .B(n438), .Z(n391) );
  XOR2_X1 U457 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n389) );
  XNOR2_X1 U458 ( .A(KEYINPUT64), .B(KEYINPUT11), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U460 ( .A(KEYINPUT75), .B(n560), .Z(n545) );
  XNOR2_X1 U461 ( .A(KEYINPUT36), .B(n545), .ZN(n463) );
  XOR2_X1 U462 ( .A(G78GAT), .B(G211GAT), .Z(n395) );
  XNOR2_X1 U463 ( .A(G183GAT), .B(G71GAT), .ZN(n394) );
  XNOR2_X1 U464 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U465 ( .A(KEYINPUT13), .B(G57GAT), .Z(n441) );
  XOR2_X1 U466 ( .A(n396), .B(n441), .Z(n398) );
  XNOR2_X1 U467 ( .A(G8GAT), .B(G64GAT), .ZN(n397) );
  XNOR2_X1 U468 ( .A(n398), .B(n397), .ZN(n413) );
  XOR2_X1 U469 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U470 ( .A1(G231GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U471 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U472 ( .A(KEYINPUT80), .B(KEYINPUT76), .Z(n404) );
  XNOR2_X1 U473 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U475 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U476 ( .A(KEYINPUT68), .B(G1GAT), .Z(n430) );
  XOR2_X1 U477 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n408) );
  XNOR2_X1 U478 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n407) );
  XNOR2_X1 U479 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U480 ( .A(n430), .B(n409), .ZN(n410) );
  XNOR2_X1 U481 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U482 ( .A(n413), .B(n412), .Z(n587) );
  INV_X1 U483 ( .A(n587), .ZN(n573) );
  NAND2_X1 U484 ( .A1(n463), .A2(n573), .ZN(n414) );
  NOR2_X1 U485 ( .A1(n488), .A2(n414), .ZN(n416) );
  XNOR2_X1 U486 ( .A(KEYINPUT37), .B(KEYINPUT100), .ZN(n415) );
  XNOR2_X1 U487 ( .A(n416), .B(n415), .ZN(n520) );
  XOR2_X1 U488 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n418) );
  NAND2_X1 U489 ( .A1(G229GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U490 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U491 ( .A(n419), .B(KEYINPUT30), .Z(n427) );
  XOR2_X1 U492 ( .A(G15GAT), .B(G113GAT), .Z(n421) );
  XNOR2_X1 U493 ( .A(G50GAT), .B(G36GAT), .ZN(n420) );
  XNOR2_X1 U494 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U495 ( .A(KEYINPUT67), .B(G141GAT), .Z(n423) );
  XNOR2_X1 U496 ( .A(G197GAT), .B(G22GAT), .ZN(n422) );
  XNOR2_X1 U497 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U498 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U499 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U500 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U501 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U502 ( .A(n433), .B(n432), .ZN(n579) );
  XNOR2_X1 U503 ( .A(KEYINPUT32), .B(KEYINPUT70), .ZN(n435) );
  AND2_X1 U504 ( .A1(G230GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U505 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U506 ( .A(n436), .B(KEYINPUT71), .Z(n440) );
  XNOR2_X1 U507 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U508 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U509 ( .A(n442), .B(n441), .Z(n448) );
  XNOR2_X1 U510 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U511 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n445) );
  INV_X1 U512 ( .A(n456), .ZN(n467) );
  NOR2_X1 U513 ( .A1(n579), .A2(n456), .ZN(n449) );
  XOR2_X1 U514 ( .A(KEYINPUT72), .B(n449), .Z(n489) );
  NAND2_X1 U515 ( .A1(n504), .A2(n535), .ZN(n454) );
  XOR2_X1 U516 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n452) );
  INV_X1 U517 ( .A(n523), .ZN(n473) );
  INV_X1 U518 ( .A(KEYINPUT41), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n456), .B(n455), .ZN(n508) );
  INV_X1 U520 ( .A(n508), .ZN(n567) );
  NOR2_X1 U521 ( .A1(n579), .A2(n567), .ZN(n459) );
  NOR2_X1 U522 ( .A1(n460), .A2(n560), .ZN(n461) );
  NAND2_X1 U523 ( .A1(n461), .A2(n573), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(KEYINPUT47), .ZN(n471) );
  NAND2_X1 U525 ( .A1(n587), .A2(n463), .ZN(n466) );
  XOR2_X1 U526 ( .A(KEYINPUT112), .B(KEYINPUT45), .Z(n464) );
  AND2_X1 U527 ( .A1(n579), .A2(n467), .ZN(n468) );
  AND2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT48), .ZN(n534) );
  NOR2_X1 U531 ( .A1(n473), .A2(n534), .ZN(n475) );
  XNOR2_X1 U532 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n478), .B(KEYINPUT55), .ZN(n479) );
  NAND2_X1 U535 ( .A1(n479), .A2(n535), .ZN(n480) );
  XOR2_X1 U536 ( .A(KEYINPUT120), .B(n480), .Z(n566) );
  NAND2_X1 U537 ( .A1(n545), .A2(n566), .ZN(n484) );
  XOR2_X1 U538 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n482) );
  XOR2_X1 U539 ( .A(KEYINPUT97), .B(KEYINPUT34), .Z(n491) );
  NOR2_X1 U540 ( .A1(n545), .A2(n573), .ZN(n486) );
  XNOR2_X1 U541 ( .A(KEYINPUT16), .B(KEYINPUT81), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n486), .B(n485), .ZN(n487) );
  OR2_X1 U543 ( .A1(n488), .A2(n487), .ZN(n509) );
  NOR2_X1 U544 ( .A1(n489), .A2(n509), .ZN(n497) );
  NAND2_X1 U545 ( .A1(n497), .A2(n521), .ZN(n490) );
  XNOR2_X1 U546 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n492), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n523), .A2(n497), .ZN(n493) );
  XNOR2_X1 U549 ( .A(n493), .B(KEYINPUT98), .ZN(n494) );
  XNOR2_X1 U550 ( .A(G8GAT), .B(n494), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U552 ( .A1(n497), .A2(n535), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NAND2_X1 U554 ( .A1(n497), .A2(n537), .ZN(n498) );
  XNOR2_X1 U555 ( .A(n498), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT39), .ZN(n502) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT101), .Z(n500) );
  NAND2_X1 U558 ( .A1(n504), .A2(n521), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n504), .A2(n523), .ZN(n503) );
  XNOR2_X1 U562 ( .A(n503), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n506) );
  NAND2_X1 U564 ( .A1(n537), .A2(n504), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n507), .ZN(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT42), .B(KEYINPUT105), .Z(n511) );
  NAND2_X1 U568 ( .A1(n579), .A2(n508), .ZN(n519) );
  NOR2_X1 U569 ( .A1(n519), .A2(n509), .ZN(n515) );
  NAND2_X1 U570 ( .A1(n515), .A2(n521), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n523), .A2(n515), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n513), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n515), .A2(n535), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U578 ( .A1(n515), .A2(n537), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n520), .A2(n519), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n529), .A2(n521), .ZN(n522) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  XOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT107), .Z(n525) );
  NAND2_X1 U585 ( .A1(n529), .A2(n523), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n525), .B(n524), .ZN(G1337GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n527) );
  NAND2_X1 U588 ( .A1(n529), .A2(n535), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n528), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n531) );
  NAND2_X1 U592 ( .A1(n529), .A2(n537), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n532), .Z(G1339GAT) );
  NOR2_X1 U595 ( .A1(n534), .A2(n533), .ZN(n550) );
  NAND2_X1 U596 ( .A1(n535), .A2(n550), .ZN(n536) );
  XOR2_X1 U597 ( .A(n536), .B(KEYINPUT113), .Z(n538) );
  NOR2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n546) );
  INV_X1 U599 ( .A(n546), .ZN(n542) );
  NOR2_X1 U600 ( .A1(n579), .A2(n542), .ZN(n539) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n539), .Z(G1340GAT) );
  NOR2_X1 U602 ( .A1(n567), .A2(n542), .ZN(n541) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NOR2_X1 U605 ( .A1(n573), .A2(n542), .ZN(n543) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(n543), .Z(n544) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n548) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n577), .A2(n550), .ZN(n551) );
  XNOR2_X1 U613 ( .A(KEYINPUT115), .B(n551), .ZN(n561) );
  INV_X1 U614 ( .A(n561), .ZN(n558) );
  NOR2_X1 U615 ( .A1(n579), .A2(n558), .ZN(n552) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  NOR2_X1 U617 ( .A1(n567), .A2(n558), .ZN(n557) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n554) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT52), .B(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n573), .A2(n558), .ZN(n559) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT118), .ZN(n563) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n563), .ZN(G1347GAT) );
  INV_X1 U628 ( .A(n579), .ZN(n564) );
  AND2_X1 U629 ( .A1(n566), .A2(n564), .ZN(n565) );
  XOR2_X1 U630 ( .A(n565), .B(G169GAT), .Z(G1348GAT) );
  INV_X1 U631 ( .A(n566), .ZN(n574) );
  NOR2_X1 U632 ( .A1(n574), .A2(n567), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n569) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT56), .B(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  NOR2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U639 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1350GAT) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n584) );
  NOR2_X1 U642 ( .A1(n579), .A2(n584), .ZN(n581) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n581), .B(n580), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n582) );
  XNOR2_X1 U646 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  INV_X1 U648 ( .A(n584), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n589), .A2(n456), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n589), .A2(n587), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n591) );
  NAND2_X1 U654 ( .A1(n589), .A2(n463), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(G218GAT), .B(n592), .Z(G1355GAT) );
endmodule

