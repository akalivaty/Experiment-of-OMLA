//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n205), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n208), .B(new_n214), .C1(new_n221), .C2(KEYINPUT1), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0023(.A(G238), .B(G244), .Z(new_n224));
  XNOR2_X1  g0024(.A(G226), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XOR2_X1   g0032(.A(G87), .B(G97), .Z(new_n233));
  XOR2_X1   g0033(.A(G107), .B(G116), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G351));
  INV_X1    g0041(.A(G1), .ZN(new_n242));
  NAND3_X1  g0042(.A1(new_n242), .A2(G13), .A3(G20), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(KEYINPUT69), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT69), .ZN(new_n245));
  NAND4_X1  g0045(.A1(new_n245), .A2(new_n242), .A3(G13), .A4(G20), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n211), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(new_n212), .B2(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n242), .A2(KEYINPUT70), .A3(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G50), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n244), .A2(new_n246), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n252), .A2(new_n259), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n262));
  INV_X1    g0062(.A(G150), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n212), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT8), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G58), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT68), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT67), .B(G58), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n267), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n264), .A2(G20), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n266), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n261), .B1(new_n275), .B2(new_n250), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT9), .ZN(new_n277));
  INV_X1    g0077(.A(G200), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G222), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G77), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(G1698), .ZN(new_n283));
  INV_X1    g0083(.A(G223), .ZN(new_n284));
  OAI221_X1 g0084(.A(new_n281), .B1(new_n282), .B2(new_n279), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n211), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(G274), .B1(new_n286), .B2(new_n211), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n287), .A2(new_n291), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(G226), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n278), .B1(new_n288), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n288), .A2(new_n296), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(G190), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n277), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n301));
  OR2_X1    g0101(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT71), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n298), .A2(G169), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n275), .A2(new_n250), .ZN(new_n306));
  INV_X1    g0106(.A(new_n261), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n304), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  OAI221_X1 g0109(.A(KEYINPUT71), .B1(new_n306), .B2(new_n307), .C1(G169), .C2(new_n298), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n298), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n277), .A2(new_n299), .A3(KEYINPUT72), .A4(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n303), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G68), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n254), .B2(new_n255), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n247), .A2(new_n250), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n247), .A2(new_n317), .A3(new_n250), .A4(KEYINPUT74), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n212), .A2(G33), .A3(G77), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n322), .B1(new_n212), .B2(G68), .C1(new_n265), .C2(new_n258), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n249), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT11), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT11), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n326), .A3(new_n249), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n320), .A2(new_n321), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n247), .B2(G68), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT76), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n329), .C1(new_n247), .C2(G68), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n260), .A2(new_n316), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n331), .B(new_n333), .C1(KEYINPUT12), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT77), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n328), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n328), .B2(new_n335), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT14), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n279), .A2(G226), .A3(new_n280), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n287), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n294), .B1(G238), .B2(new_n295), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n340), .B(G169), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n345), .A2(new_n346), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT13), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G179), .A3(new_n348), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n348), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n340), .B1(new_n356), .B2(G169), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n339), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n328), .A2(new_n335), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n349), .A2(new_n350), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(G190), .ZN(new_n361));
  OAI211_X1 g0161(.A(KEYINPUT73), .B(G200), .C1(new_n349), .C2(new_n350), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT73), .B1(new_n356), .B2(G200), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n279), .A2(G232), .A3(new_n280), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT3), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G33), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G107), .ZN(new_n372));
  INV_X1    g0172(.A(G238), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n367), .B(new_n372), .C1(new_n283), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n287), .ZN(new_n375));
  INV_X1    g0175(.A(G274), .ZN(new_n376));
  INV_X1    g0176(.A(new_n211), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G41), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n291), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n378), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n292), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G244), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G169), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G20), .A2(G77), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT8), .B(G58), .ZN(new_n389));
  INV_X1    g0189(.A(new_n274), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n388), .B1(new_n389), .B2(new_n265), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(new_n249), .B1(new_n282), .B2(new_n260), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n252), .A2(G77), .A3(new_n256), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n386), .A2(new_n387), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n384), .B1(new_n374), .B2(new_n287), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n311), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n386), .A2(G200), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n375), .A2(G190), .A3(new_n385), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n394), .A4(new_n393), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n315), .A2(new_n366), .A3(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n295), .A2(G232), .B1(new_n379), .B2(new_n291), .ZN(new_n404));
  INV_X1    g0204(.A(G87), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n264), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n368), .ZN(new_n407));
  AND2_X1   g0207(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n408));
  NOR2_X1   g0208(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n407), .B1(new_n410), .B2(G33), .ZN(new_n411));
  MUX2_X1   g0211(.A(G223), .B(G226), .S(G1698), .Z(new_n412));
  AOI21_X1  g0212(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(G179), .B(new_n404), .C1(new_n413), .C2(new_n381), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT78), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n369), .ZN(new_n416));
  NAND2_X1  g0216(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(G33), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n412), .A2(new_n418), .A3(new_n368), .ZN(new_n419));
  INV_X1    g0219(.A(new_n406), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n381), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G232), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n380), .B1(new_n382), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(G169), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n414), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n271), .A2(G68), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n202), .ZN(new_n427));
  INV_X1    g0227(.A(new_n265), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n427), .A2(G20), .B1(G159), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(new_n368), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT7), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n212), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G68), .ZN(new_n433));
  AOI21_X1  g0233(.A(G20), .B1(new_n418), .B2(new_n368), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n431), .ZN(new_n435));
  OAI211_X1 g0235(.A(KEYINPUT16), .B(new_n429), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT16), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n431), .A2(G20), .ZN(new_n438));
  AOI21_X1  g0238(.A(G33), .B1(new_n416), .B2(new_n417), .ZN(new_n439));
  INV_X1    g0239(.A(new_n370), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n431), .B1(new_n279), .B2(G20), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n316), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n428), .A2(G159), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n201), .B1(new_n271), .B2(G68), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n212), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n437), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n436), .A2(new_n249), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n270), .A2(new_n272), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n257), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(new_n252), .B1(new_n260), .B2(new_n449), .ZN(new_n451));
  AOI211_X1 g0251(.A(KEYINPUT18), .B(new_n425), .C1(new_n448), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT18), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n448), .A2(new_n451), .ZN(new_n454));
  INV_X1    g0254(.A(new_n425), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(G190), .B(new_n404), .C1(new_n413), .C2(new_n381), .ZN(new_n458));
  OAI21_X1  g0258(.A(G200), .B1(new_n421), .B2(new_n423), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n448), .A2(new_n451), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT17), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n448), .A2(new_n460), .A3(KEYINPUT17), .A4(new_n451), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n457), .A2(new_n465), .A3(KEYINPUT79), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n273), .A2(new_n256), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n467), .A2(new_n251), .B1(new_n247), .B2(new_n273), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n316), .B1(new_n434), .B2(new_n431), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT7), .B1(new_n411), .B2(G20), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n446), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n250), .B1(new_n471), .B2(KEYINPUT16), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n468), .B1(new_n472), .B2(new_n447), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT18), .B1(new_n473), .B2(new_n425), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n454), .A2(new_n453), .A3(new_n455), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(new_n463), .A4(new_n464), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT79), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n403), .A2(new_n466), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n480));
  INV_X1    g0280(.A(G107), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n260), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n482), .B2(new_n483), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n251), .B1(new_n242), .B2(G33), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G107), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  MUX2_X1   g0289(.A(G250), .B(G257), .S(G1698), .Z(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n418), .A3(new_n368), .ZN(new_n491));
  INV_X1    g0291(.A(G294), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n264), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n381), .B1(new_n493), .B2(KEYINPUT90), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT90), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n491), .B(new_n495), .C1(new_n264), .C2(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G190), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n290), .A2(G1), .ZN(new_n499));
  NAND2_X1  g0299(.A1(KEYINPUT5), .A2(G41), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(KEYINPUT5), .A2(G41), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT82), .B1(new_n503), .B2(new_n293), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n242), .A2(G45), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n289), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n505), .B1(new_n507), .B2(new_n500), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT82), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n379), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n508), .A2(new_n287), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G264), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n497), .A2(new_n498), .A3(new_n511), .A4(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n511), .ZN(new_n515));
  INV_X1    g0315(.A(new_n513), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(new_n494), .C2(new_n496), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n517), .B2(G200), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT23), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n212), .B2(G107), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n481), .A2(KEYINPUT23), .A3(G20), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n520), .A2(new_n521), .B1(new_n274), .B2(G116), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n418), .A2(new_n212), .A3(G87), .A4(new_n368), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT86), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT22), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n405), .A2(KEYINPUT22), .A3(G20), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT87), .B1(new_n527), .B2(new_n371), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT87), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n279), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n524), .B1(new_n523), .B2(KEYINPUT22), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n522), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT88), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT88), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n536), .B(new_n522), .C1(new_n532), .C2(new_n533), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n535), .A2(KEYINPUT24), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n534), .A2(KEYINPUT88), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n249), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n489), .B(new_n518), .C1(new_n538), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n247), .A2(G97), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n486), .B2(G97), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n481), .B1(new_n441), .B2(new_n442), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT6), .ZN(new_n546));
  INV_X1    g0346(.A(G97), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n546), .A2(new_n547), .A3(G107), .ZN(new_n548));
  XNOR2_X1  g0348(.A(G97), .B(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(new_n546), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n550), .A2(new_n212), .B1(new_n282), .B2(new_n265), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n249), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n504), .A2(new_n510), .B1(new_n512), .B2(G257), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n418), .A2(G244), .A3(new_n280), .A4(new_n368), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n368), .A2(new_n370), .A3(G250), .A4(G1698), .ZN(new_n559));
  AND2_X1   g0359(.A1(KEYINPUT4), .A2(G244), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n368), .A2(new_n370), .A3(new_n560), .A4(new_n280), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G283), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT80), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(KEYINPUT80), .A2(G33), .A3(G283), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n559), .A2(new_n561), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n381), .B1(new_n558), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n555), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n553), .B1(G190), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(KEYINPUT81), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT81), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n567), .B1(new_n557), .B2(new_n556), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(new_n381), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n555), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(G200), .B1(new_n576), .B2(KEYINPUT83), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n572), .A2(new_n575), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n578), .A2(KEYINPUT83), .A3(new_n554), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n571), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n311), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n554), .B1(new_n574), .B2(new_n381), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n552), .A2(new_n544), .B1(new_n582), .B2(new_n387), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n411), .A2(new_n212), .A3(G68), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT19), .B1(new_n274), .B2(G97), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n212), .B1(new_n343), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n405), .A2(new_n547), .A3(new_n481), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n249), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n260), .A2(new_n391), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(G87), .B2(new_n486), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n373), .A2(G1698), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n411), .A2(new_n596), .B1(G33), .B2(G116), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n411), .A2(KEYINPUT84), .A3(G244), .A4(G1698), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n418), .A2(G244), .A3(G1698), .A4(new_n368), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT84), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n287), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n505), .A2(G250), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n379), .A2(new_n499), .B1(new_n604), .B2(new_n381), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n595), .B(new_n607), .C1(new_n498), .C2(new_n606), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n542), .A2(new_n580), .A3(new_n584), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n242), .A2(G33), .ZN(new_n610));
  INV_X1    g0410(.A(new_n391), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n252), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n592), .A2(new_n593), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n605), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n602), .B2(new_n287), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n615), .B2(G169), .ZN(new_n616));
  AOI211_X1 g0416(.A(G179), .B(new_n614), .C1(new_n602), .C2(new_n287), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n503), .A2(G270), .A3(new_n381), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n511), .A2(new_n620), .ZN(new_n621));
  MUX2_X1   g0421(.A(G257), .B(G264), .S(G1698), .Z(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(new_n418), .A3(new_n368), .ZN(new_n623));
  XOR2_X1   g0423(.A(KEYINPUT85), .B(G303), .Z(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n371), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n381), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(G169), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n247), .A2(G116), .A3(new_n250), .A4(new_n610), .ZN(new_n628));
  INV_X1    g0428(.A(G116), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n260), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(G20), .B1(new_n264), .B2(G97), .ZN(new_n631));
  INV_X1    g0431(.A(new_n565), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT80), .B1(G33), .B2(G283), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n248), .A2(new_n211), .B1(G20), .B2(new_n629), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n634), .A2(KEYINPUT20), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT20), .B1(new_n634), .B2(new_n635), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n628), .B(new_n630), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n619), .B1(new_n627), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(G200), .B1(new_n621), .B2(new_n626), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n504), .A2(new_n510), .B1(new_n512), .B2(G270), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n623), .A2(new_n625), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n287), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(G190), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n621), .A2(new_n311), .A3(new_n626), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n638), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n387), .B1(new_n642), .B2(new_n644), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(KEYINPUT21), .A3(new_n638), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n640), .A2(new_n646), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n618), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n540), .A2(new_n249), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n535), .A2(KEYINPUT24), .A3(new_n537), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n488), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n516), .B1(new_n494), .B2(new_n496), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n511), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n387), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n517), .A2(new_n311), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n652), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n479), .A2(new_n609), .A3(new_n661), .ZN(G372));
  INV_X1    g0462(.A(new_n313), .ZN(new_n663));
  INV_X1    g0463(.A(new_n358), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n386), .A2(new_n387), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n393), .A2(new_n394), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n665), .A2(new_n666), .A3(new_n397), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n664), .B1(new_n365), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n465), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n457), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n303), .A2(new_n314), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n663), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n584), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n673), .B(new_n608), .C1(new_n617), .C2(new_n616), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT91), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n606), .A2(new_n677), .A3(new_n387), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT91), .B1(new_n615), .B2(G169), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n678), .B(KEYINPUT92), .C1(new_n679), .C2(new_n617), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n603), .A2(new_n311), .A3(new_n605), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n682), .B(KEYINPUT91), .C1(G169), .C2(new_n615), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT92), .B1(new_n683), .B2(new_n678), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n613), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n685), .A2(new_n673), .A3(new_n608), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n676), .B1(new_n686), .B2(new_n675), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n655), .A2(new_n660), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n640), .A2(new_n648), .A3(new_n650), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n685), .B1(new_n690), .B2(new_n609), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n672), .B1(new_n692), .B2(new_n479), .ZN(G369));
  INV_X1    g0493(.A(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n242), .A2(new_n212), .A3(G13), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT93), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT93), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n694), .A3(new_n697), .ZN(new_n700));
  AND4_X1   g0500(.A1(G213), .A2(new_n699), .A3(G343), .A4(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n542), .B1(new_n655), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n489), .B1(new_n538), .B2(new_n541), .ZN(new_n704));
  INV_X1    g0504(.A(new_n660), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n688), .A2(new_n702), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n689), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n701), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n708), .ZN(new_n713));
  INV_X1    g0513(.A(new_n709), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n702), .A2(new_n639), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n689), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n651), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n713), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n206), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n721), .A2(KEYINPUT94), .A3(G41), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT94), .B1(new_n721), .B2(G41), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n589), .A2(G116), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n725), .A2(new_n242), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n210), .B2(new_n725), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  NAND4_X1  g0530(.A1(new_n685), .A2(KEYINPUT26), .A3(new_n673), .A4(new_n608), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n674), .A2(new_n675), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND4_X1   g0533(.A1(new_n542), .A2(new_n580), .A3(new_n584), .A4(new_n608), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n706), .A2(new_n710), .ZN(new_n735));
  INV_X1    g0535(.A(new_n684), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n680), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n734), .A2(new_n735), .B1(new_n613), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT29), .A3(new_n702), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n692), .A2(new_n701), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(KEYINPUT29), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n578), .A2(new_n554), .ZN(new_n743));
  AOI21_X1  g0543(.A(G179), .B1(new_n642), .B2(new_n644), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n743), .A2(new_n657), .A3(new_n606), .A4(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n656), .A2(new_n570), .A3(new_n615), .A4(new_n647), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n642), .A2(G179), .A3(new_n644), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n582), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(KEYINPUT30), .A3(new_n656), .A4(new_n615), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n745), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT95), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n752), .A2(new_n701), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT31), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n754), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n609), .A2(new_n661), .A3(new_n701), .ZN(new_n762));
  OAI21_X1  g0562(.A(G330), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n742), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n730), .B1(new_n765), .B2(G1), .ZN(G364));
  INV_X1    g0566(.A(new_n718), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n212), .A2(G13), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n242), .B1(new_n769), .B2(G45), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n725), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n717), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n279), .A2(new_n206), .ZN(new_n775));
  INV_X1    g0575(.A(G355), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n776), .B1(G116), .B2(new_n206), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n411), .A2(new_n721), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n290), .B2(new_n210), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n240), .A2(G45), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n211), .B1(G20), .B2(new_n387), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n772), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n212), .A2(G179), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G190), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(G329), .ZN(new_n794));
  XOR2_X1   g0594(.A(KEYINPUT33), .B(G317), .Z(new_n795));
  NOR2_X1   g0595(.A1(new_n212), .A2(new_n311), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n278), .A2(G190), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n790), .A2(new_n797), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n795), .A2(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n796), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n802), .A2(new_n498), .A3(G200), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n794), .B(new_n801), .C1(G322), .C2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n498), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n212), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G294), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n498), .A2(new_n278), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n796), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n279), .B1(new_n811), .B2(G326), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n796), .A2(new_n791), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n809), .A2(new_n790), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G311), .A2(new_n814), .B1(new_n816), .B2(G303), .ZN(new_n817));
  AND4_X1   g0617(.A1(new_n804), .A2(new_n808), .A3(new_n812), .A4(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(KEYINPUT97), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(KEYINPUT97), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n810), .A2(new_n258), .B1(new_n813), .B2(new_n282), .ZN(new_n821));
  INV_X1    g0621(.A(new_n798), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n371), .B(new_n821), .C1(G68), .C2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n824));
  NAND3_X1  g0624(.A1(new_n793), .A2(G159), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n793), .B2(G159), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G97), .B2(new_n807), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n799), .A2(new_n481), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n815), .A2(new_n405), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n271), .C2(new_n803), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n823), .A2(new_n825), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n819), .A2(new_n820), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n789), .B1(new_n832), .B2(new_n786), .ZN(new_n833));
  INV_X1    g0633(.A(new_n785), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n717), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n774), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  NAND2_X1  g0637(.A1(new_n701), .A2(new_n666), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n401), .A2(new_n838), .B1(new_n397), .B2(new_n395), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n398), .A2(new_n701), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT98), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT98), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n400), .A2(new_n394), .A3(new_n393), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n396), .A2(new_n278), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n398), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n667), .A2(new_n702), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n741), .B(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n772), .B1(new_n850), .B2(new_n763), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n763), .B2(new_n850), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n813), .A2(new_n629), .B1(new_n799), .B2(new_n405), .ZN(new_n853));
  INV_X1    g0653(.A(new_n803), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n492), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(G303), .C2(new_n811), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n807), .A2(G97), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n279), .B1(new_n816), .B2(G107), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G283), .A2(new_n822), .B1(new_n793), .B2(G311), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n815), .A2(new_n258), .B1(new_n799), .B2(new_n316), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G132), .B2(new_n793), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n430), .B1(new_n807), .B2(new_n271), .ZN(new_n863));
  INV_X1    g0663(.A(G159), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n813), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(G137), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n810), .A2(new_n866), .B1(new_n798), .B2(new_n263), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n865), .B(new_n867), .C1(G143), .C2(new_n803), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n862), .B(new_n863), .C1(new_n868), .C2(KEYINPUT34), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(KEYINPUT34), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n786), .ZN(new_n872));
  INV_X1    g0672(.A(new_n772), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n786), .A2(new_n783), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n282), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n872), .B(new_n875), .C1(new_n849), .C2(new_n784), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n852), .A2(new_n876), .ZN(G384));
  INV_X1    g0677(.A(new_n550), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n878), .A2(KEYINPUT35), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(KEYINPUT35), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(G116), .A3(new_n213), .A4(new_n880), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT36), .Z(new_n882));
  NAND3_X1  g0682(.A1(new_n210), .A2(new_n426), .A3(G77), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n258), .A2(G68), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n242), .B(G13), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n479), .ZN(new_n887));
  INV_X1    g0687(.A(new_n661), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n734), .A2(new_n888), .A3(new_n702), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT31), .B1(new_n752), .B2(new_n701), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n753), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT102), .Z(new_n894));
  INV_X1    g0694(.A(KEYINPUT101), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n429), .B1(new_n433), .B2(new_n435), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n437), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n468), .B1(new_n472), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n461), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n898), .A2(new_n425), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT37), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n454), .A2(new_n455), .ZN(new_n903));
  INV_X1    g0703(.A(new_n899), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n454), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n903), .A2(new_n905), .A3(new_n906), .A4(new_n461), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n898), .A2(new_n899), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n476), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(new_n905), .A3(new_n461), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n907), .ZN(new_n914));
  INV_X1    g0714(.A(new_n905), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n476), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT38), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n895), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n339), .A2(new_n701), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n358), .A2(new_n365), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(new_n358), .B2(new_n365), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n849), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n889), .B2(new_n891), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n913), .A2(new_n907), .B1(new_n476), .B2(new_n915), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n924), .B(KEYINPUT101), .C1(KEYINPUT38), .C2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n918), .A2(new_n923), .A3(KEYINPUT40), .A4(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT40), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n908), .B2(new_n910), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n911), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT98), .B1(new_n839), .B2(new_n840), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n846), .A2(new_n847), .A3(new_n842), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n919), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n366), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n358), .A2(new_n365), .A3(new_n919), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n760), .A2(new_n755), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n937), .B1(new_n762), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n928), .B1(new_n930), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n927), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n894), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n894), .A2(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(G330), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n920), .A2(new_n921), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n702), .B(new_n849), .C1(new_n687), .C2(new_n691), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n945), .B1(new_n946), .B2(new_n847), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT38), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n902), .A2(new_n907), .ZN(new_n949));
  INV_X1    g0749(.A(new_n909), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n457), .B2(new_n465), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n948), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n924), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n899), .B1(new_n452), .B2(new_n456), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT39), .B1(new_n911), .B2(new_n929), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT39), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n924), .B(new_n957), .C1(KEYINPUT38), .C2(new_n925), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(KEYINPUT100), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n664), .A2(new_n702), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT99), .Z(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT100), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n953), .A2(new_n963), .A3(KEYINPUT39), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n959), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n954), .A2(new_n955), .A3(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n887), .B(new_n740), .C1(new_n741), .C2(KEYINPUT29), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n672), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n966), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n944), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n242), .B2(new_n769), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n944), .A2(new_n969), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n886), .B1(new_n971), .B2(new_n972), .ZN(G367));
  NAND2_X1  g0773(.A1(new_n553), .A2(new_n701), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n580), .A2(new_n584), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n673), .A2(new_n701), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n719), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT103), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n685), .A2(new_n595), .A3(new_n702), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n685), .B(new_n608), .C1(new_n595), .C2(new_n702), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n979), .B(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n712), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n977), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n688), .A2(new_n580), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n701), .B1(new_n988), .B2(new_n584), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n986), .B2(KEYINPUT42), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n987), .A2(new_n990), .B1(KEYINPUT43), .B2(new_n982), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n984), .A2(new_n991), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n724), .B(KEYINPUT41), .ZN(new_n994));
  INV_X1    g0794(.A(new_n977), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n713), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT44), .Z(new_n997));
  NOR2_X1   g0797(.A1(new_n713), .A2(new_n995), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n719), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n709), .A2(new_n711), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT104), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1002), .A2(new_n1003), .A3(new_n767), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n767), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1005), .A2(new_n985), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n985), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n764), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n997), .B(new_n999), .C1(new_n718), .C2(new_n714), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1001), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n994), .B1(new_n1012), .B2(new_n765), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n992), .B(new_n993), .C1(new_n1013), .C2(new_n771), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n787), .B1(new_n206), .B2(new_n391), .C1(new_n779), .C2(new_n231), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n873), .B1(new_n1015), .B2(KEYINPUT105), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(KEYINPUT105), .B2(new_n1015), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n854), .A2(new_n263), .B1(new_n792), .B2(new_n866), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n799), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n371), .B(new_n1018), .C1(G77), .C2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G143), .A2(new_n811), .B1(new_n816), .B2(new_n271), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G50), .A2(new_n814), .B1(new_n822), .B2(G159), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n806), .A2(new_n316), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n799), .A2(new_n547), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G283), .B2(new_n814), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n430), .C1(new_n481), .C2(new_n806), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n816), .A2(G116), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT46), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G294), .A2(new_n822), .B1(new_n793), .B2(G317), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n803), .A2(new_n624), .B1(new_n811), .B2(G311), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1025), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT47), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1017), .B1(new_n1035), .B2(new_n786), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n982), .B2(new_n834), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1014), .A2(new_n1037), .ZN(G387));
  INV_X1    g0838(.A(new_n1010), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1009), .A2(new_n764), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n725), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n792), .A2(new_n263), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n316), .A2(new_n813), .B1(new_n815), .B2(new_n282), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G50), .C2(new_n803), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n806), .A2(new_n391), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n430), .B(new_n1026), .C1(G159), .C2(new_n811), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n273), .A2(new_n822), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G116), .A2(new_n1019), .B1(new_n793), .B2(G326), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n806), .A2(new_n800), .B1(new_n815), .B2(new_n492), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n803), .A2(G317), .B1(new_n624), .B2(new_n814), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G322), .A2(new_n811), .B1(new_n822), .B2(G311), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n430), .B(new_n1050), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n786), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n775), .A2(new_n726), .B1(G107), .B2(new_n206), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n228), .A2(new_n290), .ZN(new_n1064));
  AOI211_X1 g0864(.A(G45), .B(new_n727), .C1(G68), .C2(G77), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n389), .A2(G50), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT50), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n779), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1063), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1062), .B(new_n772), .C1(new_n788), .C2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n714), .B2(new_n785), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1009), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n771), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1041), .A2(new_n1073), .ZN(G393));
  AND2_X1   g0874(.A1(new_n1012), .A2(new_n725), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1001), .A2(new_n1011), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1076), .A2(KEYINPUT108), .A3(new_n1010), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT108), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1001), .A2(new_n1011), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n1039), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1075), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n995), .A2(new_n785), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT106), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n803), .A2(G311), .B1(new_n811), .B2(G317), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT52), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G294), .A2(new_n814), .B1(new_n822), .B2(new_n624), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n629), .B2(new_n806), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G283), .A2(new_n816), .B1(new_n793), .B2(G322), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(new_n371), .C1(new_n481), .C2(new_n799), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT107), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n803), .A2(G159), .B1(new_n811), .B2(G150), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  AOI22_X1  g0893(.A1(G50), .A2(new_n822), .B1(new_n793), .B2(G143), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n389), .B2(new_n813), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n806), .A2(new_n282), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n411), .B1(new_n316), .B2(new_n815), .C1(new_n405), .C2(new_n799), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1088), .A2(new_n1091), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n786), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n235), .A2(new_n778), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n788), .B1(G97), .B2(new_n721), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n873), .B(new_n1101), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1076), .A2(new_n771), .B1(new_n1083), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1081), .A2(new_n1105), .ZN(G390));
  INV_X1    g0906(.A(new_n874), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n811), .A2(G283), .B1(new_n793), .B2(G294), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1108), .B1(new_n316), .B2(new_n799), .C1(new_n629), .C2(new_n854), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1109), .A2(new_n279), .A3(new_n829), .A4(new_n1096), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n547), .A2(new_n813), .B1(new_n798), .B2(new_n481), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT114), .Z(new_n1112));
  NAND2_X1  g0912(.A1(new_n811), .A2(G128), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT54), .B(G143), .ZN(new_n1114));
  INV_X1    g0914(.A(G132), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1113), .B1(new_n813), .B2(new_n1114), .C1(new_n854), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n816), .A2(G150), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G137), .A2(new_n822), .B1(new_n793), .B2(G125), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n864), .B2(new_n806), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n279), .B1(new_n799), .B2(new_n258), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT113), .Z(new_n1123));
  AOI22_X1  g0923(.A1(new_n1110), .A2(new_n1112), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n772), .B1(new_n273), .B2(new_n1107), .C1(new_n1124), .C2(new_n1100), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n959), .A2(new_n964), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n783), .ZN(new_n1127));
  INV_X1    g0927(.A(G330), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n889), .B2(new_n891), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n937), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1126), .B1(new_n947), .B2(new_n962), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n945), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n701), .B(new_n933), .C1(new_n733), .C2(new_n738), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n840), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n918), .A2(new_n961), .A3(new_n926), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1130), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT109), .ZN(new_n1139));
  AOI211_X1 g0939(.A(KEYINPUT100), .B(new_n957), .C1(new_n952), .C2(new_n924), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n963), .B1(new_n953), .B2(KEYINPUT39), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n958), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n946), .A2(new_n847), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1132), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n1144), .B2(new_n961), .ZN(new_n1145));
  OR3_X1    g0945(.A1(new_n763), .A2(new_n933), .A3(new_n945), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n739), .A2(new_n702), .A3(new_n849), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n945), .B1(new_n1147), .B2(new_n847), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1148), .B2(new_n1135), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1139), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n763), .A2(new_n933), .A3(new_n945), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(KEYINPUT109), .A3(new_n1131), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1138), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1127), .B1(new_n1154), .B2(new_n771), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1147), .A2(new_n847), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1129), .A2(KEYINPUT111), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n849), .B1(new_n1129), .B2(KEYINPUT111), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n945), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n945), .B1(new_n763), .B2(new_n933), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1130), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1157), .A2(new_n1160), .B1(new_n1162), .B2(new_n1143), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n887), .A2(KEYINPUT110), .A3(new_n1129), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT110), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n892), .A2(G330), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n479), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n967), .A2(new_n672), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT112), .B1(new_n1163), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1138), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT109), .B1(new_n1152), .B2(new_n1131), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1152), .A2(KEYINPUT109), .A3(new_n1131), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1170), .B(new_n1171), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n725), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1154), .A2(new_n1170), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1155), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT115), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(KEYINPUT115), .B(new_n1155), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(G378));
  NAND3_X1  g0982(.A1(new_n927), .A2(new_n940), .A3(G330), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n308), .A2(new_n899), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n315), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n315), .A2(new_n1184), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1183), .A2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1192), .A2(G330), .A3(new_n927), .A4(new_n940), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(new_n966), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n965), .A2(new_n955), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n954), .A2(new_n1198), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT57), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1162), .A2(new_n1143), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1171), .B(new_n1203), .C1(new_n1173), .C2(new_n1172), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1169), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1200), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(KEYINPUT117), .B1(new_n1206), .B2(new_n724), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT117), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1169), .B1(new_n1154), .B2(new_n1203), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n725), .C1(new_n1209), .C2(new_n1200), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1199), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT116), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1198), .A2(new_n1194), .A3(new_n954), .A4(new_n1195), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1199), .A2(KEYINPUT116), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1211), .B1(new_n1209), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1207), .A2(new_n1210), .A3(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n411), .A2(G41), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G50), .B(new_n1220), .C1(new_n264), .C2(new_n289), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G116), .A2(new_n811), .B1(new_n822), .B2(G97), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n1220), .C1(new_n391), .C2(new_n813), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n271), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n854), .A2(new_n481), .B1(new_n1224), .B2(new_n799), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n815), .A2(new_n282), .B1(new_n792), .B2(new_n800), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1223), .A2(new_n1225), .A3(new_n1023), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1221), .B1(new_n1227), .B2(KEYINPUT58), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n822), .A2(G132), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n815), .B2(new_n1114), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n803), .A2(G128), .B1(new_n811), .B2(G125), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n866), .B2(new_n813), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(G150), .C2(new_n807), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n264), .B(new_n289), .C1(new_n799), .C2(new_n864), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G124), .B2(new_n793), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT59), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1237), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1228), .B1(KEYINPUT58), .B2(new_n1227), .C1(new_n1235), .C2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n786), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1241), .B(new_n772), .C1(G50), .C2(new_n1107), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1193), .B2(new_n783), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n771), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1219), .A2(new_n1245), .ZN(G375));
  OAI21_X1  g1046(.A(new_n772), .B1(G68), .B2(new_n1107), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1132), .A2(new_n784), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n279), .B(new_n1045), .C1(G77), .C2(new_n1019), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n481), .A2(new_n813), .B1(new_n798), .B2(new_n629), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT118), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n803), .A2(G283), .B1(new_n811), .B2(G294), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G97), .A2(new_n816), .B1(new_n793), .B2(G303), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n815), .A2(new_n864), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n854), .A2(new_n866), .B1(new_n1224), .B2(new_n799), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(G128), .C2(new_n793), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1257), .B(new_n411), .C1(new_n258), .C2(new_n806), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n814), .A2(G150), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1259), .B1(new_n1115), .B2(new_n810), .C1(new_n798), .C2(new_n1114), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1254), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1247), .B(new_n1248), .C1(new_n786), .C2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1203), .B2(new_n771), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT119), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n994), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1163), .A2(new_n1169), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(G381));
  INV_X1    g1069(.A(KEYINPUT121), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1177), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT121), .B(new_n1155), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(G375), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(G390), .A2(G387), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1041), .A2(new_n836), .A3(new_n1073), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G384), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1277), .A2(KEYINPUT120), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G381), .B1(new_n1277), .B2(KEYINPUT120), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1274), .A2(new_n1275), .A3(new_n1278), .A4(new_n1279), .ZN(G407));
  INV_X1    g1080(.A(G213), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(G343), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1274), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G407), .A2(G213), .A3(new_n1283), .ZN(G409));
  INV_X1    g1084(.A(KEYINPUT125), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1276), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n836), .B1(new_n1041), .B2(new_n1073), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1081), .A2(new_n1105), .B1(new_n1014), .B2(new_n1037), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1285), .B(new_n1288), .C1(new_n1275), .C2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G390), .A2(G387), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1081), .A2(new_n1014), .A3(new_n1037), .A4(new_n1105), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1288), .A2(new_n1285), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT125), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1219), .A2(new_n1179), .A3(new_n1180), .A4(new_n1245), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1244), .A2(new_n1266), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1243), .B1(new_n1300), .B2(new_n771), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1271), .A2(new_n1302), .A3(new_n1272), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1282), .B1(new_n1297), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1265), .A2(KEYINPUT60), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1267), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(KEYINPUT122), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT122), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1305), .A2(new_n1308), .A3(new_n1267), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1163), .A2(KEYINPUT60), .A3(new_n1169), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1307), .A2(new_n725), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT123), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n852), .A2(new_n1312), .A3(new_n876), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1311), .A2(new_n1264), .A3(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(G384), .B(new_n1312), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1311), .B2(new_n1264), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT62), .B1(new_n1304), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT126), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1297), .A2(new_n1303), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1282), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1319), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  AOI211_X1 g1122(.A(KEYINPUT126), .B(new_n1282), .C1(new_n1297), .C2(new_n1303), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1318), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(G2897), .B(new_n1282), .C1(new_n1314), .C2(new_n1316), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1311), .A2(new_n1264), .A3(new_n1313), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1282), .A2(G2897), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1311), .A2(new_n1264), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1328), .B(new_n1329), .C1(new_n1330), .C2(new_n1315), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1327), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1333), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT61), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1296), .B1(new_n1326), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT124), .ZN(new_n1338));
  OR3_X1    g1138(.A1(new_n1332), .A2(new_n1338), .A3(new_n1304), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1338), .B1(new_n1332), .B2(new_n1304), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1324), .A2(KEYINPUT63), .A3(new_n1317), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT63), .B1(new_n1304), .B2(new_n1317), .ZN(new_n1343));
  NOR3_X1   g1143(.A1(new_n1296), .A2(new_n1343), .A3(KEYINPUT61), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1341), .A2(new_n1342), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1337), .A2(new_n1345), .ZN(G405));
  MUX2_X1   g1146(.A(new_n1181), .B(new_n1273), .S(G375), .Z(new_n1347));
  OR2_X1    g1147(.A1(new_n1296), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1296), .A2(new_n1347), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1317), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1351), .A2(KEYINPUT127), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1350), .A2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1348), .A2(new_n1352), .A3(new_n1349), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(G402));
endmodule


