//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT78), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(KEYINPUT78), .A3(G125), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n188), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n187), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n197), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n189), .A2(KEYINPUT78), .A3(G125), .ZN(new_n200));
  XNOR2_X1  g014(.A(G125), .B(G140), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(new_n193), .ZN(new_n202));
  OAI211_X1 g016(.A(G146), .B(new_n199), .C1(new_n202), .C2(new_n188), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n206), .B(KEYINPUT23), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n204), .B1(G110), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n209), .B(KEYINPUT77), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  XOR2_X1   g027(.A(KEYINPUT24), .B(G110), .Z(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n213), .A2(new_n214), .B1(new_n210), .B2(G110), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n201), .A2(new_n187), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n203), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n196), .A2(new_n197), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT79), .A3(G146), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n217), .A2(new_n218), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT70), .B(G953), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(G221), .A3(G234), .ZN(new_n226));
  XOR2_X1   g040(.A(new_n226), .B(KEYINPUT22), .Z(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n216), .A2(new_n223), .A3(new_n229), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(G234), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G902), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(KEYINPUT81), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n233), .A2(new_n236), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n231), .A2(new_n236), .A3(new_n232), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n242), .A3(new_n243), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n241), .B1(new_n249), .B2(new_n237), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(G116), .B(G119), .Z(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT2), .B(G113), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  OAI21_X1  g071(.A(G128), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT65), .A2(G143), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT65), .A2(G143), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n259), .A2(new_n260), .A3(G146), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT66), .B1(new_n187), .B2(G143), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n255), .A3(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n258), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT65), .B(G143), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n256), .B1(new_n268), .B2(G146), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n257), .A3(G128), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n262), .B(new_n264), .C1(new_n268), .C2(G146), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n258), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n267), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT67), .B(G137), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT11), .A3(G134), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT11), .B1(new_n228), .B2(G134), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n228), .A2(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n276), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  OR2_X1    g095(.A1(KEYINPUT67), .A2(G137), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT67), .A2(G137), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n277), .B1(new_n285), .B2(new_n279), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n274), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(KEYINPUT0), .A2(G128), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n289), .B(KEYINPUT64), .Z(new_n290));
  OAI211_X1 g104(.A(new_n271), .B(new_n290), .C1(KEYINPUT0), .C2(G128), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n269), .A2(KEYINPUT0), .A3(G128), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n277), .B1(new_n276), .B2(new_n280), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n291), .B(new_n292), .C1(new_n281), .C2(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n288), .A2(KEYINPUT30), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n274), .A2(KEYINPUT69), .A3(new_n287), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT69), .B1(new_n274), .B2(new_n287), .ZN(new_n298));
  INV_X1    g112(.A(new_n294), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n254), .B(new_n296), .C1(new_n300), .C2(KEYINPUT30), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n288), .A2(new_n294), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(new_n254), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G237), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n225), .A2(G210), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT74), .B1(new_n305), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n314));
  AOI211_X1 g128(.A(new_n314), .B(new_n311), .C1(new_n301), .C2(new_n304), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n254), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT73), .B1(new_n300), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT69), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n288), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n274), .A2(new_n287), .A3(KEYINPUT69), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n294), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(new_n254), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n318), .A2(new_n304), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT28), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n303), .A2(KEYINPUT28), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n311), .B(KEYINPUT72), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n316), .A2(new_n331), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n295), .B1(new_n322), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n303), .B1(new_n336), .B2(new_n254), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n314), .B1(new_n337), .B2(new_n311), .ZN(new_n338));
  AOI211_X1 g152(.A(new_n317), .B(new_n295), .C1(new_n322), .C2(new_n335), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT74), .B(new_n312), .C1(new_n339), .C2(new_n303), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n333), .A3(new_n340), .ZN(new_n341));
  AOI211_X1 g155(.A(new_n327), .B(new_n329), .C1(new_n325), .C2(KEYINPUT28), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT75), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n312), .A2(new_n333), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n303), .A2(KEYINPUT76), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n302), .A2(new_n254), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n328), .B(new_n344), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n349), .A2(new_n236), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n334), .A2(new_n343), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G472), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n326), .A2(new_n328), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n301), .A2(new_n304), .A3(new_n311), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT31), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n337), .A2(KEYINPUT31), .A3(new_n311), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n353), .A2(new_n329), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(G472), .A2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT32), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n322), .A2(new_n254), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n303), .B1(new_n362), .B2(KEYINPUT73), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n348), .B1(new_n363), .B2(new_n324), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n329), .B1(new_n364), .B2(new_n327), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n356), .A2(new_n357), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(new_n359), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n251), .B1(new_n352), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n225), .A2(G227), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G140), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n281), .A2(new_n293), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G104), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G101), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(G101), .ZN(new_n386));
  INV_X1    g200(.A(G101), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n378), .A2(new_n381), .A3(new_n387), .A4(new_n382), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n291), .A2(new_n292), .A3(new_n385), .A4(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n382), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n377), .A2(G107), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n388), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n274), .A2(KEYINPUT10), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT85), .B1(new_n261), .B2(new_n257), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n398), .B(KEYINPUT1), .C1(new_n268), .C2(G146), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(G128), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n256), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n259), .A2(new_n260), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(new_n187), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n394), .B1(new_n404), .B2(new_n270), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n390), .B(new_n396), .C1(new_n405), .C2(KEYINPUT10), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT10), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n403), .A2(KEYINPUT1), .A3(new_n205), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n400), .B2(new_n403), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n411), .B2(new_n394), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n412), .A2(KEYINPUT87), .A3(new_n390), .A4(new_n396), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n376), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n412), .A2(new_n376), .A3(new_n390), .A4(new_n396), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n375), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n274), .A2(new_n395), .ZN(new_n418));
  OAI22_X1  g232(.A1(new_n405), .A2(new_n418), .B1(new_n293), .B2(new_n281), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT12), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n415), .A3(new_n374), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G469), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n236), .ZN(new_n425));
  NAND2_X1  g239(.A1(G469), .A2(G902), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n374), .B(KEYINPUT84), .Z(new_n427));
  XNOR2_X1  g241(.A(new_n419), .B(KEYINPUT12), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n428), .B2(new_n416), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n415), .A2(new_n374), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n429), .B(G469), .C1(new_n432), .C2(new_n414), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n425), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n254), .A2(new_n389), .A3(new_n385), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n252), .A2(new_n253), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT5), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n208), .A3(G116), .ZN(new_n442));
  OAI211_X1 g256(.A(G113), .B(new_n442), .C1(new_n252), .C2(new_n441), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n395), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n439), .A2(KEYINPUT88), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT88), .B1(new_n439), .B2(new_n444), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n438), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT89), .A2(KEYINPUT6), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n439), .A2(new_n444), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n451));
  INV_X1    g265(.A(new_n448), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n438), .B(new_n452), .C1(new_n445), .C2(new_n446), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n291), .A2(new_n292), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G125), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(G125), .B2(new_n274), .ZN(new_n457));
  INV_X1    g271(.A(G224), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G953), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT90), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n457), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT7), .B1(new_n458), .B2(G953), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n450), .A2(new_n437), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n443), .A2(new_n440), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n394), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n444), .A3(KEYINPUT91), .ZN(new_n468));
  OR3_X1    g282(.A1(new_n466), .A2(KEYINPUT91), .A3(new_n394), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n437), .B(KEYINPUT8), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n463), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n456), .B(new_n472), .C1(G125), .C2(new_n274), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n464), .A2(new_n465), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n474), .A2(new_n236), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n462), .A2(new_n477), .A3(new_n475), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n436), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT9), .B(G234), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT82), .ZN(new_n483));
  OAI21_X1  g297(.A(G221), .B1(new_n483), .B2(G902), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT83), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n434), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G475), .ZN(new_n488));
  AND2_X1   g302(.A1(KEYINPUT70), .A2(G953), .ZN(new_n489));
  NOR2_X1   g303(.A1(KEYINPUT70), .A2(G953), .ZN(new_n490));
  OAI211_X1 g304(.A(G214), .B(new_n306), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n402), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n225), .A2(new_n255), .A3(G214), .A4(new_n306), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n277), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n493), .A3(G131), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n497), .A2(new_n496), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n204), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n494), .B1(new_n501), .B2(new_n277), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT18), .A4(G131), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT92), .B1(new_n504), .B2(new_n218), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n504), .A2(KEYINPUT92), .A3(new_n218), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n502), .B(new_n503), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G113), .B(G122), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n377), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT93), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n500), .A2(new_n510), .A3(new_n507), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(KEYINPUT93), .A3(new_n511), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n488), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n500), .A2(new_n510), .A3(new_n507), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n495), .A2(new_n497), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT19), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n201), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n202), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n187), .B(new_n520), .C1(new_n521), .C2(new_n519), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n518), .A2(new_n222), .A3(new_n220), .A4(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n510), .B1(new_n523), .B2(new_n507), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n488), .B(new_n236), .C1(new_n517), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT20), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n507), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n511), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n513), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT20), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n488), .A4(new_n236), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n516), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n533));
  INV_X1    g347(.A(G478), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n483), .A2(new_n235), .A3(G953), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n268), .A2(G128), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n205), .A2(G143), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n539), .A2(new_n283), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n542));
  INV_X1    g356(.A(G122), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(G116), .ZN(new_n544));
  INV_X1    g358(.A(G116), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT94), .A3(G122), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(G116), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G107), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n544), .A2(new_n546), .B1(G116), .B2(new_n543), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n380), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n539), .A2(KEYINPUT96), .A3(new_n554), .ZN(new_n555));
  OR2_X1    g369(.A1(KEYINPUT65), .A2(G143), .ZN(new_n556));
  NAND2_X1  g370(.A1(KEYINPUT65), .A2(G143), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n205), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n558), .A2(new_n553), .B1(new_n205), .B2(G143), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n558), .B2(new_n553), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n555), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI221_X4 g376(.A(new_n541), .B1(new_n550), .B2(new_n552), .C1(new_n562), .C2(G134), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n380), .B1(new_n548), .B2(KEYINPUT14), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n551), .B(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n283), .B1(new_n539), .B2(new_n540), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n541), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n538), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n541), .B1(new_n562), .B2(G134), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n550), .A2(new_n552), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n567), .A3(new_n537), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n536), .B1(new_n574), .B2(new_n236), .ZN(new_n575));
  AOI211_X1 g389(.A(G902), .B(new_n535), .C1(new_n569), .C2(new_n573), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n533), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n563), .A2(new_n568), .A3(new_n538), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n537), .B1(new_n572), .B2(new_n567), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n236), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n535), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n574), .A2(new_n236), .A3(new_n536), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(KEYINPUT97), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G952), .ZN(new_n585));
  AOI211_X1 g399(.A(G953), .B(new_n585), .C1(G234), .C2(G237), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n236), .B(new_n225), .C1(G234), .C2(G237), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT21), .B(G898), .Z(new_n590));
  OAI21_X1  g404(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT98), .Z(new_n592));
  NAND3_X1  g406(.A1(new_n532), .A2(new_n584), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n487), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n371), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  NOR2_X1   g410(.A1(new_n358), .A2(new_n360), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n365), .B2(new_n366), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n597), .B1(G472), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n251), .A2(new_n485), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n600), .A2(new_n434), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n481), .A2(new_n592), .ZN(new_n603));
  INV_X1    g417(.A(new_n532), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n605));
  OR3_X1    g419(.A1(new_n574), .A2(new_n605), .A3(KEYINPUT33), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n605), .A2(KEYINPUT33), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(KEYINPUT33), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n574), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(G478), .A3(new_n236), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n580), .A2(new_n534), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT100), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n604), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n603), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n602), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n525), .B2(KEYINPUT20), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n526), .A2(new_n531), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(new_n620), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n584), .ZN(new_n624));
  INV_X1    g438(.A(new_n516), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(new_n481), .A3(new_n625), .A4(new_n592), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n602), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G107), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n628), .B(new_n630), .ZN(G9));
  XOR2_X1   g445(.A(new_n224), .B(KEYINPUT103), .Z(new_n632));
  OR2_X1    g446(.A1(new_n230), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n635), .A2(new_n239), .B1(new_n249), .B2(new_n237), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n594), .A2(new_n637), .A3(new_n600), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  AOI21_X1  g456(.A(new_n636), .B1(new_n352), .B2(new_n370), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n587), .B1(new_n589), .B2(G900), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR4_X1   g459(.A1(new_n623), .A2(new_n584), .A3(new_n516), .A4(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n646), .A2(new_n481), .A3(new_n434), .A4(new_n486), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT106), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n643), .A2(new_n651), .A3(new_n648), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  NOR2_X1   g468(.A1(new_n347), .A2(new_n330), .ZN(new_n655));
  INV_X1    g469(.A(new_n354), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n236), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G472), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n370), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT108), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n370), .A2(new_n661), .A3(new_n658), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n479), .A2(new_n480), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(KEYINPUT107), .Z(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(KEYINPUT38), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(KEYINPUT38), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n584), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n604), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n664), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n434), .A2(new_n486), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n644), .B(KEYINPUT39), .Z(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n636), .B1(new_n677), .B2(KEYINPUT40), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n436), .B(new_n678), .C1(KEYINPUT40), .C2(new_n677), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n402), .ZN(G45));
  INV_X1    g495(.A(new_n487), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n615), .A2(new_n645), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n643), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  NAND2_X1  g499(.A1(new_n423), .A2(new_n236), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G469), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n687), .A2(new_n486), .A3(new_n425), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n371), .A2(new_n616), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  AOI22_X1  g505(.A1(new_n351), .A2(G472), .B1(new_n361), .B2(new_n369), .ZN(new_n692));
  INV_X1    g506(.A(new_n688), .ZN(new_n693));
  NOR4_X1   g507(.A1(new_n692), .A2(new_n693), .A3(new_n251), .A4(new_n626), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n545), .ZN(G18));
  INV_X1    g509(.A(new_n593), .ZN(new_n696));
  INV_X1    g510(.A(new_n481), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n643), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n328), .B1(new_n347), .B2(new_n348), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n329), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n360), .B1(new_n703), .B2(new_n366), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n705));
  INV_X1    g519(.A(G472), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n705), .B1(new_n598), .B2(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(KEYINPUT109), .B(G472), .C1(new_n358), .C2(G902), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n250), .A3(new_n688), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n603), .A2(new_n671), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n701), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  AOI211_X1 g527(.A(new_n704), .B(new_n251), .C1(new_n707), .C2(new_n708), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(KEYINPUT110), .A3(new_n688), .A4(new_n711), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  NAND4_X1  g531(.A1(new_n698), .A2(new_n637), .A3(new_n683), .A4(new_n709), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  XNOR2_X1  g533(.A(new_n426), .B(KEYINPUT111), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n425), .A2(new_n433), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(KEYINPUT112), .A3(new_n486), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT112), .B1(new_n721), .B2(new_n486), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n665), .A2(new_n436), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n371), .A2(new_n727), .A3(new_n683), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n371), .A2(new_n727), .A3(KEYINPUT42), .A4(new_n683), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  NAND3_X1  g547(.A1(new_n371), .A2(new_n727), .A3(new_n646), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT113), .B(G134), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G36));
  AND2_X1   g550(.A1(new_n614), .A2(KEYINPUT114), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n532), .B1(new_n614), .B2(KEYINPUT114), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT43), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n532), .B(KEYINPUT115), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n614), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n739), .B1(KEYINPUT43), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n600), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n637), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n726), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n429), .B1(new_n432), .B2(new_n414), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n429), .B(KEYINPUT45), .C1(new_n432), .C2(new_n414), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(G469), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT46), .B1(new_n751), .B2(new_n720), .ZN(new_n752));
  INV_X1    g566(.A(new_n425), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n720), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n485), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n676), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n746), .B(new_n758), .C1(new_n745), .C2(new_n744), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  NAND4_X1  g574(.A1(new_n692), .A2(new_n251), .A3(new_n683), .A4(new_n725), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT116), .Z(new_n762));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n754), .A2(new_n755), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(new_n485), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n756), .A2(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n189), .ZN(G42));
  AOI21_X1  g583(.A(new_n694), .B1(new_n713), .B2(new_n715), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n689), .A2(new_n699), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n732), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n575), .A2(new_n576), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n625), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n623), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n725), .A2(new_n775), .A3(KEYINPUT117), .A4(new_n644), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n674), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n352), .A2(new_n370), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n726), .A2(new_n623), .A3(new_n645), .A4(new_n774), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n777), .B(new_n778), .C1(KEYINPUT117), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n727), .A2(new_n683), .A3(new_n709), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n637), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n532), .B1(new_n575), .B2(new_n576), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n615), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n603), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n434), .A3(new_n601), .A4(new_n600), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n595), .A2(new_n788), .A3(new_n638), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n734), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n772), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n651), .B1(new_n643), .B2(new_n648), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n692), .A2(KEYINPUT106), .A3(new_n636), .A4(new_n647), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n684), .B(new_n718), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n481), .A2(new_n604), .A3(new_n670), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n486), .A2(new_n636), .A3(new_n644), .A4(new_n721), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n663), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n793), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n684), .A2(new_n718), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n653), .A2(new_n803), .A3(new_n800), .A4(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT53), .B1(new_n792), .B2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n802), .A2(KEYINPUT118), .A3(new_n804), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT118), .B1(new_n802), .B2(new_n804), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n772), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n783), .A2(KEYINPUT119), .A3(new_n790), .A4(new_n734), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n636), .B1(new_n780), .B2(new_n781), .ZN(new_n813));
  INV_X1    g627(.A(new_n734), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n789), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT53), .B1(new_n815), .B2(KEYINPUT119), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n806), .B1(new_n809), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT121), .B1(new_n585), .B2(G953), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n687), .A2(new_n425), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n485), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n765), .A2(new_n766), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n742), .A2(new_n586), .A3(new_n714), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n725), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT120), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n693), .A2(new_n587), .A3(new_n726), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n742), .A2(new_n637), .A3(new_n709), .A4(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n664), .A2(new_n250), .A3(new_n831), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n604), .A2(new_n614), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n827), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n825), .A2(new_n693), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n436), .B1(new_n667), .B2(new_n668), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT50), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n825), .A2(new_n838), .A3(new_n841), .A4(new_n693), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n830), .A2(new_n836), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n827), .A2(new_n835), .A3(new_n832), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n829), .B(new_n828), .C1(new_n846), .C2(new_n843), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n742), .A2(new_n371), .A3(new_n831), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT48), .Z(new_n849));
  INV_X1    g663(.A(new_n615), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n833), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n821), .A2(new_n845), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n805), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n802), .A2(KEYINPUT118), .A3(new_n804), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n792), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n805), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n810), .A2(new_n815), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT53), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n857), .A2(new_n860), .A3(KEYINPUT54), .ZN(new_n861));
  OR2_X1    g675(.A1(KEYINPUT121), .A2(G953), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n820), .A2(new_n852), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n825), .A2(new_n697), .A3(new_n693), .ZN(new_n864));
  OAI22_X1  g678(.A1(new_n863), .A2(new_n864), .B1(G952), .B2(G953), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n822), .B(KEYINPUT49), .Z(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(new_n436), .A3(new_n741), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n664), .A3(new_n601), .A4(new_n669), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(G75));
  INV_X1    g683(.A(new_n225), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n585), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT125), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n855), .B1(new_n791), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n772), .B1(KEYINPUT119), .B2(new_n815), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n854), .A2(new_n856), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n236), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT56), .B1(new_n878), .B2(G210), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n454), .B(new_n461), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT122), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n872), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n818), .B2(new_n236), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n876), .A2(new_n877), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(KEYINPUT123), .A3(G902), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n478), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n882), .A2(KEYINPUT124), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(KEYINPUT124), .B2(new_n882), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n883), .B1(new_n888), .B2(new_n891), .ZN(G51));
  INV_X1    g706(.A(new_n872), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n720), .A2(KEYINPUT57), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n720), .A2(KEYINPUT57), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n876), .A2(new_n877), .A3(new_n819), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n819), .B1(new_n876), .B2(new_n877), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n894), .B(new_n895), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n423), .ZN(new_n899));
  INV_X1    g713(.A(new_n751), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n885), .A2(new_n900), .A3(new_n887), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n893), .B1(new_n899), .B2(new_n901), .ZN(G54));
  AND2_X1   g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n885), .A2(new_n887), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n529), .ZN(new_n905));
  INV_X1    g719(.A(new_n529), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n885), .A2(new_n906), .A3(new_n887), .A4(new_n903), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n893), .B1(new_n905), .B2(new_n907), .ZN(G60));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT59), .Z(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n820), .B2(new_n861), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n872), .B1(new_n911), .B2(new_n610), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n610), .B1(new_n896), .B2(new_n897), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n910), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT60), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n886), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n234), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n886), .A2(new_n635), .A3(new_n917), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n872), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n919), .A2(KEYINPUT61), .A3(new_n872), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G66));
  NAND3_X1  g739(.A1(new_n770), .A2(new_n790), .A3(new_n771), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n590), .A2(G224), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n926), .A2(new_n225), .B1(G953), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n454), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(G898), .B2(new_n225), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT126), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n928), .B(new_n931), .ZN(G69));
  OAI21_X1  g746(.A(new_n520), .B1(new_n521), .B2(new_n519), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n336), .B(new_n933), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(G227), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n870), .A2(G900), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n796), .B1(new_n672), .B2(new_n679), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT62), .ZN(new_n939));
  INV_X1    g753(.A(new_n768), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n371), .ZN(new_n942));
  NOR4_X1   g756(.A1(new_n942), .A2(new_n677), .A3(new_n726), .A4(new_n786), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT127), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(new_n759), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n225), .ZN(new_n946));
  OAI221_X1 g760(.A(new_n935), .B1(new_n936), .B2(new_n937), .C1(new_n941), .C2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n940), .A2(new_n732), .A3(new_n734), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n758), .A2(new_n371), .A3(new_n798), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n759), .A2(new_n653), .A3(new_n803), .A4(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n225), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n951), .B(new_n934), .C1(G227), .C2(new_n937), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n947), .A2(new_n952), .ZN(G72));
  NAND2_X1  g767(.A1(G472), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT63), .Z(new_n955));
  INV_X1    g769(.A(new_n926), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n945), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n941), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n337), .A2(new_n312), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n893), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n948), .A2(new_n926), .A3(new_n950), .ZN(new_n961));
  INV_X1    g775(.A(new_n955), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n312), .B(new_n337), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n316), .A2(new_n354), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n857), .A2(new_n860), .A3(new_n955), .A4(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n960), .A2(new_n963), .A3(new_n965), .ZN(G57));
endmodule


