//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT64), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n202), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n239), .B(new_n245), .ZN(G351));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G107), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G232), .A2(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G238), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(new_n248), .A3(G274), .ZN(new_n267));
  INV_X1    g0067(.A(G244), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n248), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(G200), .B1(new_n263), .B2(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n263), .A2(new_n271), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n216), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  XOR2_X1   g0078(.A(KEYINPUT8), .B(G58), .Z(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n207), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n255), .A2(G20), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT15), .B(G87), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n285), .A2(KEYINPUT67), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n283), .B(new_n290), .C1(new_n207), .C2(new_n284), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n278), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT68), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n295), .A2(new_n206), .A3(G13), .A4(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n277), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n284), .B1(new_n206), .B2(G20), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n299), .A2(new_n284), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n275), .A2(new_n292), .A3(new_n302), .ZN(new_n303));
  OR3_X1    g0103(.A1(new_n263), .A2(G179), .A3(new_n271), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n263), .B2(new_n271), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n288), .A2(new_n286), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n291), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n277), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n311), .B2(new_n301), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n260), .B1(new_n256), .B2(new_n257), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G223), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n258), .A2(G222), .A3(new_n260), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n316), .C1(new_n284), .C2(new_n258), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n270), .ZN(new_n320));
  INV_X1    g0120(.A(G274), .ZN(new_n321));
  AND2_X1   g0121(.A1(G1), .A2(G13), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(new_n247), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n320), .A2(G226), .B1(new_n323), .B2(new_n266), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G200), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n319), .A2(G190), .A3(new_n324), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(KEYINPUT69), .A2(KEYINPUT10), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n293), .A2(G50), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n277), .B1(new_n206), .B2(G20), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(G50), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n203), .A2(G20), .ZN(new_n333));
  INV_X1    g0133(.A(G150), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n207), .A2(new_n255), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G58), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(KEYINPUT8), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT65), .B(G58), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(KEYINPUT8), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n336), .B1(new_n341), .B2(new_n286), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n332), .B1(new_n342), .B2(new_n278), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT9), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n329), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT69), .A2(KEYINPUT10), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(new_n344), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n328), .A2(new_n346), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n326), .A3(new_n327), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n347), .B1(new_n351), .B2(new_n345), .ZN(new_n352));
  INV_X1    g0152(.A(new_n343), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n305), .B2(new_n325), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(G179), .B2(new_n325), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n313), .A2(new_n350), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT70), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n356), .B(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(G223), .B(new_n260), .C1(new_n249), .C2(new_n250), .ZN(new_n359));
  OAI211_X1 g0159(.A(G226), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n318), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n320), .A2(G232), .B1(new_n323), .B2(new_n266), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT75), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT75), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n363), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  INV_X1    g0170(.A(new_n365), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n369), .A2(new_n305), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT65), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(G58), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n337), .A2(KEYINPUT65), .ZN(new_n375));
  OAI21_X1  g0175(.A(G68), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n207), .B1(new_n376), .B2(new_n213), .ZN(new_n377));
  INV_X1    g0177(.A(G159), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n335), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT74), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n256), .A2(new_n207), .A3(new_n257), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n257), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n381), .B1(new_n386), .B2(G68), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n337), .A2(KEYINPUT65), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n373), .A2(G58), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n241), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n390), .B2(new_n201), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT74), .ZN(new_n392));
  INV_X1    g0192(.A(new_n379), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n380), .A2(new_n387), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n393), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n241), .B1(new_n384), .B2(new_n385), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n381), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(new_n277), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n340), .A2(new_n331), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n340), .B2(new_n293), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n372), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n372), .B2(new_n403), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n365), .A2(G190), .ZN(new_n410));
  INV_X1    g0210(.A(G200), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n369), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n409), .B1(new_n412), .B2(new_n403), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n363), .A2(new_n364), .A3(new_n367), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n367), .B1(new_n363), .B2(new_n364), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n410), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n399), .A4(new_n402), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  OR2_X1    g0221(.A1(G226), .A2(G1698), .ZN(new_n422));
  INV_X1    g0222(.A(G232), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G1698), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n422), .B(new_n424), .C1(new_n249), .C2(new_n250), .ZN(new_n425));
  INV_X1    g0225(.A(G97), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n255), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n318), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n248), .A2(G238), .A3(new_n269), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n267), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n421), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(new_n370), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n432), .A3(new_n421), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT71), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n248), .B1(new_n425), .B2(new_n428), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n267), .A2(new_n431), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT13), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT71), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n434), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT13), .B1(new_n438), .B2(new_n439), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT14), .B1(new_n444), .B2(G169), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT14), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n446), .B(new_n305), .C1(new_n435), .C2(new_n443), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n442), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n331), .A2(G68), .A3(new_n297), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT12), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n293), .B2(G68), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n294), .A2(KEYINPUT12), .A3(new_n241), .A4(new_n296), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT73), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT11), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n207), .A2(G33), .A3(G77), .ZN(new_n457));
  OAI221_X1 g0257(.A(new_n457), .B1(new_n207), .B2(G68), .C1(new_n335), .C2(new_n202), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT72), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n458), .A2(new_n459), .A3(new_n277), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n459), .B1(new_n458), .B2(new_n277), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n277), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT72), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n458), .A2(new_n459), .A3(new_n277), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(KEYINPUT11), .A3(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n449), .A2(KEYINPUT73), .A3(new_n451), .A4(new_n452), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n455), .A2(new_n462), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n411), .B1(new_n435), .B2(new_n443), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n437), .A2(new_n441), .A3(G190), .A4(new_n443), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n448), .A2(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n408), .A2(new_n420), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n358), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n258), .A2(G238), .A3(new_n260), .ZN(new_n476));
  OAI211_X1 g0276(.A(G244), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n318), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n206), .A2(G45), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n323), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n248), .A2(G250), .A3(new_n481), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n480), .A2(new_n274), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n479), .B2(new_n318), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(G200), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n278), .B(new_n293), .C1(G1), .C2(new_n255), .ZN(new_n490));
  INV_X1    g0290(.A(G87), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT19), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT78), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT78), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT19), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT79), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n258), .A2(new_n207), .A3(G68), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT79), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n493), .A2(new_n495), .A3(new_n497), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n496), .A2(KEYINPUT19), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n494), .A2(KEYINPUT78), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n427), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(G97), .A2(G107), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n506), .A2(new_n207), .B1(new_n491), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n277), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n298), .A2(new_n287), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n509), .A2(KEYINPUT80), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT80), .B1(new_n509), .B2(new_n510), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n489), .B(new_n492), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n490), .A2(new_n287), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n509), .A2(new_n510), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT80), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n509), .A2(KEYINPUT80), .A3(new_n510), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n480), .A2(new_n486), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n305), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(G179), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n513), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT81), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT81), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n513), .B(new_n525), .C1(new_n519), .C2(new_n522), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT76), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n528), .A2(new_n252), .A3(KEYINPUT6), .A4(G97), .ZN(new_n529));
  NAND2_X1  g0329(.A1(KEYINPUT6), .A2(G97), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT76), .B1(new_n530), .B2(G107), .ZN(new_n531));
  AND2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n507), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n529), .B(new_n531), .C1(new_n533), .C2(KEYINPUT6), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n386), .A2(G107), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n278), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n293), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n426), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n490), .B2(new_n426), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(KEYINPUT5), .B(G41), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n318), .B1(new_n482), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G257), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n323), .A2(new_n482), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(new_n260), .C1(new_n249), .C2(new_n250), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT77), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT4), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT4), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n314), .A2(G250), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G283), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n550), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n546), .B1(new_n555), .B2(new_n318), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n370), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n541), .B(new_n557), .C1(G169), .C2(new_n556), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(G190), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n537), .A2(new_n540), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n411), .C2(new_n556), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n527), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n542), .A2(new_n482), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(G270), .A3(new_n248), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n545), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n314), .A2(G264), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n258), .A2(G257), .A3(new_n260), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n251), .A2(G303), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n318), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G200), .ZN(new_n574));
  INV_X1    g0374(.A(G116), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n206), .B2(G33), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n297), .A2(new_n278), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G116), .B2(new_n297), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n554), .B(new_n207), .C1(G33), .C2(new_n426), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(G20), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n277), .A2(KEYINPUT82), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT82), .B1(new_n277), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(KEYINPUT20), .B(new_n579), .C1(new_n581), .C2(new_n582), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n578), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n574), .B(new_n587), .C1(new_n274), .C2(new_n573), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n573), .A2(G169), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(new_n587), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n585), .A2(new_n586), .ZN(new_n592));
  INV_X1    g0392(.A(new_n578), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n594), .A2(KEYINPUT21), .A3(G169), .A4(new_n573), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n567), .A2(G179), .A3(new_n572), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n588), .A2(new_n591), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(G250), .B(new_n260), .C1(new_n249), .C2(new_n250), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT84), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n258), .A2(new_n602), .A3(G250), .A4(new_n260), .ZN(new_n603));
  NAND2_X1  g0403(.A1(G33), .A2(G294), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n258), .A2(G257), .A3(G1698), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n318), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n564), .A2(G264), .A3(new_n248), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n545), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n305), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n606), .B2(new_n318), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n370), .A3(new_n545), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n207), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n614));
  AND2_X1   g0414(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n615));
  NOR2_X1   g0415(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n258), .A2(new_n207), .A3(G87), .A4(new_n615), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n478), .A2(G20), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT23), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n207), .B2(G107), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n252), .A2(KEYINPUT23), .A3(G20), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT24), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT24), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n618), .A2(new_n619), .A3(new_n624), .A4(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n278), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n538), .A2(KEYINPUT25), .A3(new_n252), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT25), .B1(new_n538), .B2(new_n252), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n490), .A2(new_n252), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n611), .B(new_n613), .C1(new_n629), .C2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n629), .A2(new_n632), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n612), .A2(new_n274), .A3(new_n545), .ZN(new_n635));
  AOI21_X1  g0435(.A(G200), .B1(new_n612), .B2(new_n545), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n633), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n633), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n599), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n475), .A2(new_n563), .A3(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n468), .ZN(new_n643));
  INV_X1    g0443(.A(new_n469), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n471), .A3(new_n644), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n645), .A2(new_n312), .B1(new_n448), .B2(new_n468), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT87), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n420), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  INV_X1    g0449(.A(new_n407), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n405), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n352), .B(new_n350), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n355), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n520), .A2(G179), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n521), .A2(KEYINPUT86), .ZN(new_n656));
  OR3_X1    g0456(.A1(new_n488), .A2(KEYINPUT86), .A3(G169), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI22_X1  g0458(.A1(new_n511), .A2(new_n512), .B1(new_n287), .B2(new_n490), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n591), .A2(new_n595), .A3(new_n597), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n613), .B1(new_n629), .B2(new_n632), .ZN(new_n662));
  INV_X1    g0462(.A(new_n611), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n558), .A2(new_n561), .A3(new_n637), .A4(new_n513), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n660), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n660), .A2(new_n513), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n558), .ZN(new_n670));
  INV_X1    g0470(.A(new_n558), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n524), .A2(KEYINPUT26), .A3(new_n526), .A4(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n667), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n654), .B1(new_n475), .B2(new_n673), .ZN(G369));
  INV_X1    g0474(.A(new_n640), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n633), .A2(new_n637), .A3(new_n638), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT88), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n629), .B2(new_n632), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n677), .A2(new_n686), .B1(new_n664), .B2(new_n685), .ZN(new_n687));
  INV_X1    g0487(.A(new_n685), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n587), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n598), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n661), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(KEYINPUT89), .B(G330), .Z(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n687), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n661), .A2(new_n688), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n677), .A2(new_n698), .B1(new_n664), .B2(new_n688), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n210), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n507), .A2(new_n491), .A3(new_n575), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT90), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n703), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n214), .B2(new_n703), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n673), .B2(new_n685), .ZN(new_n710));
  AND4_X1   g0510(.A1(KEYINPUT26), .A2(new_n671), .A3(new_n660), .A4(new_n513), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n524), .A2(new_n526), .A3(new_n671), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n668), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n688), .C1(new_n713), .C2(new_n667), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n524), .A2(new_n526), .A3(new_n562), .A4(new_n688), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n566), .B1(new_n318), .B2(new_n571), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n612), .A3(G179), .A4(new_n488), .ZN(new_n719));
  INV_X1    g0519(.A(new_n556), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n717), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n718), .A2(G179), .A3(new_n488), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n720), .A3(new_n610), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n612), .A2(new_n488), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(KEYINPUT30), .A3(new_n556), .A4(new_n596), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n716), .B1(new_n726), .B2(new_n685), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n726), .A2(new_n716), .A3(new_n685), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n715), .A2(new_n641), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n710), .A2(new_n714), .B1(new_n694), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n708), .B1(new_n730), .B2(G1), .ZN(G364));
  AND2_X1   g0531(.A1(new_n207), .A2(G13), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n206), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n702), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT91), .Z(new_n736));
  NAND3_X1  g0536(.A1(new_n690), .A2(new_n693), .A3(new_n691), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(new_n695), .B2(new_n737), .ZN(new_n738));
  OR3_X1    g0538(.A1(KEYINPUT92), .A2(G13), .A3(G33), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT92), .B1(G13), .B2(G33), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n216), .B1(G20), .B2(new_n305), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n210), .A2(new_n251), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n265), .B2(new_n215), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n245), .B2(new_n265), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n701), .A2(new_n251), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n750), .A2(G355), .B1(new_n575), .B2(new_n701), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n746), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(G20), .A2(G179), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n274), .A2(new_n411), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n274), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n202), .A2(new_n757), .B1(new_n759), .B2(new_n339), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n207), .A2(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G87), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n411), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n761), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n764), .B(new_n258), .C1(new_n252), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G190), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n755), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n767), .B1(G77), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n758), .A2(new_n370), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n426), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n761), .A2(new_n768), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G159), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n779));
  AOI21_X1  g0579(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n771), .B(new_n780), .C1(new_n778), .C2(new_n779), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n755), .A2(new_n765), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n760), .B(new_n781), .C1(G68), .C2(new_n783), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n786));
  INV_X1    g0586(.A(new_n759), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G311), .A2(new_n770), .B1(new_n787), .B2(G322), .ZN(new_n788));
  INV_X1    g0588(.A(new_n757), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT33), .B(G317), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G326), .A2(new_n789), .B1(new_n783), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G303), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n762), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n251), .B1(new_n766), .B2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n793), .B(new_n795), .C1(G329), .C2(new_n777), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n773), .A2(G294), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n788), .A2(new_n791), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n785), .A2(new_n786), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n752), .B1(new_n799), .B2(new_n744), .ZN(new_n800));
  INV_X1    g0600(.A(new_n743), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n692), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n738), .B1(new_n802), .B2(new_n736), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT96), .Z(G396));
  NAND2_X1  g0604(.A1(new_n672), .A2(new_n670), .ZN(new_n805));
  INV_X1    g0605(.A(new_n667), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n685), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n685), .B1(new_n292), .B2(new_n302), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT100), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n306), .B(new_n304), .C1(new_n292), .C2(new_n302), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(new_n688), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n312), .A2(KEYINPUT100), .A3(new_n685), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n313), .A2(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n807), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n729), .A2(new_n694), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n736), .B1(new_n815), .B2(new_n816), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G137), .A2(new_n789), .B1(new_n783), .B2(G150), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT99), .ZN(new_n821));
  INV_X1    g0621(.A(G143), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n822), .B2(new_n759), .C1(new_n378), .C2(new_n769), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n766), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G68), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n202), .B2(new_n762), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n774), .A2(new_n339), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n776), .A2(new_n831), .ZN(new_n832));
  NOR4_X1   g0632(.A1(new_n829), .A2(new_n830), .A3(new_n251), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n824), .B2(KEYINPUT34), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G107), .A2(new_n763), .B1(new_n827), .B2(G87), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n258), .B1(new_n777), .B2(G311), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(new_n426), .C2(new_n774), .ZN(new_n837));
  XOR2_X1   g0637(.A(KEYINPUT98), .B(G283), .Z(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G116), .A2(new_n770), .B1(new_n783), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G294), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n841), .B2(new_n759), .C1(new_n792), .C2(new_n757), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n826), .A2(new_n834), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n744), .ZN(new_n844));
  INV_X1    g0644(.A(new_n736), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n741), .A2(new_n744), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT97), .Z(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n845), .B1(new_n284), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n741), .B2(new_n813), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n819), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G384));
  OR2_X1    g0653(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n217), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  NAND3_X1  g0657(.A1(new_n215), .A2(G77), .A3(new_n376), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n206), .B(G13), .C1(new_n858), .C2(new_n240), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n448), .A2(new_n468), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n685), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n372), .A2(new_n403), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n418), .A2(new_n399), .A3(new_n402), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n403), .A2(new_n682), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n213), .B1(new_n339), .B2(new_n241), .ZN(new_n868));
  AOI211_X1 g0668(.A(KEYINPUT74), .B(new_n379), .C1(new_n868), .C2(G20), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n392), .B1(new_n391), .B2(new_n393), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n278), .B1(new_n871), .B2(new_n387), .ZN(new_n872));
  INV_X1    g0672(.A(new_n397), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n380), .A2(new_n394), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n381), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n401), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT102), .B1(new_n876), .B2(new_n683), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT16), .B1(new_n871), .B2(new_n873), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n395), .A2(new_n277), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n402), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(new_n682), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n372), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n877), .A2(new_n882), .A3(new_n864), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n867), .B1(new_n884), .B2(KEYINPUT37), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n876), .A2(KEYINPUT102), .A3(new_n683), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n881), .B1(new_n880), .B2(new_n682), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n408), .B2(new_n420), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n413), .A2(new_n419), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n651), .A2(new_n895), .B1(new_n886), .B2(new_n887), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(KEYINPUT103), .B(KEYINPUT39), .C1(new_n891), .C2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n883), .A2(new_n864), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n899), .B1(new_n888), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n896), .B(KEYINPUT38), .C1(new_n901), .C2(new_n867), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n895), .A2(KEYINPUT104), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n413), .A2(new_n905), .A3(new_n419), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n408), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n865), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n907), .A2(new_n908), .B1(new_n893), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n902), .B(new_n903), .C1(new_n910), .C2(KEYINPUT38), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n898), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n890), .B1(new_n885), .B2(new_n889), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n902), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT103), .B1(new_n914), .B2(KEYINPUT39), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n862), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n810), .A2(new_n685), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n807), .B2(new_n814), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n685), .A2(new_n468), .ZN(new_n919));
  OAI21_X1  g0719(.A(G169), .B1(new_n433), .B2(new_n440), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n446), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n444), .A2(KEYINPUT14), .A3(G169), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n438), .A2(new_n439), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT71), .B1(new_n923), .B2(new_n421), .ZN(new_n924));
  NOR4_X1   g0724(.A1(new_n438), .A2(new_n439), .A3(new_n436), .A4(KEYINPUT13), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n921), .A2(new_n922), .B1(new_n926), .B2(new_n434), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n645), .B(new_n919), .C1(new_n927), .C2(new_n643), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT101), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n472), .A2(KEYINPUT101), .A3(new_n919), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n448), .A2(new_n468), .A3(new_n685), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n918), .A2(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n936), .A2(new_n914), .B1(new_n651), .B2(new_n683), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n916), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n710), .A2(new_n714), .A3(new_n474), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT105), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT105), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n710), .A2(new_n714), .A3(new_n474), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n654), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n938), .B(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n891), .A2(new_n897), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n813), .B1(new_n932), .B2(new_n933), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n729), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n946), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n902), .B1(new_n910), .B2(KEYINPUT38), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n948), .A2(KEYINPUT40), .A3(new_n729), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n729), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n954), .B1(new_n475), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n950), .A2(new_n474), .A3(new_n729), .A4(new_n953), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n694), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n945), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n206), .B2(new_n732), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n945), .A2(new_n958), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n860), .B1(new_n960), .B2(new_n961), .ZN(G367));
  OAI21_X1  g0762(.A(new_n562), .B1(new_n560), .B2(new_n688), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n671), .A2(new_n685), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(new_n677), .A3(new_n698), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT42), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n558), .B1(new_n963), .B2(new_n633), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n966), .A2(KEYINPUT42), .B1(new_n688), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n492), .B1(new_n511), .B2(new_n512), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n685), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n660), .A2(new_n513), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n660), .B2(new_n971), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n967), .A2(new_n969), .B1(KEYINPUT43), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n696), .A2(new_n965), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n702), .B(new_n979), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n699), .A2(new_n965), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT45), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT107), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n699), .A2(new_n965), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(KEYINPUT44), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n984), .A2(KEYINPUT44), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n987), .A2(new_n985), .A3(new_n983), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n696), .ZN(new_n990));
  MUX2_X1   g0790(.A(new_n687), .B(new_n677), .S(new_n698), .Z(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(new_n695), .Z(new_n992));
  NAND3_X1  g0792(.A1(new_n986), .A2(new_n697), .A3(new_n988), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n730), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n980), .B1(new_n994), .B2(new_n730), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n978), .B1(new_n995), .B2(new_n734), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n235), .A2(new_n747), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n745), .B1(new_n210), .B2(new_n287), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n841), .A2(new_n782), .B1(new_n759), .B2(new_n792), .ZN(new_n999));
  INV_X1    g0799(.A(G311), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n1000), .A2(new_n757), .B1(new_n769), .B2(new_n838), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n827), .A2(G97), .ZN(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n251), .C1(new_n1004), .C2(new_n776), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT108), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n762), .A2(new_n575), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n774), .A2(new_n252), .B1(new_n1008), .B2(KEYINPUT46), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(KEYINPUT46), .B2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1002), .A2(new_n1007), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n202), .A2(new_n769), .B1(new_n782), .B2(new_n378), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT109), .Z(new_n1014));
  NAND2_X1  g0814(.A1(new_n827), .A2(G77), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n339), .B2(new_n762), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n251), .B(new_n1016), .C1(G137), .C2(new_n777), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n773), .A2(G68), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G143), .A2(new_n789), .B1(new_n787), .B2(G150), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1012), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT110), .Z(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT47), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n744), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n736), .B1(new_n997), .B2(new_n998), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT111), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(KEYINPUT111), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n801), .C2(new_n973), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n996), .A2(new_n1028), .ZN(G387));
  NOR2_X1   g0829(.A1(new_n231), .A2(new_n265), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n750), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1030), .A2(new_n747), .B1(new_n705), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n279), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n1033), .A2(G50), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n1033), .B2(G50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n705), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1032), .A2(new_n1038), .B1(new_n252), .B2(new_n701), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n202), .A2(new_n759), .B1(new_n757), .B2(new_n378), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n241), .A2(new_n769), .B1(new_n782), .B2(new_n340), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n763), .A2(G77), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n777), .A2(G150), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1042), .A2(new_n1003), .A3(new_n1043), .A4(new_n258), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n774), .A2(new_n287), .ZN(new_n1045));
  NOR4_X1   g0845(.A1(new_n1040), .A2(new_n1041), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT113), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n251), .B1(new_n766), .B2(new_n575), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G311), .A2(new_n783), .B1(new_n789), .B2(G322), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n792), .B2(new_n769), .C1(new_n1004), .C2(new_n759), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n773), .A2(new_n839), .B1(new_n763), .B2(G294), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT49), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1048), .B(new_n1057), .C1(G326), .C2(new_n777), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1047), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n736), .B1(new_n746), .B2(new_n1039), .C1(new_n1060), .C2(new_n1024), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n687), .B2(new_n743), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n992), .B2(new_n734), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n992), .A2(new_n730), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n702), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n992), .A2(new_n730), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(G393));
  INV_X1    g0867(.A(KEYINPUT114), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n990), .A2(new_n1068), .A3(new_n993), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n993), .A2(new_n1068), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n1064), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n702), .A3(new_n994), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n965), .A2(new_n801), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1000), .A2(new_n759), .B1(new_n757), .B2(new_n1004), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n251), .B1(new_n766), .B2(new_n252), .ZN(new_n1076));
  INV_X1    g0876(.A(G322), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n838), .A2(new_n762), .B1(new_n776), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(G116), .C2(new_n773), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G294), .A2(new_n770), .B1(new_n783), .B2(G303), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1075), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n334), .A2(new_n757), .B1(new_n759), .B2(new_n378), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n774), .A2(new_n284), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n258), .B1(new_n766), .B2(new_n491), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n762), .A2(new_n241), .B1(new_n776), .B2(new_n822), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G50), .A2(new_n783), .B1(new_n770), .B2(new_n279), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1083), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1024), .B1(new_n1081), .B2(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n745), .B1(new_n426), .B2(new_n210), .C1(new_n239), .C2(new_n747), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n736), .A2(new_n1091), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1073), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n734), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT115), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1072), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1072), .B2(new_n1095), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G390));
  AND2_X1   g0900(.A1(new_n729), .A2(G330), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n934), .B1(new_n1101), .B2(new_n814), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n688), .B(new_n814), .C1(new_n713), .C2(new_n667), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n729), .A2(new_n934), .A3(new_n814), .A4(new_n694), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n917), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT116), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n729), .A2(new_n814), .A3(new_n694), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1101), .A2(new_n948), .B1(new_n1109), .B2(new_n935), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1110), .B2(new_n918), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n935), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n948), .A2(G330), .A3(new_n729), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n918), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1115), .A3(KEYINPUT116), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1107), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1101), .A2(new_n474), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n943), .A2(new_n1119), .A3(new_n654), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT103), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n947), .B2(new_n903), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n862), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n918), .B2(new_n935), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1123), .A2(new_n1125), .A3(new_n911), .A4(new_n898), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n934), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1128), .A2(new_n1124), .A3(new_n951), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1126), .A2(new_n1104), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n951), .A2(new_n1124), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n934), .B2(new_n1127), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n912), .A2(new_n915), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n1125), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1121), .B(new_n1130), .C1(new_n1134), .C2(new_n1113), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1107), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1110), .A2(new_n1108), .A3(new_n918), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT116), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1118), .B(new_n653), .C1(new_n940), .C2(new_n942), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1130), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1113), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1135), .A2(new_n1144), .A3(new_n702), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n734), .B(new_n1130), .C1(new_n1134), .C2(new_n1113), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT120), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1133), .A2(new_n741), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n762), .B2(new_n334), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n763), .A2(G150), .A3(new_n1149), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(new_n378), .C2(new_n774), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n769), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n251), .B1(new_n777), .B2(G125), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n202), .B2(new_n766), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1153), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G128), .A2(new_n789), .B1(new_n787), .B2(G132), .ZN(new_n1159));
  INV_X1    g0959(.A(G137), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(new_n1159), .C1(new_n1160), .C2(new_n782), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G107), .A2(new_n783), .B1(new_n789), .B2(G283), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n426), .B2(new_n769), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT118), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n777), .A2(G294), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n764), .A2(new_n828), .A3(new_n1165), .A4(new_n251), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1166), .A2(new_n1084), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n575), .B2(new_n759), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1161), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT119), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1024), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1170), .B2(new_n1169), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n845), .B1(new_n340), .B2(new_n848), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1148), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1146), .A2(new_n1147), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1147), .B1(new_n1146), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1145), .B1(new_n1175), .B2(new_n1176), .ZN(G378));
  INV_X1    g0977(.A(KEYINPUT122), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n949), .B1(new_n902), .B2(new_n913), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n953), .B(G330), .C1(new_n1179), .C2(KEYINPUT40), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n350), .A2(new_n352), .A3(new_n355), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n353), .A2(new_n683), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1185), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n950), .A2(G330), .A3(new_n953), .A4(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1186), .A2(new_n916), .A3(new_n1188), .A4(new_n937), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1186), .A2(new_n1188), .B1(new_n916), .B2(new_n937), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1178), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n938), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(KEYINPUT122), .A3(new_n1189), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1192), .A2(new_n734), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1187), .A2(new_n742), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n846), .A2(new_n202), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n773), .A2(G150), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n762), .B2(new_n1154), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G125), .A2(new_n789), .B1(new_n787), .B2(G128), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n831), .B2(new_n782), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G137), .C2(new_n770), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(G33), .A2(G41), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT121), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n766), .A2(new_n378), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(G124), .C2(new_n777), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1205), .A2(new_n1206), .A3(new_n1210), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n252), .A2(new_n759), .B1(new_n769), .B2(new_n287), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n426), .A2(new_n782), .B1(new_n757), .B2(new_n575), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n766), .A2(new_n339), .B1(new_n776), .B2(new_n794), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n258), .A2(G41), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1215), .A2(new_n1018), .A3(new_n1042), .A4(new_n1216), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1212), .A2(new_n1213), .A3(new_n1217), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT58), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(KEYINPUT58), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1208), .B(new_n202), .C1(G41), .C2(new_n258), .ZN(new_n1221));
  AND4_X1   g1021(.A1(new_n1211), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n736), .B(new_n1198), .C1(new_n1222), .C2(new_n1024), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1197), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1196), .A2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1130), .B1(new_n1134), .B2(new_n1113), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1140), .B1(new_n1227), .B2(new_n1141), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n1195), .A3(new_n1192), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT57), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1194), .B2(new_n1189), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n703), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1226), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(G375));
  AOI21_X1  g1035(.A(new_n845), .B1(new_n241), .B2(new_n848), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n252), .A2(new_n769), .B1(new_n759), .B2(new_n794), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n575), .A2(new_n782), .B1(new_n757), .B2(new_n841), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1015), .A2(new_n251), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n762), .A2(new_n426), .B1(new_n776), .B2(new_n792), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1045), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1160), .A2(new_n759), .B1(new_n769), .B2(new_n334), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n831), .A2(new_n757), .B1(new_n782), .B2(new_n1154), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n258), .B1(new_n766), .B2(new_n339), .ZN(new_n1246));
  INV_X1    g1046(.A(G128), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n762), .A2(new_n378), .B1(new_n776), .B2(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(G50), .C2(new_n773), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1239), .A2(new_n1242), .B1(new_n1245), .B2(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1236), .B1(new_n1024), .B2(new_n1250), .C1(new_n934), .C2(new_n742), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1139), .B2(new_n734), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1121), .A2(new_n980), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1254), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(G381));
  AND2_X1   g1059(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1260), .A2(new_n1261), .A3(G378), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(G387), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1099), .A3(new_n1258), .A4(new_n1263), .ZN(G407));
  NAND2_X1  g1064(.A1(new_n684), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G407), .A2(G213), .A3(new_n1267), .ZN(G409));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1194), .A2(KEYINPUT122), .A3(new_n1189), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT122), .B1(new_n1194), .B2(new_n1189), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1224), .B1(new_n1272), .B2(new_n734), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT57), .B1(new_n1272), .B2(new_n1228), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1233), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G378), .B(new_n1273), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G378), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1194), .A2(new_n1189), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1224), .B1(new_n1278), .B2(new_n734), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1229), .B2(new_n980), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1266), .B1(new_n1276), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT60), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(new_n1256), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1117), .A2(new_n1120), .A3(KEYINPUT60), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n702), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1253), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n852), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G384), .B(new_n1253), .C1(new_n1285), .C2(new_n1287), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1266), .A2(G2897), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1289), .A2(new_n1290), .A3(new_n1292), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT124), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT124), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1289), .A2(new_n1296), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1282), .A2(new_n1293), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1269), .B1(new_n1299), .B2(KEYINPUT61), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1276), .A2(new_n1281), .ZN(new_n1301));
  OR2_X1    g1101(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(new_n1265), .A3(new_n1291), .A4(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1282), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1291), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  XOR2_X1   g1107(.A(G393), .B(G396), .Z(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1099), .A2(G387), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1099), .A2(G387), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1309), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1312), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1293), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n980), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1272), .A2(new_n1319), .A3(new_n1228), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G378), .B1(new_n1320), .B2(new_n1279), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(G378), .B2(new_n1234), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1317), .B(new_n1318), .C1(new_n1322), .C2(new_n1266), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(KEYINPUT125), .A3(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1300), .A2(new_n1307), .A3(new_n1316), .A4(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1282), .A2(new_n1291), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1282), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1329), .A2(new_n1324), .A3(new_n1323), .A4(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1316), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1326), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(KEYINPUT127), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1326), .A2(new_n1333), .A3(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(G405));
  XNOR2_X1  g1138(.A(new_n1234), .B(G378), .ZN(new_n1339));
  XOR2_X1   g1139(.A(new_n1339), .B(new_n1291), .Z(new_n1340));
  XNOR2_X1  g1140(.A(new_n1340), .B(new_n1332), .ZN(G402));
endmodule


