//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XOR2_X1   g002(.A(G211gat), .B(G218gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT22), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n206), .B(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G141gat), .B(G148gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n215), .B1(G155gat), .B2(G162gat), .ZN(new_n216));
  AND2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  OAI22_X1  g016(.A1(new_n214), .A2(new_n216), .B1(KEYINPUT75), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n218), .A2(new_n220), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n213), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G228gat), .A2(G233gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n221), .A2(new_n222), .ZN(new_n232));
  INV_X1    g031(.A(new_n213), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n229), .B(new_n231), .C1(new_n232), .C2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n207), .A2(KEYINPUT81), .A3(new_n211), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n204), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT81), .B1(new_n207), .B2(new_n211), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n228), .B1(new_n238), .B2(new_n239), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n225), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT82), .ZN(new_n243));
  OR3_X1    g042(.A1(new_n242), .A2(new_n243), .A3(new_n232), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n242), .B2(new_n232), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n229), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n230), .B(KEYINPUT80), .Z(new_n248));
  AND3_X1   g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n236), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G22gat), .ZN(new_n252));
  INV_X1    g051(.A(G22gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n253), .B(new_n236), .C1(new_n249), .C2(new_n250), .ZN(new_n254));
  XNOR2_X1  g053(.A(G78gat), .B(G106gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(KEYINPUT79), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n252), .B2(new_n254), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n203), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n252), .A2(new_n254), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n256), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(new_n202), .A3(new_n258), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G127gat), .B(G134gat), .Z(new_n266));
  XNOR2_X1  g065(.A(G113gat), .B(G120gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n266), .B1(KEYINPUT1), .B2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n268), .B(KEYINPUT67), .Z(new_n269));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270));
  INV_X1    g069(.A(G120gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(G113gat), .ZN(new_n272));
  INV_X1    g071(.A(G113gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n272), .B(new_n274), .C1(new_n273), .C2(G120gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n269), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT23), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(G169gat), .ZN(new_n286));
  INV_X1    g085(.A(G176gat), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n283), .B(new_n285), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT24), .B1(new_n291), .B2(KEYINPUT64), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(KEYINPUT64), .B2(new_n291), .ZN(new_n293));
  INV_X1    g092(.A(G183gat), .ZN(new_n294));
  INV_X1    g093(.A(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n297), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n291), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n289), .B1(new_n302), .B2(new_n288), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n299), .A2(new_n303), .A3(KEYINPUT65), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n295), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n282), .A2(KEYINPUT26), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n286), .B2(new_n287), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n282), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n312), .A2(new_n313), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n281), .B1(new_n308), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(G227gat), .A2(G233gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n306), .B2(new_n307), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n280), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT32), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT70), .B(G71gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(G99gat), .ZN(new_n326));
  XOR2_X1   g125(.A(G15gat), .B(G43gat), .Z(new_n327));
  XOR2_X1   g126(.A(new_n326), .B(new_n327), .Z(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT33), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n320), .B1(new_n319), .B2(new_n322), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT34), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI211_X1 g133(.A(KEYINPUT34), .B(new_n320), .C1(new_n319), .C2(new_n322), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n331), .A2(new_n334), .A3(new_n335), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n324), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n331), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n332), .A2(new_n333), .ZN(new_n341));
  INV_X1    g140(.A(new_n335), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n324), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n336), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n339), .A2(KEYINPUT87), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT87), .B1(new_n339), .B2(new_n345), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n269), .A2(new_n232), .A3(new_n279), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n232), .A2(new_n224), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n280), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n269), .A2(new_n232), .A3(KEYINPUT4), .A4(new_n279), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n355), .A2(KEYINPUT5), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n354), .A3(new_n357), .ZN(new_n359));
  INV_X1    g158(.A(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n280), .A2(new_n223), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n356), .B1(new_n361), .B2(new_n349), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT5), .ZN(new_n363));
  OAI22_X1  g162(.A1(new_n359), .A2(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G1gat), .B(G29gat), .Z(new_n366));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT6), .B1(new_n365), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n358), .A2(new_n364), .A3(new_n370), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT85), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n364), .A3(new_n375), .A4(new_n370), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n372), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(new_n373), .ZN(new_n379));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n304), .A2(new_n317), .ZN(new_n384));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n385), .B(KEYINPUT72), .Z(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT74), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n386), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n321), .B2(new_n228), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n233), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n321), .A2(new_n393), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n386), .B1(new_n384), .B2(new_n234), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n396), .A2(new_n213), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n383), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n394), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n213), .B1(new_n400), .B2(new_n391), .ZN(new_n401));
  INV_X1    g200(.A(new_n398), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n382), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n403), .A3(KEYINPUT30), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n395), .A2(new_n398), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n382), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n409));
  AND2_X1   g208(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n379), .B(new_n408), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n265), .A2(new_n348), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n408), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n373), .A2(new_n378), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n372), .A2(new_n373), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n372), .A2(KEYINPUT78), .A3(new_n373), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n343), .A2(new_n344), .A3(new_n336), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n344), .B1(new_n343), .B2(new_n336), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n420), .A2(new_n261), .A3(new_n264), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT35), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n413), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n261), .A2(new_n264), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n418), .A2(new_n419), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n408), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(KEYINPUT36), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT36), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n421), .B2(new_n422), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n427), .A2(new_n429), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n374), .A2(new_n376), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n415), .B1(new_n434), .B2(new_n372), .ZN(new_n435));
  INV_X1    g234(.A(new_n399), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT37), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n382), .A2(new_n437), .ZN(new_n438));
  OAI22_X1  g237(.A1(new_n436), .A2(new_n438), .B1(new_n405), .B2(new_n437), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT38), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n396), .A2(new_n397), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT86), .B1(new_n441), .B2(new_n233), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n392), .A2(new_n394), .A3(new_n233), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n441), .A2(KEYINPUT86), .A3(new_n233), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT37), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT38), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n446), .B(new_n447), .C1(new_n436), .C2(new_n438), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n435), .A2(new_n440), .A3(new_n403), .A4(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n361), .A2(new_n356), .A3(new_n349), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT84), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n359), .A2(new_n360), .ZN(new_n453));
  OR3_X1    g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n370), .B1(new_n453), .B2(new_n452), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT40), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(KEYINPUT40), .A3(new_n455), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n414), .A2(new_n458), .A3(new_n434), .A4(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n449), .A2(new_n264), .A3(new_n261), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n433), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n426), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G113gat), .B(G141gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(G169gat), .B(G197gat), .Z(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT12), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT93), .ZN(new_n471));
  INV_X1    g270(.A(G1gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n253), .A2(G15gat), .ZN(new_n473));
  INV_X1    g272(.A(G15gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G22gat), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT91), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT91), .B1(new_n473), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n475), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT91), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n472), .A2(KEYINPUT16), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI211_X1 g283(.A(KEYINPUT92), .B(G8gat), .C1(new_n478), .C2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n488));
  AND4_X1   g287(.A1(new_n487), .A2(new_n478), .A3(new_n484), .A4(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n471), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G36gat), .ZN(new_n491));
  AND2_X1   g290(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G29gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498));
  OR2_X1    g297(.A1(G43gat), .A2(G50gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(G43gat), .A2(G50gat), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n504));
  OR2_X1    g303(.A1(KEYINPUT90), .A2(G50gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(KEYINPUT90), .A2(G50gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n504), .B1(new_n507), .B2(G43gat), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n501), .B1(new_n508), .B2(new_n497), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n478), .A2(new_n484), .A3(new_n488), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n486), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n478), .A2(new_n484), .A3(new_n487), .A4(new_n488), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(KEYINPUT93), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n490), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n508), .A2(new_n497), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n502), .B1(new_n517), .B2(new_n501), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT17), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n510), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n519), .B(new_n521), .C1(new_n485), .C2(new_n489), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n512), .A2(KEYINPUT93), .A3(new_n513), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT93), .B1(new_n512), .B2(new_n513), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n518), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n515), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n516), .B(KEYINPUT13), .Z(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n523), .A2(KEYINPUT94), .A3(new_n524), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n515), .A2(KEYINPUT18), .A3(new_n522), .A4(new_n516), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n470), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n533), .A2(new_n525), .A3(new_n469), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n536), .B(KEYINPUT95), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G57gat), .B(G64gat), .Z(new_n544));
  INV_X1    g343(.A(KEYINPUT9), .ZN(new_n545));
  INV_X1    g344(.A(G71gat), .ZN(new_n546));
  INV_X1    g345(.A(G78gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G71gat), .B(G78gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n544), .A2(new_n550), .A3(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n528), .B2(new_n529), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT98), .B(KEYINPUT19), .Z(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n557), .B(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G127gat), .B(G155gat), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT20), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT97), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n564), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n562), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT7), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n572), .A2(new_n575), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G99gat), .B(G106gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n571), .B1(new_n576), .B2(new_n577), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n585), .A2(new_n581), .A3(new_n575), .A4(new_n579), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n575), .A2(new_n579), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n588), .A2(KEYINPUT99), .A3(new_n581), .A4(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT100), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(KEYINPUT100), .A3(new_n589), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n510), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n519), .A2(new_n521), .A3(new_n592), .A4(new_n593), .ZN(new_n596));
  AND2_X1   g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT41), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G190gat), .B(G218gat), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n597), .A2(KEYINPUT41), .ZN(new_n602));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n600), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n595), .A2(new_n596), .A3(new_n605), .A4(new_n598), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n601), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n604), .B1(new_n601), .B2(new_n606), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n570), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n552), .A2(new_n553), .A3(new_n586), .A4(new_n583), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n555), .B2(new_n590), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G120gat), .B(G148gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT103), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n621), .B(new_n611), .C1(new_n555), .C2(new_n590), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n554), .A2(new_n621), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n587), .A2(KEYINPUT100), .A3(new_n589), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT100), .B1(new_n587), .B2(new_n589), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(KEYINPUT101), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n623), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n613), .B1(new_n631), .B2(KEYINPUT102), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n633));
  AOI211_X1 g432(.A(new_n633), .B(new_n623), .C1(new_n629), .C2(new_n630), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n615), .B(new_n620), .C1(new_n632), .C2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n615), .B1(new_n631), .B2(new_n614), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n619), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n463), .A2(new_n543), .A3(new_n610), .A4(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(new_n428), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(new_n472), .ZN(G1324gat));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n414), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n644), .A2(G8gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT16), .B(G8gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(KEYINPUT42), .B2(new_n647), .ZN(G1325gat));
  AOI21_X1  g448(.A(G15gat), .B1(new_n643), .B2(new_n348), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n430), .A2(new_n432), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n474), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT104), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n650), .B1(new_n643), .B2(new_n653), .ZN(G1326gat));
  OR3_X1    g453(.A1(new_n640), .A2(KEYINPUT105), .A3(new_n265), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT105), .B1(new_n640), .B2(new_n265), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  AOI22_X1  g458(.A1(new_n425), .A2(new_n413), .B1(new_n433), .B2(new_n461), .ZN(new_n660));
  INV_X1    g459(.A(new_n543), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n639), .A2(new_n570), .ZN(new_n663));
  INV_X1    g462(.A(new_n609), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT106), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n667), .A2(G29gat), .A3(new_n428), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT45), .Z(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n660), .B2(new_n664), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n463), .A2(KEYINPUT44), .A3(new_n609), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n661), .A2(new_n663), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675), .B2(new_n428), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n669), .A2(new_n676), .ZN(G1328gat));
  NOR3_X1   g476(.A1(new_n667), .A2(G36gat), .A3(new_n408), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT46), .ZN(new_n679));
  OAI21_X1  g478(.A(G36gat), .B1(new_n675), .B2(new_n408), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(G1329gat));
  NAND3_X1  g480(.A1(new_n662), .A2(new_n348), .A3(new_n666), .ZN(new_n682));
  INV_X1    g481(.A(G43gat), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n682), .A2(new_n683), .B1(new_n684), .B2(KEYINPUT47), .ZN(new_n685));
  INV_X1    g484(.A(new_n651), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(G43gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n675), .B2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n684), .A2(KEYINPUT47), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1330gat));
  OAI211_X1 g489(.A(new_n505), .B(new_n506), .C1(new_n667), .C2(new_n265), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n427), .A2(new_n507), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n675), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g493(.A1(new_n463), .A2(new_n661), .A3(new_n610), .A4(new_n638), .ZN(new_n695));
  INV_X1    g494(.A(new_n428), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g497(.A(new_n408), .B(KEYINPUT108), .Z(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n702), .B(new_n703), .Z(G1333gat));
  AOI21_X1  g503(.A(new_n546), .B1(new_n695), .B2(new_n686), .ZN(new_n705));
  INV_X1    g504(.A(new_n348), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(G71gat), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n695), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g508(.A1(new_n695), .A2(new_n427), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G78gat), .ZN(G1335gat));
  INV_X1    g510(.A(new_n570), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n543), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n638), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT109), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n673), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G85gat), .B1(new_n716), .B2(new_n428), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n427), .A2(new_n429), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n461), .A2(new_n718), .A3(new_n651), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n411), .A2(new_n346), .A3(new_n347), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n720), .A2(new_n265), .B1(new_n424), .B2(KEYINPUT35), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n609), .B(new_n713), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n664), .B1(new_n426), .B2(new_n462), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT51), .B1(new_n725), .B2(new_n713), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n724), .A2(new_n726), .A3(KEYINPUT110), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT110), .B1(new_n724), .B2(new_n726), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n638), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n696), .A2(new_n576), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n717), .B1(new_n729), .B2(new_n730), .ZN(G1336gat));
  NOR2_X1   g530(.A1(new_n700), .A2(G92gat), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n638), .B(new_n732), .C1(new_n724), .C2(new_n726), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n671), .A2(new_n672), .A3(new_n414), .A4(new_n715), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(G92gat), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT52), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n723), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n725), .A2(KEYINPUT51), .A3(new_n713), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n639), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT52), .B1(new_n740), .B2(new_n732), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n671), .A2(new_n672), .A3(new_n699), .A4(new_n715), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G92gat), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT111), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745));
  AND4_X1   g544(.A1(KEYINPUT111), .A2(new_n733), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n737), .B1(new_n744), .B2(new_n746), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n716), .B2(new_n651), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n706), .A2(G99gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n729), .B2(new_n749), .ZN(G1338gat));
  NOR2_X1   g549(.A1(new_n265), .A2(G106gat), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n671), .A2(new_n672), .A3(new_n427), .A4(new_n715), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n740), .A2(new_n751), .B1(new_n752), .B2(G106gat), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1339gat));
  NOR2_X1   g554(.A1(new_n632), .A2(new_n634), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n620), .A2(new_n615), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n631), .A2(new_n614), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n620), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n622), .A2(new_n614), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n629), .B2(new_n630), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n760), .B1(new_n763), .B2(KEYINPUT112), .ZN(new_n764));
  INV_X1    g563(.A(new_n762), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT101), .B1(new_n594), .B2(new_n624), .ZN(new_n766));
  INV_X1    g565(.A(new_n630), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n761), .B1(new_n756), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n758), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n631), .A2(KEYINPUT54), .A3(new_n614), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n776), .A2(new_n773), .A3(new_n620), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n770), .B(new_n764), .C1(new_n632), .C2(new_n634), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n777), .A2(new_n778), .A3(new_n775), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n774), .B(new_n543), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n532), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n530), .A2(new_n515), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT114), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n530), .A2(new_n515), .A3(new_n785), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n515), .A2(new_n522), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(G229gat), .A3(G233gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n784), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n540), .A2(new_n541), .B1(new_n789), .B2(new_n468), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n638), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n781), .A2(KEYINPUT116), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT116), .B1(new_n781), .B2(new_n791), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(new_n609), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n780), .A2(new_n779), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n789), .A2(new_n468), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n542), .A2(new_n609), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n795), .A2(KEYINPUT115), .A3(new_n774), .A4(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n774), .B(new_n797), .C1(new_n779), .C2(new_n780), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n570), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n610), .A2(new_n639), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n543), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n427), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n699), .A2(new_n428), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n348), .A3(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n809), .A2(new_n273), .A3(new_n661), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n781), .A2(new_n791), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n609), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n781), .A2(KEYINPUT116), .A3(new_n791), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n802), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n806), .B1(new_n815), .B2(new_n712), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n427), .A2(new_n421), .A3(new_n422), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n696), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n543), .A3(new_n700), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n810), .B1(new_n820), .B2(new_n273), .ZN(G1340gat));
  OAI21_X1  g620(.A(G120gat), .B1(new_n809), .B2(new_n639), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n700), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n638), .A2(new_n271), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT117), .ZN(G1341gat));
  OAI21_X1  g625(.A(G127gat), .B1(new_n809), .B2(new_n570), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n570), .A2(G127gat), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n823), .B2(new_n828), .ZN(G1342gat));
  INV_X1    g628(.A(G134gat), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n414), .A2(new_n664), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n819), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n809), .B2(new_n664), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n686), .A2(new_n265), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n816), .A2(new_n696), .A3(new_n837), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n661), .A2(G141gat), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n838), .A2(new_n699), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n791), .A2(KEYINPUT118), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n790), .A2(new_n638), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n781), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n664), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n801), .A3(new_n798), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n805), .B1(new_n848), .B2(new_n570), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT57), .B1(new_n849), .B2(new_n265), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n811), .A2(new_n812), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n664), .A3(new_n814), .ZN(new_n853));
  INV_X1    g652(.A(new_n802), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n712), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n851), .B(new_n427), .C1(new_n855), .C2(new_n805), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n808), .A2(new_n651), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n850), .A2(new_n856), .A3(new_n543), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT58), .B1(new_n858), .B2(G141gat), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n841), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n858), .A2(new_n862), .A3(G141gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n858), .B2(G141gat), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n863), .A2(new_n864), .A3(new_n840), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(G1344gat));
  NOR2_X1   g666(.A1(new_n838), .A2(new_n699), .ZN(new_n868));
  INV_X1    g667(.A(G148gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n638), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT121), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n850), .A2(new_n856), .A3(new_n857), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n639), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(KEYINPUT59), .A3(new_n869), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n427), .A2(new_n851), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n847), .A2(new_n799), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n570), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(new_n806), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n427), .B1(new_n855), .B2(new_n805), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(KEYINPUT57), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n638), .A3(new_n857), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n875), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n871), .B1(new_n874), .B2(new_n883), .ZN(G1345gat));
  OAI21_X1  g683(.A(G155gat), .B1(new_n872), .B2(new_n570), .ZN(new_n885));
  INV_X1    g684(.A(new_n868), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n570), .A2(G155gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n872), .B2(new_n664), .ZN(new_n889));
  INV_X1    g688(.A(new_n831), .ZN(new_n890));
  OR3_X1    g689(.A1(new_n838), .A2(G162gat), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n696), .A2(new_n408), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(new_n348), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n807), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n896), .A2(new_n286), .A3(new_n661), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n696), .B1(new_n803), .B2(new_n806), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n817), .A3(new_n699), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n543), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n897), .B1(new_n901), .B2(new_n286), .ZN(G1348gat));
  OAI21_X1  g701(.A(G176gat), .B1(new_n896), .B2(new_n639), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n638), .A2(new_n287), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n899), .B2(new_n904), .ZN(G1349gat));
  NAND3_X1  g704(.A1(new_n900), .A2(new_n309), .A3(new_n712), .ZN(new_n906));
  OAI21_X1  g705(.A(G183gat), .B1(new_n896), .B2(new_n570), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT60), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n906), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n900), .A2(new_n295), .A3(new_n609), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n807), .A2(new_n609), .A3(new_n895), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n916));
  AND4_X1   g715(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(G190gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n295), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n915), .A2(new_n918), .B1(new_n914), .B2(new_n916), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n913), .B1(new_n917), .B2(new_n919), .ZN(G1351gat));
  AOI21_X1  g719(.A(new_n851), .B1(new_n816), .B2(new_n427), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT124), .B1(new_n921), .B2(new_n879), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  INV_X1    g722(.A(new_n879), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n265), .B1(new_n803), .B2(new_n806), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n851), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n894), .A2(new_n651), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n922), .A2(new_n926), .A3(new_n543), .A4(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n927), .B1(new_n881), .B2(new_n923), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n932), .A2(KEYINPUT125), .A3(new_n543), .A4(new_n922), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(G197gat), .A3(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n686), .A2(new_n265), .A3(new_n700), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n898), .A2(new_n935), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n936), .A2(G197gat), .A3(new_n661), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(G1352gat));
  INV_X1    g737(.A(new_n936), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  AOI21_X1  g739(.A(G204gat), .B1(new_n940), .B2(KEYINPUT62), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n638), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n940), .A2(KEYINPUT62), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n932), .A2(new_n922), .ZN(new_n945));
  OAI21_X1  g744(.A(G204gat), .B1(new_n945), .B2(new_n639), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n939), .A2(new_n209), .A3(new_n712), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n928), .A2(new_n712), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n921), .A2(new_n879), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n209), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n949), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n881), .B2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n957), .A2(new_n951), .A3(new_n924), .A4(new_n953), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G211gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(new_n954), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n948), .B1(new_n956), .B2(new_n961), .ZN(G1354gat));
  NOR3_X1   g761(.A1(new_n945), .A2(new_n210), .A3(new_n664), .ZN(new_n963));
  AOI21_X1  g762(.A(G218gat), .B1(new_n939), .B2(new_n609), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


