

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756;

  OR2_X1 U369 ( .A1(n512), .A2(n507), .ZN(n566) );
  XNOR2_X2 U370 ( .A(n426), .B(n425), .ZN(n731) );
  INV_X1 U371 ( .A(G953), .ZN(n750) );
  XNOR2_X2 U372 ( .A(n406), .B(n483), .ZN(n745) );
  XNOR2_X2 U373 ( .A(n663), .B(G146), .ZN(n431) );
  XNOR2_X2 U374 ( .A(n412), .B(n636), .ZN(n495) );
  NOR2_X1 U375 ( .A1(n756), .A2(n755), .ZN(n565) );
  OR2_X2 U376 ( .A1(n638), .A2(G902), .ZN(n412) );
  INV_X1 U377 ( .A(n724), .ZN(n348) );
  XNOR2_X1 U378 ( .A(n370), .B(n369), .ZN(n368) );
  NAND2_X1 U379 ( .A1(n372), .A2(n371), .ZN(n370) );
  NOR2_X1 U380 ( .A1(n588), .A2(n587), .ZN(n371) );
  AND2_X1 U381 ( .A1(n627), .A2(n609), .ZN(n530) );
  XNOR2_X1 U382 ( .A(n565), .B(KEYINPUT46), .ZN(n372) );
  AND2_X1 U383 ( .A1(n378), .A2(n384), .ZN(n383) );
  NOR2_X1 U384 ( .A1(n691), .A2(n495), .ZN(n497) );
  XNOR2_X2 U385 ( .A(n407), .B(G104), .ZN(n732) );
  XNOR2_X2 U386 ( .A(G110), .B(G107), .ZN(n407) );
  XNOR2_X1 U387 ( .A(n746), .B(n364), .ZN(n395) );
  XNOR2_X1 U388 ( .A(n366), .B(n365), .ZN(n364) );
  NOR2_X1 U389 ( .A1(n380), .A2(n379), .ZN(n552) );
  NAND2_X1 U390 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U391 ( .A1(n383), .A2(n350), .ZN(n379) );
  INV_X1 U392 ( .A(KEYINPUT22), .ZN(n356) );
  NAND2_X1 U393 ( .A1(n348), .A2(G217), .ZN(n377) );
  NAND2_X1 U394 ( .A1(n348), .A2(G210), .ZN(n361) );
  NAND2_X1 U395 ( .A1(n586), .A2(n388), .ZN(n587) );
  XNOR2_X1 U396 ( .A(KEYINPUT77), .B(n584), .ZN(n586) );
  INV_X1 U397 ( .A(KEYINPUT48), .ZN(n369) );
  XNOR2_X1 U398 ( .A(n392), .B(n391), .ZN(n366) );
  XNOR2_X1 U399 ( .A(n390), .B(KEYINPUT73), .ZN(n365) );
  XNOR2_X1 U400 ( .A(G128), .B(G137), .ZN(n390) );
  XNOR2_X1 U401 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U402 ( .A(n431), .B(G140), .ZN(n367) );
  AND2_X1 U403 ( .A1(n572), .A2(n387), .ZN(n591) );
  NAND2_X1 U404 ( .A1(n558), .A2(KEYINPUT72), .ZN(n384) );
  XNOR2_X1 U405 ( .A(n550), .B(n385), .ZN(n378) );
  XNOR2_X1 U406 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n385) );
  NAND2_X1 U407 ( .A1(n549), .A2(KEYINPUT72), .ZN(n382) );
  OR2_X1 U408 ( .A1(n549), .A2(n349), .ZN(n381) );
  XNOR2_X1 U409 ( .A(n475), .B(n474), .ZN(n512) );
  OR2_X1 U410 ( .A1(n525), .A2(n524), .ZN(n526) );
  OR2_X1 U411 ( .A1(n517), .A2(n575), .ZN(n518) );
  INV_X1 U412 ( .A(KEYINPUT124), .ZN(n373) );
  XNOR2_X1 U413 ( .A(n361), .B(n354), .ZN(n360) );
  OR2_X1 U414 ( .A1(n558), .A2(KEYINPUT72), .ZN(n349) );
  XNOR2_X1 U415 ( .A(KEYINPUT38), .B(n593), .ZN(n350) );
  OR2_X1 U416 ( .A1(G953), .A2(G237), .ZN(n351) );
  BUF_X1 U417 ( .A(n551), .Z(n593) );
  AND2_X1 U418 ( .A1(n382), .A2(n383), .ZN(n352) );
  XOR2_X1 U419 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n353) );
  XOR2_X1 U420 ( .A(n626), .B(n625), .Z(n354) );
  XNOR2_X1 U421 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n355) );
  AND2_X1 U422 ( .A1(n608), .A2(G953), .ZN(n730) );
  INV_X1 U423 ( .A(n730), .ZN(n359) );
  INV_X1 U424 ( .A(n516), .ZN(n529) );
  XNOR2_X2 U425 ( .A(n357), .B(n356), .ZN(n516) );
  NAND2_X2 U426 ( .A1(n514), .A2(n513), .ZN(n357) );
  XNOR2_X2 U427 ( .A(n462), .B(n461), .ZN(n514) );
  XNOR2_X1 U428 ( .A(n358), .B(n355), .ZN(G51) );
  NAND2_X1 U429 ( .A1(n360), .A2(n359), .ZN(n358) );
  XNOR2_X2 U430 ( .A(n363), .B(n362), .ZN(n426) );
  XNOR2_X2 U431 ( .A(KEYINPUT3), .B(G119), .ZN(n362) );
  XNOR2_X2 U432 ( .A(G116), .B(G113), .ZN(n363) );
  AND2_X2 U433 ( .A1(n668), .A2(n544), .ZN(n601) );
  XNOR2_X2 U434 ( .A(n430), .B(G134), .ZN(n483) );
  XNOR2_X2 U435 ( .A(n367), .B(n389), .ZN(n746) );
  NAND2_X2 U436 ( .A1(n368), .A2(n599), .ZN(n667) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(G66) );
  NAND2_X1 U438 ( .A1(n375), .A2(n359), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n375) );
  INV_X1 U440 ( .A(n607), .ZN(n376) );
  NAND2_X1 U441 ( .A1(n352), .A2(n381), .ZN(n579) );
  XNOR2_X1 U442 ( .A(n445), .B(n444), .ZN(n551) );
  NAND2_X1 U443 ( .A1(n440), .A2(n604), .ZN(n445) );
  XNOR2_X1 U444 ( .A(n732), .B(n408), .ZN(n427) );
  XNOR2_X1 U445 ( .A(n428), .B(n427), .ZN(n439) );
  XNOR2_X1 U446 ( .A(n439), .B(n438), .ZN(n622) );
  XNOR2_X2 U447 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n434) );
  BUF_X1 U448 ( .A(n519), .Z(n556) );
  OR2_X2 U449 ( .A1(n630), .A2(G902), .ZN(n422) );
  XNOR2_X1 U450 ( .A(n401), .B(n400), .ZN(n519) );
  XOR2_X1 U451 ( .A(n465), .B(n464), .Z(n386) );
  XOR2_X1 U452 ( .A(n448), .B(n447), .Z(n387) );
  OR2_X1 U453 ( .A1(n585), .A2(KEYINPUT47), .ZN(n388) );
  BUF_X1 U454 ( .A(n671), .Z(n713) );
  NOR2_X1 U455 ( .A1(n558), .A2(n557), .ZN(n567) );
  XNOR2_X1 U456 ( .A(n746), .B(n386), .ZN(n472) );
  XNOR2_X1 U457 ( .A(n472), .B(n471), .ZN(n617) );
  XNOR2_X1 U458 ( .A(n473), .B(n615), .ZN(n474) );
  AND2_X1 U459 ( .A1(n580), .A2(n581), .ZN(n653) );
  NOR2_X1 U460 ( .A1(n579), .A2(n578), .ZN(n610) );
  XOR2_X1 U461 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n389) );
  INV_X2 U462 ( .A(G125), .ZN(n663) );
  XOR2_X1 U463 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n391) );
  XOR2_X1 U464 ( .A(G119), .B(G110), .Z(n392) );
  NAND2_X1 U465 ( .A1(G234), .A2(n750), .ZN(n393) );
  XOR2_X1 U466 ( .A(KEYINPUT8), .B(n393), .Z(n481) );
  NAND2_X1 U467 ( .A1(G221), .A2(n481), .ZN(n394) );
  XNOR2_X1 U468 ( .A(n395), .B(n394), .ZN(n607) );
  NOR2_X1 U469 ( .A1(n607), .A2(G902), .ZN(n401) );
  XNOR2_X1 U470 ( .A(KEYINPUT15), .B(G902), .ZN(n604) );
  NAND2_X1 U471 ( .A1(n604), .A2(G234), .ZN(n397) );
  XNOR2_X1 U472 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n396) );
  XNOR2_X1 U473 ( .A(n397), .B(n396), .ZN(n402) );
  NAND2_X1 U474 ( .A1(G217), .A2(n402), .ZN(n399) );
  INV_X1 U475 ( .A(KEYINPUT25), .ZN(n398) );
  NAND2_X1 U476 ( .A1(n402), .A2(G221), .ZN(n404) );
  XNOR2_X1 U477 ( .A(KEYINPUT95), .B(KEYINPUT21), .ZN(n403) );
  XNOR2_X1 U478 ( .A(n404), .B(n403), .ZN(n555) );
  INV_X1 U479 ( .A(n555), .ZN(n685) );
  OR2_X2 U480 ( .A1(n519), .A2(n685), .ZN(n691) );
  XNOR2_X1 U481 ( .A(G137), .B(G131), .ZN(n405) );
  XNOR2_X1 U482 ( .A(n434), .B(n405), .ZN(n406) );
  XNOR2_X2 U483 ( .A(G143), .B(G128), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n745), .B(G146), .ZN(n413) );
  XNOR2_X2 U485 ( .A(KEYINPUT65), .B(G101), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n417), .B(KEYINPUT68), .ZN(n408) );
  NAND2_X1 U487 ( .A1(n750), .A2(G227), .ZN(n409) );
  XNOR2_X1 U488 ( .A(n409), .B(G140), .ZN(n410) );
  XNOR2_X1 U489 ( .A(n427), .B(n410), .ZN(n411) );
  XNOR2_X1 U490 ( .A(n413), .B(n411), .ZN(n638) );
  INV_X1 U491 ( .A(G469), .ZN(n636) );
  INV_X1 U492 ( .A(n495), .ZN(n562) );
  XNOR2_X2 U493 ( .A(n562), .B(KEYINPUT1), .ZN(n575) );
  INV_X1 U494 ( .A(n575), .ZN(n589) );
  NOR2_X1 U495 ( .A1(n691), .A2(n589), .ZN(n423) );
  INV_X1 U496 ( .A(n413), .ZN(n421) );
  XNOR2_X1 U497 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n414) );
  XNOR2_X1 U498 ( .A(n414), .B(KEYINPUT70), .ZN(n415) );
  XNOR2_X1 U499 ( .A(n426), .B(n415), .ZN(n419) );
  XNOR2_X1 U500 ( .A(KEYINPUT71), .B(n351), .ZN(n466) );
  NAND2_X1 U501 ( .A1(n466), .A2(G210), .ZN(n416) );
  XNOR2_X1 U502 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U503 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U504 ( .A(n421), .B(n420), .ZN(n630) );
  INV_X1 U505 ( .A(G472), .ZN(n628) );
  XNOR2_X2 U506 ( .A(n422), .B(n628), .ZN(n687) );
  XNOR2_X1 U507 ( .A(n687), .B(KEYINPUT6), .ZN(n569) );
  NAND2_X1 U508 ( .A1(n423), .A2(n569), .ZN(n424) );
  XNOR2_X2 U509 ( .A(n424), .B(KEYINPUT33), .ZN(n671) );
  XNOR2_X1 U510 ( .A(KEYINPUT16), .B(G122), .ZN(n425) );
  INV_X1 U511 ( .A(n731), .ZN(n428) );
  XNOR2_X1 U512 ( .A(KEYINPUT85), .B(KEYINPUT17), .ZN(n429) );
  XNOR2_X1 U513 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U514 ( .A(n432), .B(n431), .ZN(n437) );
  NAND2_X1 U515 ( .A1(n750), .A2(G224), .ZN(n433) );
  XNOR2_X1 U516 ( .A(n433), .B(KEYINPUT18), .ZN(n435) );
  XNOR2_X1 U517 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U518 ( .A(n437), .B(n436), .ZN(n438) );
  INV_X1 U519 ( .A(n622), .ZN(n440) );
  INV_X1 U520 ( .A(G902), .ZN(n486) );
  INV_X1 U521 ( .A(G237), .ZN(n441) );
  NAND2_X1 U522 ( .A1(n486), .A2(n441), .ZN(n446) );
  NAND2_X1 U523 ( .A1(n446), .A2(G210), .ZN(n443) );
  INV_X1 U524 ( .A(KEYINPUT75), .ZN(n442) );
  XNOR2_X1 U525 ( .A(n443), .B(n442), .ZN(n444) );
  INV_X1 U526 ( .A(n551), .ZN(n449) );
  NAND2_X1 U527 ( .A1(n446), .A2(G214), .ZN(n448) );
  INV_X1 U528 ( .A(KEYINPUT88), .ZN(n447) );
  NAND2_X1 U529 ( .A1(n449), .A2(n387), .ZN(n450) );
  XNOR2_X1 U530 ( .A(n450), .B(KEYINPUT19), .ZN(n580) );
  NOR2_X1 U531 ( .A1(G898), .A2(n750), .ZN(n451) );
  XOR2_X1 U532 ( .A(KEYINPUT90), .B(n451), .Z(n734) );
  NAND2_X1 U533 ( .A1(G237), .A2(G234), .ZN(n452) );
  XNOR2_X1 U534 ( .A(n452), .B(KEYINPUT14), .ZN(n455) );
  NAND2_X1 U535 ( .A1(n455), .A2(G902), .ZN(n453) );
  XOR2_X1 U536 ( .A(KEYINPUT91), .B(n453), .Z(n545) );
  NOR2_X1 U537 ( .A1(n734), .A2(n545), .ZN(n454) );
  XNOR2_X1 U538 ( .A(n454), .B(KEYINPUT92), .ZN(n457) );
  NAND2_X1 U539 ( .A1(n455), .A2(G952), .ZN(n456) );
  XOR2_X1 U540 ( .A(KEYINPUT89), .B(n456), .Z(n720) );
  NOR2_X1 U541 ( .A1(G953), .A2(n720), .ZN(n548) );
  OR2_X1 U542 ( .A1(n457), .A2(n548), .ZN(n459) );
  INV_X1 U543 ( .A(KEYINPUT93), .ZN(n458) );
  XNOR2_X1 U544 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U545 ( .A1(n580), .A2(n460), .ZN(n462) );
  INV_X1 U546 ( .A(KEYINPUT0), .ZN(n461) );
  BUF_X1 U547 ( .A(n514), .Z(n502) );
  NAND2_X1 U548 ( .A1(n671), .A2(n502), .ZN(n463) );
  XNOR2_X1 U549 ( .A(n463), .B(n353), .ZN(n491) );
  XOR2_X1 U550 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n465) );
  XNOR2_X1 U551 ( .A(G143), .B(KEYINPUT101), .ZN(n464) );
  NAND2_X1 U552 ( .A1(n466), .A2(G214), .ZN(n470) );
  XNOR2_X1 U553 ( .A(G113), .B(G122), .ZN(n468) );
  XOR2_X1 U554 ( .A(G131), .B(G104), .Z(n467) );
  XNOR2_X1 U555 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U556 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U557 ( .A1(G902), .A2(n617), .ZN(n475) );
  XNOR2_X1 U558 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n473) );
  INV_X1 U559 ( .A(G475), .ZN(n615) );
  XOR2_X1 U560 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n477) );
  XNOR2_X1 U561 ( .A(G107), .B(KEYINPUT9), .ZN(n476) );
  XNOR2_X1 U562 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U563 ( .A(n478), .B(KEYINPUT104), .Z(n480) );
  XNOR2_X1 U564 ( .A(G116), .B(G122), .ZN(n479) );
  XNOR2_X1 U565 ( .A(n480), .B(n479), .ZN(n485) );
  NAND2_X1 U566 ( .A1(G217), .A2(n481), .ZN(n482) );
  XNOR2_X1 U567 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U568 ( .A(n485), .B(n484), .ZN(n726) );
  NAND2_X1 U569 ( .A1(n726), .A2(n486), .ZN(n487) );
  INV_X1 U570 ( .A(G478), .ZN(n725) );
  XNOR2_X1 U571 ( .A(n487), .B(n725), .ZN(n511) );
  OR2_X1 U572 ( .A1(n512), .A2(n511), .ZN(n489) );
  INV_X1 U573 ( .A(KEYINPUT107), .ZN(n488) );
  XNOR2_X1 U574 ( .A(n489), .B(n488), .ZN(n577) );
  INV_X1 U575 ( .A(n577), .ZN(n490) );
  NAND2_X1 U576 ( .A1(n491), .A2(n490), .ZN(n493) );
  INV_X1 U577 ( .A(KEYINPUT35), .ZN(n492) );
  XNOR2_X2 U578 ( .A(n493), .B(n492), .ZN(n627) );
  INV_X1 U579 ( .A(KEYINPUT44), .ZN(n494) );
  OR2_X1 U580 ( .A1(n627), .A2(n494), .ZN(n510) );
  INV_X1 U581 ( .A(KEYINPUT96), .ZN(n496) );
  XNOR2_X1 U582 ( .A(n497), .B(n496), .ZN(n549) );
  INV_X1 U583 ( .A(n502), .ZN(n498) );
  OR2_X1 U584 ( .A1(n549), .A2(n498), .ZN(n499) );
  XNOR2_X1 U585 ( .A(n499), .B(KEYINPUT97), .ZN(n500) );
  NAND2_X1 U586 ( .A1(n500), .A2(n687), .ZN(n647) );
  NOR2_X1 U587 ( .A1(n691), .A2(n687), .ZN(n501) );
  AND2_X1 U588 ( .A1(n501), .A2(n575), .ZN(n698) );
  NAND2_X1 U589 ( .A1(n502), .A2(n698), .ZN(n506) );
  XOR2_X1 U590 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n504) );
  INV_X1 U591 ( .A(KEYINPUT99), .ZN(n503) );
  XNOR2_X1 U592 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U593 ( .A(n506), .B(n505), .ZN(n659) );
  NAND2_X1 U594 ( .A1(n647), .A2(n659), .ZN(n508) );
  INV_X1 U595 ( .A(n511), .ZN(n507) );
  AND2_X1 U596 ( .A1(n512), .A2(n507), .ZN(n650) );
  XNOR2_X1 U597 ( .A(KEYINPUT105), .B(n650), .ZN(n597) );
  NAND2_X1 U598 ( .A1(n597), .A2(n566), .ZN(n707) );
  NAND2_X1 U599 ( .A1(n508), .A2(n707), .ZN(n509) );
  NAND2_X1 U600 ( .A1(n510), .A2(n509), .ZN(n522) );
  NAND2_X1 U601 ( .A1(n512), .A2(n511), .ZN(n706) );
  NOR2_X1 U602 ( .A1(n706), .A2(n685), .ZN(n513) );
  INV_X1 U603 ( .A(n569), .ZN(n515) );
  NAND2_X1 U604 ( .A1(n516), .A2(n515), .ZN(n525) );
  XNOR2_X1 U605 ( .A(n525), .B(KEYINPUT80), .ZN(n517) );
  XNOR2_X1 U606 ( .A(n518), .B(KEYINPUT81), .ZN(n521) );
  XNOR2_X1 U607 ( .A(n556), .B(KEYINPUT106), .ZN(n684) );
  INV_X1 U608 ( .A(n684), .ZN(n520) );
  AND2_X2 U609 ( .A1(n521), .A2(n520), .ZN(n614) );
  NOR2_X2 U610 ( .A1(n522), .A2(n614), .ZN(n523) );
  XNOR2_X1 U611 ( .A(n523), .B(KEYINPUT82), .ZN(n539) );
  NAND2_X1 U612 ( .A1(n684), .A2(n575), .ZN(n524) );
  XNOR2_X1 U613 ( .A(n526), .B(KEYINPUT32), .ZN(n613) );
  NAND2_X1 U614 ( .A1(n556), .A2(n687), .ZN(n527) );
  OR2_X1 U615 ( .A1(n527), .A2(n575), .ZN(n528) );
  OR2_X1 U616 ( .A1(n529), .A2(n528), .ZN(n609) );
  NAND2_X1 U617 ( .A1(n613), .A2(n530), .ZN(n531) );
  INV_X1 U618 ( .A(KEYINPUT69), .ZN(n533) );
  XNOR2_X1 U619 ( .A(n531), .B(n533), .ZN(n532) );
  NAND2_X1 U620 ( .A1(n532), .A2(n494), .ZN(n537) );
  AND2_X1 U621 ( .A1(n533), .A2(KEYINPUT44), .ZN(n534) );
  AND2_X1 U622 ( .A1(n609), .A2(n534), .ZN(n535) );
  NAND2_X1 U623 ( .A1(n613), .A2(n535), .ZN(n536) );
  NAND2_X1 U624 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n539), .A2(n538), .ZN(n543) );
  XNOR2_X1 U626 ( .A(KEYINPUT79), .B(KEYINPUT45), .ZN(n541) );
  INV_X1 U627 ( .A(KEYINPUT64), .ZN(n540) );
  XNOR2_X1 U628 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X2 U629 ( .A(n543), .B(n542), .ZN(n668) );
  INV_X1 U630 ( .A(KEYINPUT2), .ZN(n544) );
  OR2_X1 U631 ( .A1(n750), .A2(n545), .ZN(n546) );
  NOR2_X1 U632 ( .A1(G900), .A2(n546), .ZN(n547) );
  NOR2_X1 U633 ( .A1(n548), .A2(n547), .ZN(n558) );
  INV_X1 U634 ( .A(n687), .ZN(n559) );
  NAND2_X1 U635 ( .A1(n559), .A2(n387), .ZN(n550) );
  XNOR2_X1 U636 ( .A(KEYINPUT39), .B(n552), .ZN(n596) );
  NOR2_X1 U637 ( .A1(n596), .A2(n566), .ZN(n553) );
  XNOR2_X1 U638 ( .A(n553), .B(KEYINPUT40), .ZN(n756) );
  NAND2_X1 U639 ( .A1(n350), .A2(n387), .ZN(n708) );
  NOR2_X1 U640 ( .A1(n706), .A2(n708), .ZN(n554) );
  XNOR2_X1 U641 ( .A(n554), .B(KEYINPUT41), .ZN(n703) );
  INV_X1 U642 ( .A(n703), .ZN(n672) );
  NAND2_X1 U643 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U644 ( .A1(n567), .A2(n559), .ZN(n561) );
  INV_X1 U645 ( .A(KEYINPUT28), .ZN(n560) );
  XNOR2_X1 U646 ( .A(n561), .B(n560), .ZN(n563) );
  AND2_X1 U647 ( .A1(n563), .A2(n562), .ZN(n581) );
  AND2_X1 U648 ( .A1(n672), .A2(n581), .ZN(n564) );
  XNOR2_X1 U649 ( .A(n564), .B(KEYINPUT42), .ZN(n755) );
  XNOR2_X1 U650 ( .A(KEYINPUT112), .B(KEYINPUT36), .ZN(n574) );
  XNOR2_X2 U651 ( .A(KEYINPUT108), .B(n566), .ZN(n656) );
  INV_X1 U652 ( .A(n567), .ZN(n568) );
  NOR2_X1 U653 ( .A1(n656), .A2(n568), .ZN(n570) );
  NAND2_X1 U654 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U655 ( .A(n571), .B(KEYINPUT109), .ZN(n572) );
  NAND2_X1 U656 ( .A1(n591), .A2(n449), .ZN(n573) );
  XOR2_X1 U657 ( .A(n574), .B(n573), .Z(n576) );
  NAND2_X1 U658 ( .A1(n576), .A2(n575), .ZN(n662) );
  INV_X1 U659 ( .A(n662), .ZN(n588) );
  OR2_X1 U660 ( .A1(n577), .A2(n593), .ZN(n578) );
  INV_X1 U661 ( .A(n610), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n707), .A2(n653), .ZN(n585) );
  NAND2_X1 U663 ( .A1(n585), .A2(KEYINPUT47), .ZN(n582) );
  NAND2_X1 U664 ( .A1(n583), .A2(n582), .ZN(n584) );
  BUF_X1 U665 ( .A(n589), .Z(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT43), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U669 ( .A(n595), .B(KEYINPUT110), .ZN(n754) );
  NOR2_X1 U670 ( .A1(n596), .A2(n597), .ZN(n665) );
  INV_X1 U671 ( .A(n665), .ZN(n598) );
  AND2_X1 U672 ( .A1(n754), .A2(n598), .ZN(n599) );
  INV_X1 U673 ( .A(KEYINPUT78), .ZN(n600) );
  XNOR2_X2 U674 ( .A(n667), .B(n600), .ZN(n666) );
  NAND2_X1 U675 ( .A1(n601), .A2(n666), .ZN(n678) );
  INV_X1 U676 ( .A(n667), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n602), .A2(n668), .ZN(n681) );
  NAND2_X1 U678 ( .A1(n681), .A2(KEYINPUT2), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n678), .A2(n603), .ZN(n606) );
  INV_X1 U680 ( .A(n604), .ZN(n605) );
  NAND2_X2 U681 ( .A1(n606), .A2(n605), .ZN(n724) );
  INV_X1 U682 ( .A(G952), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n609), .B(G110), .ZN(G12) );
  XOR2_X1 U684 ( .A(G143), .B(KEYINPUT115), .Z(n611) );
  XOR2_X1 U685 ( .A(n611), .B(n610), .Z(G45) );
  XOR2_X1 U686 ( .A(G119), .B(KEYINPUT127), .Z(n612) );
  XNOR2_X1 U687 ( .A(n613), .B(n612), .ZN(G21) );
  XOR2_X1 U688 ( .A(n614), .B(G101), .Z(G3) );
  NOR2_X1 U689 ( .A1(n724), .A2(n615), .ZN(n619) );
  XOR2_X1 U690 ( .A(KEYINPUT87), .B(KEYINPUT59), .Z(n616) );
  XNOR2_X1 U691 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X1 U693 ( .A1(n620), .A2(n730), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT60), .ZN(G60) );
  BUF_X1 U695 ( .A(n622), .Z(n626) );
  XOR2_X1 U696 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n624) );
  XNOR2_X1 U697 ( .A(KEYINPUT55), .B(KEYINPUT84), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n627), .B(G122), .ZN(G24) );
  NOR2_X1 U700 ( .A1(n724), .A2(n628), .ZN(n632) );
  XOR2_X1 U701 ( .A(KEYINPUT86), .B(KEYINPUT62), .Z(n629) );
  XNOR2_X1 U702 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n633), .A2(n730), .ZN(n635) );
  XNOR2_X1 U705 ( .A(KEYINPUT83), .B(KEYINPUT63), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(G57) );
  NOR2_X1 U707 ( .A1(n724), .A2(n636), .ZN(n640) );
  XNOR2_X1 U708 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(n641) );
  NOR2_X1 U711 ( .A1(n641), .A2(n730), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n642), .B(KEYINPUT122), .ZN(G54) );
  NOR2_X1 U713 ( .A1(n647), .A2(n656), .ZN(n644) );
  XNOR2_X1 U714 ( .A(G104), .B(KEYINPUT113), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n646) );
  XNOR2_X1 U717 ( .A(G107), .B(KEYINPUT114), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n649) );
  INV_X1 U719 ( .A(n650), .ZN(n658) );
  NOR2_X1 U720 ( .A1(n647), .A2(n658), .ZN(n648) );
  XOR2_X1 U721 ( .A(n649), .B(n648), .Z(G9) );
  XOR2_X1 U722 ( .A(G128), .B(KEYINPUT29), .Z(n652) );
  NAND2_X1 U723 ( .A1(n653), .A2(n650), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(G30) );
  INV_X1 U725 ( .A(n656), .ZN(n654) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n655), .B(G146), .ZN(G48) );
  NOR2_X1 U728 ( .A1(n656), .A2(n659), .ZN(n657) );
  XOR2_X1 U729 ( .A(G113), .B(n657), .Z(G15) );
  NOR2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U731 ( .A(KEYINPUT116), .B(n660), .Z(n661) );
  XNOR2_X1 U732 ( .A(G116), .B(n661), .ZN(G18) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U735 ( .A(G134), .B(n665), .Z(G36) );
  NAND2_X1 U736 ( .A1(n666), .A2(n667), .ZN(n670) );
  BUF_X1 U737 ( .A(n668), .Z(n669) );
  INV_X1 U738 ( .A(n669), .ZN(n736) );
  NOR2_X1 U739 ( .A1(n670), .A2(n736), .ZN(n677) );
  NAND2_X1 U740 ( .A1(n672), .A2(n713), .ZN(n675) );
  NOR2_X1 U741 ( .A1(KEYINPUT2), .A2(KEYINPUT76), .ZN(n673) );
  NOR2_X1 U742 ( .A1(G953), .A2(n673), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n679) );
  AND2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n683) );
  AND2_X1 U746 ( .A1(KEYINPUT2), .A2(KEYINPUT76), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n722) );
  NAND2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U750 ( .A(KEYINPUT49), .B(n686), .Z(n688) );
  AND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n697) );
  XOR2_X1 U752 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n692) );
  INV_X1 U753 ( .A(n692), .ZN(n689) );
  AND2_X1 U754 ( .A1(n691), .A2(n689), .ZN(n690) );
  NAND2_X1 U755 ( .A1(n690), .A2(n590), .ZN(n695) );
  NAND2_X1 U756 ( .A1(n590), .A2(n691), .ZN(n693) );
  NAND2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n700) );
  INV_X1 U760 ( .A(n698), .ZN(n699) );
  AND2_X1 U761 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U762 ( .A(KEYINPUT51), .B(n701), .Z(n702) );
  NOR2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U764 ( .A(n704), .B(KEYINPUT118), .ZN(n717) );
  NOR2_X1 U765 ( .A1(n350), .A2(n387), .ZN(n705) );
  NOR2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n712) );
  INV_X1 U767 ( .A(n707), .ZN(n709) );
  NOR2_X1 U768 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U769 ( .A(KEYINPUT119), .B(n710), .Z(n711) );
  NOR2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n715) );
  INV_X1 U771 ( .A(n713), .ZN(n714) );
  NOR2_X1 U772 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U774 ( .A(n718), .B(KEYINPUT52), .ZN(n719) );
  NOR2_X1 U775 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U778 ( .A1(n724), .A2(n725), .ZN(n728) );
  XOR2_X1 U779 ( .A(KEYINPUT123), .B(n726), .Z(n727) );
  XNOR2_X1 U780 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U781 ( .A1(n730), .A2(n729), .ZN(G63) );
  XOR2_X1 U782 ( .A(n732), .B(G101), .Z(n733) );
  XNOR2_X1 U783 ( .A(n731), .B(n733), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n735), .A2(n734), .ZN(n743) );
  NOR2_X1 U785 ( .A1(n736), .A2(G953), .ZN(n741) );
  NAND2_X1 U786 ( .A1(G953), .A2(G224), .ZN(n737) );
  XNOR2_X1 U787 ( .A(KEYINPUT61), .B(n737), .ZN(n738) );
  NAND2_X1 U788 ( .A1(n738), .A2(G898), .ZN(n739) );
  XNOR2_X1 U789 ( .A(n739), .B(KEYINPUT125), .ZN(n740) );
  NOR2_X1 U790 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U791 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U792 ( .A(KEYINPUT126), .B(n744), .ZN(G69) );
  XOR2_X1 U793 ( .A(n745), .B(n746), .Z(n749) );
  XOR2_X1 U794 ( .A(G227), .B(n749), .Z(n747) );
  NAND2_X1 U795 ( .A1(G900), .A2(n747), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(G953), .ZN(n753) );
  XNOR2_X1 U797 ( .A(n666), .B(n749), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n753), .A2(n752), .ZN(G72) );
  XNOR2_X1 U800 ( .A(G140), .B(n754), .ZN(G42) );
  XOR2_X1 U801 ( .A(G137), .B(n755), .Z(G39) );
  XOR2_X1 U802 ( .A(G131), .B(n756), .Z(G33) );
endmodule

