//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n660, new_n661, new_n664, new_n666, new_n667, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AND2_X1   g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n452), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n465), .A2(new_n467), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT70), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n471), .B(new_n477), .C1(new_n472), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n466), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n470), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n470), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n480), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(G113), .A2(G2104), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n479), .A2(new_n488), .ZN(G160));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G112), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n465), .A2(new_n470), .A3(new_n467), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n493), .B(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n496), .B2(G124), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n473), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G136), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n497), .B2(new_n501), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(G162));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(G114), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(G2105), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n473), .A2(KEYINPUT73), .A3(G114), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G126), .A2(G2105), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n493), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G138), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(G2105), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n465), .A2(new_n467), .A3(new_n516), .A4(new_n470), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT4), .ZN(new_n518));
  NOR3_X1   g093(.A1(new_n515), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n519));
  INV_X1    g094(.A(new_n485), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n484), .B1(new_n470), .B2(new_n481), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n514), .B1(new_n518), .B2(new_n522), .ZN(G164));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT76), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(G543), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT75), .B(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n526), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT75), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(new_n525), .A3(KEYINPUT5), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n524), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n537));
  NAND2_X1  g112(.A1(G75), .A2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n538), .B1(new_n536), .B2(KEYINPUT77), .ZN(new_n539));
  OAI21_X1  g114(.A(G651), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(KEYINPUT6), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT6), .ZN(new_n543));
  OAI21_X1  g118(.A(KEYINPUT74), .B1(new_n543), .B2(G651), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n545), .A2(new_n541), .A3(KEYINPUT6), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(G50), .A2(G543), .ZN(new_n548));
  OAI21_X1  g123(.A(KEYINPUT76), .B1(new_n530), .B2(KEYINPUT5), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n534), .B2(KEYINPUT5), .ZN(new_n550));
  AOI211_X1 g125(.A(KEYINPUT76), .B(new_n526), .C1(new_n531), .C2(new_n533), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G88), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n548), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n540), .A2(KEYINPUT78), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n556), .B(G651), .C1(new_n537), .C2(new_n539), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(G303));
  INV_X1    g133(.A(G303), .ZN(G166));
  INV_X1    g134(.A(new_n542), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n545), .B1(KEYINPUT6), .B2(new_n541), .ZN(new_n561));
  NOR3_X1   g136(.A1(new_n543), .A2(KEYINPUT74), .A3(G651), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT79), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n565), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n564), .A2(G51), .A3(G543), .A4(new_n566), .ZN(new_n567));
  OAI211_X1 g142(.A(G63), .B(G651), .C1(new_n550), .C2(new_n551), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT80), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n567), .A2(KEYINPUT80), .A3(new_n568), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT81), .B(KEYINPUT7), .ZN(new_n573));
  NAND3_X1  g148(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n563), .B1(new_n529), .B2(new_n535), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(G89), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(G286));
  INV_X1    g153(.A(G286), .ZN(G168));
  NAND2_X1  g154(.A1(new_n529), .A2(new_n535), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n541), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n564), .A2(G52), .A3(G543), .A4(new_n566), .ZN(new_n583));
  OAI211_X1 g158(.A(G90), .B(new_n547), .C1(new_n550), .C2(new_n551), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n583), .A2(KEYINPUT82), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT82), .B1(new_n583), .B2(new_n584), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(G301));
  INV_X1    g162(.A(G301), .ZN(G171));
  INV_X1    g163(.A(G56), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n529), .B2(new_n535), .ZN(new_n590));
  AND2_X1   g165(.A1(G68), .A2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n530), .B1(new_n563), .B2(KEYINPUT79), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT83), .B(G43), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n593), .A2(new_n566), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n576), .A2(G81), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G860), .ZN(G153));
  NAND4_X1  g173(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g174(.A1(G1), .A2(G3), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT8), .ZN(new_n601));
  NAND4_X1  g176(.A1(G319), .A2(G483), .A3(G661), .A4(new_n601), .ZN(G188));
  NAND4_X1  g177(.A1(new_n564), .A2(G53), .A3(G543), .A4(new_n566), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT9), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(KEYINPUT84), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n605), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n593), .A2(G53), .A3(new_n566), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n576), .A2(G91), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n611));
  OAI21_X1  g186(.A(G65), .B1(new_n550), .B2(new_n551), .ZN(new_n612));
  NAND2_X1  g187(.A1(G78), .A2(G543), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n611), .B1(new_n614), .B2(G651), .ZN(new_n615));
  INV_X1    g190(.A(G65), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n529), .B2(new_n535), .ZN(new_n617));
  INV_X1    g192(.A(new_n613), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n611), .B(G651), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n609), .B(new_n610), .C1(new_n615), .C2(new_n620), .ZN(G299));
  NAND4_X1  g196(.A1(new_n564), .A2(G49), .A3(G543), .A4(new_n566), .ZN(new_n622));
  INV_X1    g197(.A(G74), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n529), .A2(new_n535), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G651), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n580), .A2(G87), .A3(new_n547), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n622), .A2(new_n625), .A3(new_n626), .ZN(G288));
  AOI22_X1  g202(.A1(new_n580), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(new_n563), .ZN(new_n629));
  INV_X1    g204(.A(G61), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n529), .B2(new_n535), .ZN(new_n631));
  AND2_X1   g206(.A1(G73), .A2(G543), .ZN(new_n632));
  OAI21_X1  g207(.A(G651), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g210(.A(KEYINPUT86), .B(G651), .C1(new_n631), .C2(new_n632), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n629), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G305));
  AOI22_X1  g213(.A1(new_n580), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(new_n541), .ZN(new_n640));
  OAI21_X1  g215(.A(G543), .B1(new_n547), .B2(new_n565), .ZN(new_n641));
  INV_X1    g216(.A(new_n566), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G47), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n576), .A2(G85), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n640), .A2(new_n644), .A3(new_n645), .ZN(G290));
  NAND2_X1  g221(.A1(G301), .A2(G868), .ZN(new_n647));
  NAND2_X1  g222(.A1(G79), .A2(G543), .ZN(new_n648));
  INV_X1    g223(.A(G66), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n552), .B2(new_n649), .ZN(new_n650));
  AOI22_X1  g225(.A1(new_n650), .A2(G651), .B1(new_n643), .B2(G54), .ZN(new_n651));
  AOI21_X1  g226(.A(KEYINPUT10), .B1(new_n576), .B2(G92), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n576), .A2(G92), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n651), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n647), .B1(new_n657), .B2(G868), .ZN(G321));
  XOR2_X1   g233(.A(G321), .B(KEYINPUT87), .Z(G284));
  INV_X1    g234(.A(G868), .ZN(new_n660));
  NAND2_X1  g235(.A1(G299), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(G168), .B2(new_n660), .ZN(G297));
  OAI21_X1  g237(.A(new_n661), .B1(G168), .B2(new_n660), .ZN(G280));
  INV_X1    g238(.A(G559), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n657), .B1(new_n664), .B2(G860), .ZN(G148));
  NAND2_X1  g240(.A1(new_n657), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G868), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(G868), .B2(new_n597), .ZN(G323));
  XNOR2_X1  g243(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n669));
  XNOR2_X1  g244(.A(G323), .B(new_n669), .ZN(G282));
  NAND2_X1  g245(.A1(new_n483), .A2(new_n485), .ZN(new_n671));
  INV_X1    g246(.A(new_n474), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT12), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT13), .ZN(new_n676));
  AOI22_X1  g251(.A1(new_n675), .A2(new_n676), .B1(KEYINPUT89), .B2(G2100), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(new_n676), .B2(new_n675), .ZN(new_n678));
  NOR2_X1   g253(.A1(KEYINPUT89), .A2(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n500), .A2(G135), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n496), .A2(G123), .ZN(new_n682));
  OR2_X1    g257(.A1(G99), .A2(G2105), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n683), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G2096), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n686), .ZN(G156));
  XNOR2_X1  g262(.A(KEYINPUT15), .B(G2435), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT91), .B(G2438), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2427), .B(G2430), .Z(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n692), .A2(KEYINPUT14), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G2443), .B(G2446), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G2451), .B(G2454), .Z(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT90), .B(KEYINPUT16), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n696), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1341), .B(G1348), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT92), .Z(new_n703));
  INV_X1    g278(.A(G14), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n700), .B2(new_n701), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n703), .A2(new_n705), .ZN(G401));
  XOR2_X1   g281(.A(G2084), .B(G2090), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G2072), .A2(G2078), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n442), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G2067), .B(G2678), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n708), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT18), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n710), .A2(KEYINPUT93), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n710), .A2(KEYINPUT93), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n715), .A2(new_n716), .A3(new_n712), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n710), .B(KEYINPUT17), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n717), .B(new_n708), .C1(new_n718), .C2(new_n712), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n718), .A2(new_n712), .A3(new_n707), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n714), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(G2096), .B(G2100), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(G227));
  XOR2_X1   g298(.A(G1956), .B(G2474), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT95), .ZN(new_n725));
  XNOR2_X1  g300(.A(G1961), .B(G1966), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n728));
  XNOR2_X1  g303(.A(G1971), .B(G1976), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT20), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n725), .A2(new_n726), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n727), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n732), .B(new_n734), .C1(new_n730), .C2(new_n733), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT96), .ZN(new_n736));
  XNOR2_X1  g311(.A(G1991), .B(G1996), .ZN(new_n737));
  XNOR2_X1  g312(.A(G1981), .B(G1986), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n740));
  XOR2_X1   g315(.A(new_n739), .B(new_n740), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n735), .A2(KEYINPUT96), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n735), .A2(KEYINPUT96), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n744), .A2(new_n745), .A3(new_n741), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n746), .ZN(G229));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n748), .A2(G32), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT26), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n752), .A2(new_n753), .B1(G105), .B2(new_n672), .ZN(new_n754));
  INV_X1    g329(.A(G141), .ZN(new_n755));
  INV_X1    g330(.A(G129), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n495), .A2(G2105), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n754), .B1(new_n499), .B2(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n749), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(G160), .A2(G29), .ZN(new_n762));
  INV_X1    g337(.A(G34), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n763), .B2(KEYINPUT24), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT24), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G2084), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G16), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(G5), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G301), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT104), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n497), .A2(new_n501), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(KEYINPUT72), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n748), .B1(new_n779), .B2(new_n502), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n748), .A2(G35), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n780), .A2(KEYINPUT29), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n784));
  OAI21_X1  g359(.A(G29), .B1(new_n503), .B2(new_n504), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n781), .ZN(new_n786));
  OAI21_X1  g361(.A(G2090), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n770), .A2(G21), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G168), .B2(new_n770), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G1966), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT103), .ZN(new_n791));
  OAI21_X1  g366(.A(KEYINPUT29), .B1(new_n780), .B2(new_n782), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n785), .A2(new_n784), .A3(new_n781), .ZN(new_n793));
  INV_X1    g368(.A(G2090), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n777), .A2(new_n787), .A3(new_n791), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G27), .A2(G29), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G164), .B2(G29), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G2078), .ZN(new_n799));
  INV_X1    g374(.A(new_n685), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT31), .B(G11), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT30), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(G28), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n748), .B1(new_n803), .B2(G28), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n798), .B2(G2078), .ZN(new_n807));
  INV_X1    g382(.A(G2084), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n801), .B(new_n807), .C1(new_n808), .C2(new_n766), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n748), .A2(G33), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n671), .A2(G127), .ZN(new_n811));
  INV_X1    g386(.A(G115), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n464), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n473), .B1(new_n813), .B2(KEYINPUT102), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(KEYINPUT102), .B2(new_n813), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT25), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n500), .B2(G139), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  AOI211_X1 g394(.A(G2072), .B(new_n810), .C1(new_n819), .C2(G29), .ZN(new_n820));
  NOR2_X1   g395(.A1(G16), .A2(G19), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n597), .B2(G16), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(G1341), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n809), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n759), .A2(new_n760), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n822), .A2(G1341), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n810), .B1(new_n819), .B2(G29), .ZN(new_n827));
  INV_X1    g402(.A(G2072), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n825), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n772), .A2(new_n773), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n748), .A2(G26), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT28), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n834));
  INV_X1    g409(.A(G116), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(G2105), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n496), .B2(G128), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n500), .A2(G140), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n837), .A2(KEYINPUT101), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT101), .B1(new_n837), .B2(new_n838), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g417(.A(G2067), .B(new_n833), .C1(new_n842), .C2(new_n748), .ZN(new_n843));
  INV_X1    g418(.A(G2067), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n837), .A2(new_n838), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n748), .B1(new_n847), .B2(new_n839), .ZN(new_n848));
  INV_X1    g423(.A(new_n833), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n770), .A2(G4), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n657), .B2(new_n770), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT100), .B(G1348), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n824), .A2(new_n831), .A3(new_n851), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n769), .A2(KEYINPUT104), .A3(new_n774), .ZN(new_n857));
  NAND2_X1  g432(.A1(G299), .A2(G16), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n770), .A2(G20), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT23), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT105), .B(G1956), .Z(new_n862));
  OR2_X1    g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n789), .A2(G1966), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n862), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n857), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n796), .A2(new_n856), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n770), .A2(G23), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G288), .B2(G16), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI211_X1 g447(.A(KEYINPUT33), .B(new_n869), .C1(G288), .C2(G16), .ZN(new_n873));
  OAI21_X1  g448(.A(G1976), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n576), .A2(G87), .B1(new_n624), .B2(G651), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n770), .B1(new_n875), .B2(new_n622), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT33), .B1(new_n876), .B2(new_n869), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n870), .A2(new_n871), .ZN(new_n878));
  INV_X1    g453(.A(G1976), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n770), .A2(G6), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n637), .B2(new_n770), .ZN(new_n883));
  XNOR2_X1  g458(.A(KEYINPUT32), .B(G1981), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n881), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n555), .A2(G16), .A3(new_n557), .ZN(new_n888));
  OR2_X1    g463(.A1(G16), .A2(G22), .ZN(new_n889));
  AOI21_X1  g464(.A(G1971), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(G1971), .A3(new_n889), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n887), .A2(KEYINPUT34), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT34), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n881), .A2(new_n892), .A3(new_n885), .A4(new_n886), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G1991), .Z(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n500), .A2(G131), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n496), .A2(G119), .ZN(new_n902));
  OAI21_X1  g477(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n903));
  INV_X1    g478(.A(G107), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(G2105), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G29), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n748), .A2(G25), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT97), .Z(new_n910));
  AOI21_X1  g485(.A(new_n900), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n905), .B1(new_n496), .B2(G119), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n748), .B1(new_n912), .B2(new_n901), .ZN(new_n913));
  INV_X1    g488(.A(new_n910), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n913), .A2(KEYINPUT98), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n899), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n908), .A2(new_n900), .A3(new_n910), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT98), .B1(new_n913), .B2(new_n914), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n898), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n640), .A2(G16), .A3(new_n644), .A4(new_n645), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT99), .ZN(new_n922));
  OR2_X1    g497(.A1(G16), .A2(G24), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(G1986), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  INV_X1    g503(.A(G1986), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n924), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n920), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n868), .B1(new_n897), .B2(new_n933), .ZN(new_n934));
  AOI211_X1 g509(.A(KEYINPUT36), .B(new_n932), .C1(new_n893), .C2(new_n896), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n867), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(G311));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n936), .B(new_n938), .ZN(G150));
  NAND4_X1  g514(.A1(new_n564), .A2(G55), .A3(G543), .A4(new_n566), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n580), .A2(G93), .A3(new_n547), .ZN(new_n941));
  AND2_X1   g516(.A1(G80), .A2(G543), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n580), .B2(G67), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n940), .B(new_n941), .C1(new_n943), .C2(new_n541), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n947));
  INV_X1    g522(.A(G67), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n529), .B2(new_n535), .ZN(new_n949));
  OAI21_X1  g524(.A(G651), .B1(new_n949), .B2(new_n942), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n950), .A2(KEYINPUT107), .A3(new_n940), .A4(new_n941), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n947), .A3(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n950), .A2(new_n940), .A3(new_n941), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n597), .A2(new_n953), .A3(KEYINPUT107), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT38), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n657), .A2(G559), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n956), .B(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT39), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT108), .Z(new_n961));
  AOI21_X1  g536(.A(G860), .B1(new_n958), .B2(new_n959), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n944), .A2(G860), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT109), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT37), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n966), .ZN(G145));
  INV_X1    g542(.A(KEYINPUT40), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n500), .A2(G142), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n496), .A2(G130), .ZN(new_n970));
  OR2_X1    g545(.A1(G106), .A2(G2105), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n971), .B(G2104), .C1(G118), .C2(new_n473), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n674), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n973), .A2(new_n674), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n907), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n973), .A2(new_n674), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(new_n901), .A3(new_n912), .A4(new_n974), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n977), .B2(new_n979), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n522), .A2(new_n518), .ZN(new_n984));
  INV_X1    g559(.A(new_n514), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n840), .A2(new_n986), .A3(new_n841), .ZN(new_n987));
  AOI21_X1  g562(.A(G164), .B1(new_n847), .B2(new_n839), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n758), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(new_n840), .B2(new_n841), .ZN(new_n990));
  INV_X1    g565(.A(new_n758), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n847), .A2(G164), .A3(new_n839), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n819), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n819), .B1(new_n989), .B2(new_n993), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n983), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OR3_X1    g572(.A1(new_n503), .A2(G160), .A3(new_n504), .ZN(new_n998));
  OAI21_X1  g573(.A(G160), .B1(new_n503), .B2(new_n504), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n998), .A2(new_n800), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n800), .B1(new_n998), .B2(new_n999), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n989), .A2(new_n993), .ZN(new_n1003));
  INV_X1    g578(.A(new_n819), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n982), .A3(new_n994), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n997), .A2(new_n1002), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G37), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1002), .B1(new_n997), .B2(new_n1006), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n968), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1010), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(KEYINPUT40), .A3(new_n1008), .A4(new_n1007), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1011), .A2(new_n1013), .ZN(G395));
  NAND2_X1  g589(.A1(new_n944), .A2(new_n660), .ZN(new_n1015));
  INV_X1    g590(.A(G288), .ZN(new_n1016));
  XNOR2_X1  g591(.A(G290), .B(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(G305), .A2(new_n555), .A3(new_n557), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(G305), .B1(new_n555), .B2(new_n557), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G303), .A2(new_n637), .ZN(new_n1022));
  XNOR2_X1  g597(.A(G290), .B(G288), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n1018), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n1026));
  XNOR2_X1  g601(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n666), .B(new_n955), .ZN(new_n1028));
  INV_X1    g603(.A(new_n610), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n617), .A2(new_n618), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT85), .B1(new_n1030), .B2(new_n541), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1029), .B1(new_n1031), .B2(new_n619), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n653), .B(new_n654), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1032), .A2(new_n609), .A3(new_n1033), .A4(new_n651), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G299), .A2(new_n656), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT41), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT41), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1037), .B1(new_n1042), .B2(new_n1028), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1027), .B(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1015), .B1(new_n1044), .B2(new_n660), .ZN(G295));
  OAI21_X1  g620(.A(new_n1015), .B1(new_n1044), .B2(new_n660), .ZN(G331));
  NAND2_X1  g621(.A1(new_n583), .A2(new_n584), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT82), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n583), .A2(KEYINPUT82), .A3(new_n584), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n572), .A2(new_n577), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(new_n571), .A4(new_n582), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G301), .A2(G286), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1035), .B(new_n1034), .C1(new_n1055), .C2(new_n955), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1053), .A2(new_n1054), .B1(new_n952), .B2(new_n954), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT114), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1059));
  INV_X1    g634(.A(new_n955), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1036), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  AND2_X1   g637(.A1(G301), .A2(G286), .ZN(new_n1063));
  NOR2_X1   g638(.A1(G301), .A2(G286), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n955), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1055), .A2(new_n1067), .A3(new_n955), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1055), .B2(new_n955), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1055), .A2(new_n955), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1058), .B(new_n1066), .C1(new_n1071), .C2(new_n1041), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1025), .ZN(new_n1073));
  AOI21_X1  g648(.A(G37), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1065), .A2(KEYINPUT112), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1057), .A2(new_n1067), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1061), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1039), .B(new_n1040), .C1(new_n1070), .C2(new_n1057), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1025), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1077), .A2(new_n1025), .A3(KEYINPUT113), .A4(new_n1078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1074), .A2(new_n1083), .A3(KEYINPUT43), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1085));
  AOI21_X1  g660(.A(G37), .B1(new_n1085), .B2(new_n1073), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT43), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT44), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT44), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT43), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1074), .A2(new_n1083), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1088), .A2(new_n1093), .ZN(G397));
  INV_X1    g669(.A(KEYINPUT45), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(G164), .B2(G1384), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n479), .A2(G40), .A3(new_n488), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n842), .B(G2067), .ZN(new_n1099));
  INV_X1    g674(.A(G1996), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n758), .B(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n907), .B(new_n898), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(G290), .B(G1986), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1098), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n479), .A2(G40), .A3(new_n488), .ZN(new_n1106));
  INV_X1    g681(.A(G1384), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n986), .A2(KEYINPUT45), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1096), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(G2078), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT53), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1109), .B2(G2078), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n986), .A2(new_n1115), .A3(new_n1107), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1106), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n773), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  INV_X1    g695(.A(G1966), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1109), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1106), .A2(new_n1114), .A3(new_n1116), .A4(new_n808), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(G8), .B1(new_n1124), .B2(G286), .ZN(new_n1125));
  AOI21_X1  g700(.A(G168), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT51), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT51), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(G8), .C1(new_n1124), .C2(G286), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1120), .B1(new_n1130), .B2(KEYINPUT62), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT55), .ZN(new_n1133));
  INV_X1    g708(.A(G8), .ZN(new_n1134));
  AOI211_X1 g709(.A(new_n1133), .B(new_n1134), .C1(new_n555), .C2(new_n557), .ZN(new_n1135));
  INV_X1    g710(.A(G1971), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1109), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1106), .A2(new_n1114), .A3(new_n1116), .A4(new_n794), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1134), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1132), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G164), .A2(G1384), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1106), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1016), .A2(G1976), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(G8), .ZN(new_n1144));
  NAND2_X1  g719(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1145), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1142), .A2(new_n1143), .A3(G8), .A4(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1149));
  NAND2_X1  g724(.A1(G288), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT118), .B(G1981), .Z(new_n1152));
  OAI21_X1  g727(.A(new_n633), .B1(new_n628), .B2(new_n563), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n637), .A2(new_n1152), .B1(new_n1153), .B2(G1981), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT49), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(G8), .B(new_n1142), .C1(new_n1154), .C2(KEYINPUT49), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1151), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(KEYINPUT120), .B(new_n1151), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1140), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1132), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1135), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT116), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT116), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT115), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1138), .A2(new_n1169), .B1(new_n1109), .B2(new_n1136), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n1138), .A2(new_n1169), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1134), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1127), .A2(new_n1174), .A3(new_n1129), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1131), .A2(new_n1162), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1142), .A2(G8), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n879), .B(new_n1016), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n637), .A2(new_n1152), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT119), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1177), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1172), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1153), .A2(G1981), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT49), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1177), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI22_X1  g762(.A1(new_n1144), .A2(new_n1145), .B1(G288), .B2(new_n1149), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1187), .A2(new_n1155), .B1(new_n1188), .B2(new_n1148), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1181), .B1(new_n1183), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1110), .B2(KEYINPUT53), .ZN(new_n1192));
  NOR4_X1   g767(.A1(new_n1109), .A2(KEYINPUT126), .A3(new_n1112), .A4(G2078), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1113), .B(new_n1118), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(G171), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1111), .A2(G301), .A3(new_n1113), .A4(new_n1118), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1196), .A2(KEYINPUT54), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1195), .A2(new_n1197), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1120), .B1(new_n1194), .B2(G171), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT54), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1162), .A2(new_n1198), .A3(new_n1173), .A4(new_n1201), .ZN(new_n1202));
  XOR2_X1   g777(.A(KEYINPUT56), .B(G2072), .Z(new_n1203));
  OR2_X1    g778(.A1(new_n1109), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(KEYINPUT123), .A2(KEYINPUT57), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT57), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(G299), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1032), .A2(new_n1206), .A3(new_n1207), .A4(new_n609), .ZN(new_n1210));
  INV_X1    g785(.A(G1956), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1117), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1204), .A2(new_n1209), .A3(new_n1210), .A4(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1215), .A2(KEYINPUT124), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1204), .A2(new_n1212), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1209), .A2(new_n1210), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1216), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  NOR3_X1   g795(.A1(new_n1097), .A2(G1384), .A3(G164), .ZN(new_n1221));
  AOI22_X1  g796(.A1(new_n1117), .A2(new_n854), .B1(new_n1221), .B2(new_n844), .ZN(new_n1222));
  OR2_X1    g797(.A1(new_n1222), .A2(new_n656), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1214), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1217), .A2(new_n1215), .ZN(new_n1225));
  AOI21_X1  g800(.A(KEYINPUT61), .B1(new_n1225), .B2(new_n1213), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT60), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1222), .A2(new_n656), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1227), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1222), .A2(new_n1227), .A3(new_n657), .ZN(new_n1230));
  NAND2_X1  g805(.A1(KEYINPUT125), .A2(KEYINPUT59), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n597), .A2(new_n1231), .ZN(new_n1232));
  XOR2_X1   g807(.A(KEYINPUT58), .B(G1341), .Z(new_n1233));
  NAND2_X1  g808(.A1(new_n1142), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g809(.A1(new_n1106), .A2(new_n1096), .A3(new_n1108), .A4(new_n1100), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1232), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g811(.A1(KEYINPUT125), .A2(KEYINPUT59), .ZN(new_n1237));
  NOR2_X1   g812(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g813(.A(new_n1237), .ZN(new_n1239));
  AOI211_X1 g814(.A(new_n1239), .B(new_n1232), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1230), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  NOR3_X1   g816(.A1(new_n1226), .A2(new_n1229), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g817(.A1(new_n1220), .A2(KEYINPUT61), .A3(new_n1213), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1224), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g819(.A(new_n1176), .B(new_n1190), .C1(new_n1202), .C2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g820(.A1(new_n1124), .A2(G8), .A3(G168), .ZN(new_n1246));
  INV_X1    g821(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1162), .A2(new_n1173), .A3(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g823(.A(KEYINPUT121), .B(KEYINPUT63), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1250));
  OAI21_X1  g825(.A(new_n1189), .B1(new_n1250), .B2(new_n1172), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1251), .A2(KEYINPUT122), .ZN(new_n1252));
  INV_X1    g827(.A(KEYINPUT122), .ZN(new_n1253));
  OAI211_X1 g828(.A(new_n1189), .B(new_n1253), .C1(new_n1250), .C2(new_n1172), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g830(.A(KEYINPUT63), .ZN(new_n1256));
  NOR3_X1   g831(.A1(new_n1183), .A2(new_n1256), .A3(new_n1246), .ZN(new_n1257));
  AOI22_X1  g832(.A1(new_n1248), .A2(new_n1249), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g833(.A(new_n1105), .B1(new_n1245), .B2(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g834(.A(new_n842), .B(new_n844), .ZN(new_n1260));
  OAI21_X1  g835(.A(new_n1098), .B1(new_n1260), .B2(new_n758), .ZN(new_n1261));
  NAND2_X1  g836(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1262));
  XNOR2_X1  g837(.A(new_n1262), .B(KEYINPUT46), .ZN(new_n1263));
  NAND2_X1  g838(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g839(.A(KEYINPUT47), .ZN(new_n1265));
  NAND2_X1  g840(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g841(.A1(new_n1261), .A2(KEYINPUT47), .A3(new_n1263), .ZN(new_n1267));
  AND3_X1   g842(.A1(new_n1266), .A2(KEYINPUT127), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g843(.A(KEYINPUT127), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1269));
  INV_X1    g844(.A(new_n1098), .ZN(new_n1270));
  NOR3_X1   g845(.A1(new_n1270), .A2(G1986), .A3(G290), .ZN(new_n1271));
  XNOR2_X1  g846(.A(new_n1271), .B(KEYINPUT48), .ZN(new_n1272));
  AOI21_X1  g847(.A(new_n1272), .B1(new_n1103), .B2(new_n1098), .ZN(new_n1273));
  NOR2_X1   g848(.A1(new_n907), .A2(new_n899), .ZN(new_n1274));
  NAND3_X1  g849(.A1(new_n1099), .A2(new_n1101), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g850(.A1(new_n842), .A2(new_n844), .ZN(new_n1276));
  AOI21_X1  g851(.A(new_n1270), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  OR2_X1    g852(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1278));
  NOR3_X1   g853(.A1(new_n1268), .A2(new_n1269), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g854(.A1(new_n1259), .A2(new_n1279), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g855(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1282));
  NOR2_X1   g856(.A1(G227), .A2(new_n461), .ZN(new_n1283));
  NAND3_X1  g857(.A1(new_n743), .A2(new_n746), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g858(.A(new_n1284), .B1(new_n703), .B2(new_n705), .ZN(new_n1285));
  OAI21_X1  g859(.A(new_n1285), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1286));
  NOR2_X1   g860(.A1(new_n1282), .A2(new_n1286), .ZN(G308));
  OAI221_X1 g861(.A(new_n1285), .B1(new_n1009), .B2(new_n1010), .C1(new_n1091), .C2(new_n1092), .ZN(G225));
endmodule


