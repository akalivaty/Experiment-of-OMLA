

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596;

  XOR2_X1 U323 ( .A(n364), .B(n363), .Z(n520) );
  XOR2_X1 U324 ( .A(n420), .B(n324), .Z(n291) );
  XOR2_X1 U325 ( .A(KEYINPUT89), .B(n427), .Z(n292) );
  INV_X1 U326 ( .A(KEYINPUT93), .ZN(n368) );
  XNOR2_X1 U327 ( .A(n368), .B(KEYINPUT25), .ZN(n369) );
  XNOR2_X1 U328 ( .A(n370), .B(n369), .ZN(n371) );
  INV_X1 U329 ( .A(KEYINPUT11), .ZN(n326) );
  XNOR2_X1 U330 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U331 ( .A(n477), .B(KEYINPUT120), .ZN(n478) );
  XNOR2_X1 U332 ( .A(n329), .B(n328), .ZN(n330) );
  NAND2_X1 U333 ( .A1(n397), .A2(n396), .ZN(n486) );
  XNOR2_X1 U334 ( .A(n479), .B(n478), .ZN(n480) );
  INV_X1 U335 ( .A(G190GAT), .ZN(n481) );
  INV_X1 U336 ( .A(KEYINPUT102), .ZN(n455) );
  XNOR2_X1 U337 ( .A(KEYINPUT38), .B(n454), .ZN(n504) );
  XNOR2_X1 U338 ( .A(n481), .B(KEYINPUT58), .ZN(n482) );
  XNOR2_X1 U339 ( .A(n455), .B(G50GAT), .ZN(n456) );
  XNOR2_X1 U340 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n457), .B(n456), .ZN(G1331GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT21), .B(G218GAT), .Z(n294) );
  XNOR2_X1 U343 ( .A(KEYINPUT83), .B(G211GAT), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U345 ( .A(G197GAT), .B(n295), .Z(n350) );
  XOR2_X1 U346 ( .A(KEYINPUT24), .B(KEYINPUT82), .Z(n297) );
  XNOR2_X1 U347 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U349 ( .A(G50GAT), .B(G162GAT), .Z(n324) );
  XOR2_X1 U350 ( .A(n298), .B(n324), .Z(n305) );
  XOR2_X1 U351 ( .A(G141GAT), .B(G22GAT), .Z(n441) );
  XOR2_X1 U352 ( .A(G106GAT), .B(G78GAT), .Z(n299) );
  XOR2_X1 U353 ( .A(G148GAT), .B(n299), .Z(n421) );
  INV_X1 U354 ( .A(n421), .ZN(n300) );
  XNOR2_X1 U355 ( .A(KEYINPUT22), .B(n300), .ZN(n302) );
  NAND2_X1 U356 ( .A1(G228GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n441), .B(n303), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n350), .B(n306), .ZN(n311) );
  XOR2_X1 U361 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n308) );
  XNOR2_X1 U362 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U364 ( .A(KEYINPUT2), .B(n309), .ZN(n388) );
  INV_X1 U365 ( .A(n388), .ZN(n310) );
  XOR2_X1 U366 ( .A(n311), .B(n310), .Z(n476) );
  XOR2_X1 U367 ( .A(KEYINPUT28), .B(n476), .Z(n527) );
  XOR2_X1 U368 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n313) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G29GAT), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U371 ( .A(KEYINPUT7), .B(n314), .Z(n450) );
  XOR2_X1 U372 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n316) );
  XNOR2_X1 U373 ( .A(G134GAT), .B(G106GAT), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U375 ( .A(n450), .B(n317), .Z(n331) );
  INV_X1 U376 ( .A(KEYINPUT72), .ZN(n318) );
  NAND2_X1 U377 ( .A1(n318), .A2(G85GAT), .ZN(n321) );
  INV_X1 U378 ( .A(G85GAT), .ZN(n319) );
  NAND2_X1 U379 ( .A1(n319), .A2(KEYINPUT72), .ZN(n320) );
  NAND2_X1 U380 ( .A1(n321), .A2(n320), .ZN(n323) );
  XNOR2_X1 U381 ( .A(G99GAT), .B(G92GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n420) );
  NAND2_X1 U383 ( .A1(G232GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n291), .B(n325), .ZN(n329) );
  XOR2_X1 U385 ( .A(G36GAT), .B(G190GAT), .Z(n359) );
  XNOR2_X1 U386 ( .A(G218GAT), .B(n359), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n562) );
  XOR2_X1 U388 ( .A(n562), .B(KEYINPUT36), .Z(n592) );
  XOR2_X1 U389 ( .A(G120GAT), .B(G71GAT), .Z(n431) );
  XOR2_X1 U390 ( .A(G127GAT), .B(KEYINPUT0), .Z(n333) );
  XNOR2_X1 U391 ( .A(G113GAT), .B(G134GAT), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n389) );
  XOR2_X1 U393 ( .A(n431), .B(n389), .Z(n335) );
  XNOR2_X1 U394 ( .A(G43GAT), .B(G99GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U396 ( .A(KEYINPUT81), .B(G176GAT), .Z(n337) );
  NAND2_X1 U397 ( .A1(G227GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U399 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U400 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n341) );
  XNOR2_X1 U401 ( .A(G15GAT), .B(G190GAT), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n342), .B(KEYINPUT65), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U405 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n346) );
  XNOR2_X1 U406 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U408 ( .A(G169GAT), .B(n347), .Z(n351) );
  XOR2_X1 U409 ( .A(n348), .B(n351), .Z(n536) );
  INV_X1 U410 ( .A(n536), .ZN(n523) );
  NAND2_X1 U411 ( .A1(n476), .A2(n523), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n349), .B(KEYINPUT26), .ZN(n581) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n364) );
  INV_X1 U414 ( .A(KEYINPUT74), .ZN(n352) );
  NAND2_X1 U415 ( .A1(G64GAT), .A2(n352), .ZN(n355) );
  INV_X1 U416 ( .A(G64GAT), .ZN(n353) );
  NAND2_X1 U417 ( .A1(n353), .A2(KEYINPUT74), .ZN(n354) );
  NAND2_X1 U418 ( .A1(n355), .A2(n354), .ZN(n357) );
  XNOR2_X1 U419 ( .A(G176GAT), .B(G204GAT), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n427) );
  NAND2_X1 U421 ( .A1(G226GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n292), .B(n358), .ZN(n360) );
  XOR2_X1 U423 ( .A(n360), .B(n359), .Z(n362) );
  XNOR2_X1 U424 ( .A(G8GAT), .B(G92GAT), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n520), .B(KEYINPUT27), .ZN(n393) );
  NOR2_X1 U427 ( .A1(n581), .A2(n393), .ZN(n365) );
  XNOR2_X1 U428 ( .A(KEYINPUT91), .B(n365), .ZN(n372) );
  INV_X1 U429 ( .A(n520), .ZN(n471) );
  NAND2_X1 U430 ( .A1(n536), .A2(n471), .ZN(n366) );
  XOR2_X1 U431 ( .A(KEYINPUT92), .B(n366), .Z(n367) );
  NOR2_X1 U432 ( .A1(n476), .A2(n367), .ZN(n370) );
  NAND2_X1 U433 ( .A1(n372), .A2(n371), .ZN(n392) );
  XOR2_X1 U434 ( .A(G57GAT), .B(G148GAT), .Z(n374) );
  XNOR2_X1 U435 ( .A(G1GAT), .B(G141GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U437 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n376) );
  XNOR2_X1 U438 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U440 ( .A(n378), .B(n377), .Z(n383) );
  XOR2_X1 U441 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n380) );
  NAND2_X1 U442 ( .A1(G225GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U444 ( .A(KEYINPUT88), .B(n381), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U446 ( .A(G85GAT), .B(G162GAT), .Z(n385) );
  XNOR2_X1 U447 ( .A(G29GAT), .B(G120GAT), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U449 ( .A(n387), .B(n386), .Z(n391) );
  XOR2_X1 U450 ( .A(n389), .B(n388), .Z(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n517) );
  NAND2_X1 U452 ( .A1(n392), .A2(n517), .ZN(n397) );
  INV_X1 U453 ( .A(n527), .ZN(n534) );
  NOR2_X1 U454 ( .A1(n536), .A2(n534), .ZN(n395) );
  NOR2_X1 U455 ( .A1(n393), .A2(n517), .ZN(n394) );
  XNOR2_X1 U456 ( .A(n394), .B(KEYINPUT90), .ZN(n532) );
  NAND2_X1 U457 ( .A1(n395), .A2(n532), .ZN(n396) );
  XOR2_X1 U458 ( .A(G78GAT), .B(G71GAT), .Z(n399) );
  XNOR2_X1 U459 ( .A(G183GAT), .B(G127GAT), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U461 ( .A(G64GAT), .B(G155GAT), .Z(n401) );
  XNOR2_X1 U462 ( .A(G22GAT), .B(G211GAT), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U464 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U465 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n405) );
  NAND2_X1 U466 ( .A1(G231GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U468 ( .A(KEYINPUT15), .B(n406), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U470 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n410) );
  XNOR2_X1 U471 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U473 ( .A(n412), .B(n411), .Z(n416) );
  XNOR2_X1 U474 ( .A(G15GAT), .B(G8GAT), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n413), .B(G1GAT), .ZN(n445) );
  XNOR2_X1 U476 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n414), .B(KEYINPUT13), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n445), .B(n426), .ZN(n415) );
  XOR2_X1 U479 ( .A(n416), .B(n415), .Z(n589) );
  INV_X1 U480 ( .A(n589), .ZN(n574) );
  NAND2_X1 U481 ( .A1(n486), .A2(n574), .ZN(n417) );
  NOR2_X1 U482 ( .A1(n592), .A2(n417), .ZN(n419) );
  XNOR2_X1 U483 ( .A(KEYINPUT37), .B(KEYINPUT97), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n516) );
  XOR2_X1 U485 ( .A(n420), .B(n421), .Z(n435) );
  XOR2_X1 U486 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n423) );
  NAND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n425) );
  INV_X1 U489 ( .A(KEYINPUT71), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U493 ( .A(KEYINPUT73), .B(n430), .Z(n433) );
  XNOR2_X1 U494 ( .A(n431), .B(KEYINPUT32), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U496 ( .A(n435), .B(n434), .Z(n586) );
  INV_X1 U497 ( .A(n586), .ZN(n459) );
  XOR2_X1 U498 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n437) );
  XNOR2_X1 U499 ( .A(G197GAT), .B(KEYINPUT66), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n449) );
  XOR2_X1 U501 ( .A(G113GAT), .B(G36GAT), .Z(n439) );
  XNOR2_X1 U502 ( .A(G169GAT), .B(G50GAT), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U504 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U505 ( .A1(G229GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U507 ( .A(n444), .B(KEYINPUT68), .Z(n447) );
  XNOR2_X1 U508 ( .A(n445), .B(KEYINPUT30), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U511 ( .A(n451), .B(n450), .Z(n565) );
  INV_X1 U512 ( .A(n565), .ZN(n583) );
  NAND2_X1 U513 ( .A1(n459), .A2(n583), .ZN(n452) );
  XNOR2_X1 U514 ( .A(n452), .B(KEYINPUT75), .ZN(n487) );
  NAND2_X1 U515 ( .A1(n516), .A2(n487), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n453), .B(KEYINPUT98), .ZN(n454) );
  NOR2_X1 U517 ( .A1(n527), .A2(n504), .ZN(n457) );
  INV_X1 U518 ( .A(n562), .ZN(n545) );
  NOR2_X1 U519 ( .A1(n574), .A2(n592), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n458), .B(KEYINPUT45), .ZN(n461) );
  AND2_X1 U521 ( .A1(n459), .A2(n565), .ZN(n460) );
  AND2_X1 U522 ( .A1(n461), .A2(n460), .ZN(n462) );
  XOR2_X1 U523 ( .A(n462), .B(KEYINPUT108), .Z(n469) );
  XNOR2_X1 U524 ( .A(n586), .B(KEYINPUT41), .ZN(n567) );
  NOR2_X1 U525 ( .A1(n565), .A2(n567), .ZN(n464) );
  XNOR2_X1 U526 ( .A(KEYINPUT107), .B(KEYINPUT46), .ZN(n463) );
  XNOR2_X1 U527 ( .A(n464), .B(n463), .ZN(n466) );
  NOR2_X1 U528 ( .A1(n589), .A2(n562), .ZN(n465) );
  AND2_X1 U529 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n467), .B(KEYINPUT47), .ZN(n468) );
  NAND2_X1 U531 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT48), .ZN(n531) );
  NAND2_X1 U533 ( .A1(n531), .A2(n471), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n472), .B(KEYINPUT119), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n473), .B(KEYINPUT54), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n474), .A2(n517), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n475), .B(KEYINPUT64), .ZN(n580) );
  NOR2_X1 U538 ( .A1(n580), .A2(n476), .ZN(n479) );
  INV_X1 U539 ( .A(KEYINPUT55), .ZN(n477) );
  NAND2_X1 U540 ( .A1(n480), .A2(n536), .ZN(n573) );
  NOR2_X1 U541 ( .A1(n545), .A2(n573), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n545), .A2(n589), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  AND2_X1 U544 ( .A1(n486), .A2(n485), .ZN(n507) );
  NAND2_X1 U545 ( .A1(n487), .A2(n507), .ZN(n496) );
  NOR2_X1 U546 ( .A1(n517), .A2(n496), .ZN(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U549 ( .A(G1GAT), .B(n490), .Z(G1324GAT) );
  NOR2_X1 U550 ( .A1(n520), .A2(n496), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  NOR2_X1 U553 ( .A1(n523), .A2(n496), .ZN(n494) );
  XNOR2_X1 U554 ( .A(KEYINPUT35), .B(KEYINPUT96), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(n495), .ZN(G1326GAT) );
  NOR2_X1 U557 ( .A1(n527), .A2(n496), .ZN(n497) );
  XOR2_X1 U558 ( .A(G22GAT), .B(n497), .Z(G1327GAT) );
  NOR2_X1 U559 ( .A1(n504), .A2(n517), .ZN(n501) );
  XOR2_X1 U560 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n499) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT100), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n520), .A2(n504), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(KEYINPUT101), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(G1329GAT) );
  NOR2_X1 U567 ( .A1(n523), .A2(n504), .ZN(n505) );
  XOR2_X1 U568 ( .A(KEYINPUT40), .B(n505), .Z(n506) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NOR2_X1 U570 ( .A1(n583), .A2(n567), .ZN(n515) );
  NAND2_X1 U571 ( .A1(n515), .A2(n507), .ZN(n512) );
  NOR2_X1 U572 ( .A1(n517), .A2(n512), .ZN(n508) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n508), .Z(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n520), .A2(n512), .ZN(n510) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n523), .A2(n512), .ZN(n511) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n511), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n527), .A2(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n517), .A2(n526), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(KEYINPUT103), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NOR2_X1 U586 ( .A1(n520), .A2(n526), .ZN(n521) );
  XOR2_X1 U587 ( .A(KEYINPUT104), .B(n521), .Z(n522) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  NOR2_X1 U589 ( .A1(n523), .A2(n526), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT105), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1338GAT) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT106), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U595 ( .A(G106GAT), .B(n530), .Z(G1339GAT) );
  NAND2_X1 U596 ( .A1(n531), .A2(n532), .ZN(n533) );
  XOR2_X1 U597 ( .A(KEYINPUT109), .B(n533), .Z(n551) );
  NOR2_X1 U598 ( .A1(n534), .A2(n551), .ZN(n535) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n546) );
  NOR2_X1 U600 ( .A1(n565), .A2(n546), .ZN(n538) );
  XNOR2_X1 U601 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n539), .ZN(G1340GAT) );
  NOR2_X1 U604 ( .A1(n567), .A2(n546), .ZN(n541) );
  XNOR2_X1 U605 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n542), .ZN(G1341GAT) );
  NOR2_X1 U608 ( .A1(n574), .A2(n546), .ZN(n543) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(n543), .Z(n544) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n548) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT115), .Z(n553) );
  NOR2_X1 U617 ( .A1(n581), .A2(n551), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n561), .A2(n583), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XNOR2_X1 U620 ( .A(KEYINPUT116), .B(KEYINPUT52), .ZN(n558) );
  XOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .Z(n556) );
  INV_X1 U622 ( .A(n567), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n561), .A2(n554), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  XOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT117), .Z(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n589), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT118), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n573), .ZN(n566) );
  XOR2_X1 U633 ( .A(G169GAT), .B(n566), .Z(G1348GAT) );
  NOR2_X1 U634 ( .A1(n573), .A2(n567), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(KEYINPUT56), .B(n570), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1350GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT125), .B(n579), .Z(n585) );
  NOR2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U648 ( .A(n582), .B(KEYINPUT124), .Z(n593) );
  INV_X1 U649 ( .A(n593), .ZN(n590) );
  NAND2_X1 U650 ( .A1(n583), .A2(n590), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U652 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  NAND2_X1 U653 ( .A1(n586), .A2(n590), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n591), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U658 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

