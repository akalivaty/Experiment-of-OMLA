

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U319 ( .A(n388), .B(KEYINPUT48), .ZN(n543) );
  AND2_X1 U320 ( .A1(n387), .A2(n386), .ZN(n388) );
  INV_X1 U321 ( .A(KEYINPUT37), .ZN(n470) );
  XOR2_X1 U322 ( .A(n364), .B(n335), .Z(n287) );
  XOR2_X1 U323 ( .A(n369), .B(n368), .Z(n288) );
  XOR2_X1 U324 ( .A(n321), .B(n320), .Z(n289) );
  XOR2_X1 U325 ( .A(G64GAT), .B(KEYINPUT71), .Z(n290) );
  XOR2_X1 U326 ( .A(n364), .B(n437), .Z(n291) );
  INV_X1 U327 ( .A(G134GAT), .ZN(n294) );
  XNOR2_X1 U328 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U329 ( .A(n297), .B(n296), .ZN(n298) );
  INV_X1 U330 ( .A(KEYINPUT99), .ZN(n454) );
  XNOR2_X1 U331 ( .A(n322), .B(n289), .ZN(n323) );
  XNOR2_X1 U332 ( .A(n455), .B(n454), .ZN(n542) );
  XNOR2_X1 U333 ( .A(n324), .B(n323), .ZN(n328) );
  NOR2_X1 U334 ( .A1(n415), .A2(n515), .ZN(n561) );
  XNOR2_X1 U335 ( .A(n471), .B(n470), .ZN(n514) );
  XOR2_X1 U336 ( .A(n373), .B(n372), .Z(n568) );
  NOR2_X1 U337 ( .A1(n450), .A2(n527), .ZN(n557) );
  XOR2_X1 U338 ( .A(n449), .B(n448), .Z(n521) );
  XNOR2_X1 U339 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n451) );
  XNOR2_X1 U340 ( .A(n474), .B(G43GAT), .ZN(n475) );
  XNOR2_X1 U341 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n476), .B(n475), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n293) );
  XNOR2_X1 U344 ( .A(KEYINPUT73), .B(KEYINPUT78), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n297) );
  NAND2_X1 U346 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U347 ( .A(n298), .B(KEYINPUT9), .Z(n305) );
  XOR2_X1 U348 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n302) );
  XOR2_X1 U349 ( .A(G50GAT), .B(G162GAT), .Z(n417) );
  XOR2_X1 U350 ( .A(KEYINPUT77), .B(G218GAT), .Z(n300) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n319) );
  XNOR2_X1 U353 ( .A(n417), .B(n319), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n303), .B(KEYINPUT75), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n314) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(KEYINPUT68), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n306), .B(G29GAT), .ZN(n307) );
  XOR2_X1 U359 ( .A(n307), .B(KEYINPUT67), .Z(n309) );
  XNOR2_X1 U360 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n359) );
  XOR2_X1 U362 ( .A(KEYINPUT70), .B(G92GAT), .Z(n311) );
  XNOR2_X1 U363 ( .A(G99GAT), .B(G85GAT), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U365 ( .A(G106GAT), .B(n312), .Z(n373) );
  XNOR2_X1 U366 ( .A(n359), .B(n373), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n376) );
  XNOR2_X1 U368 ( .A(KEYINPUT79), .B(n376), .ZN(n538) );
  XNOR2_X1 U369 ( .A(G176GAT), .B(G204GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n290), .B(n315), .ZN(n364) );
  XOR2_X1 U371 ( .A(G8GAT), .B(G183GAT), .Z(n335) );
  NAND2_X1 U372 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n287), .B(n316), .ZN(n324) );
  XOR2_X1 U374 ( .A(G211GAT), .B(KEYINPUT21), .Z(n318) );
  XNOR2_X1 U375 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n418) );
  XNOR2_X1 U377 ( .A(n418), .B(n319), .ZN(n322) );
  XOR2_X1 U378 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n321) );
  XNOR2_X1 U379 ( .A(G92GAT), .B(KEYINPUT98), .ZN(n320) );
  XOR2_X1 U380 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n326) );
  XNOR2_X1 U381 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U383 ( .A(G169GAT), .B(n327), .Z(n449) );
  XOR2_X1 U384 ( .A(n328), .B(n449), .Z(n453) );
  XOR2_X1 U385 ( .A(KEYINPUT47), .B(KEYINPUT116), .Z(n379) );
  XOR2_X1 U386 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n330) );
  XNOR2_X1 U387 ( .A(G64GAT), .B(KEYINPUT83), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U389 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n332) );
  XNOR2_X1 U390 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n346) );
  XOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT13), .Z(n370) );
  XOR2_X1 U394 ( .A(n370), .B(n335), .Z(n337) );
  XNOR2_X1 U395 ( .A(G78GAT), .B(G211GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U397 ( .A(G22GAT), .B(G155GAT), .Z(n420) );
  XNOR2_X1 U398 ( .A(G15GAT), .B(G1GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n338), .B(KEYINPUT69), .ZN(n355) );
  XOR2_X1 U400 ( .A(n420), .B(n355), .Z(n340) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U403 ( .A(n342), .B(n341), .Z(n344) );
  XNOR2_X1 U404 ( .A(G127GAT), .B(G71GAT), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U406 ( .A(n346), .B(n345), .Z(n573) );
  INV_X1 U407 ( .A(n573), .ZN(n556) );
  XOR2_X1 U408 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n348) );
  XNOR2_X1 U409 ( .A(KEYINPUT64), .B(KEYINPUT30), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n363) );
  XOR2_X1 U411 ( .A(G113GAT), .B(G50GAT), .Z(n350) );
  XNOR2_X1 U412 ( .A(G169GAT), .B(G36GAT), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U414 ( .A(G8GAT), .B(G197GAT), .Z(n352) );
  XNOR2_X1 U415 ( .A(G141GAT), .B(G22GAT), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U417 ( .A(n354), .B(n353), .Z(n361) );
  XOR2_X1 U418 ( .A(n355), .B(KEYINPUT66), .Z(n357) );
  NAND2_X1 U419 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n554) );
  INV_X1 U424 ( .A(n554), .ZN(n562) );
  XOR2_X1 U425 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n291), .B(n365), .ZN(n369) );
  XOR2_X1 U428 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n367) );
  XNOR2_X1 U429 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U431 ( .A(G148GAT), .B(G78GAT), .Z(n416) );
  XNOR2_X1 U432 ( .A(n416), .B(n370), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n288), .B(n371), .ZN(n372) );
  XOR2_X1 U434 ( .A(KEYINPUT41), .B(n568), .Z(n546) );
  NOR2_X1 U435 ( .A1(n562), .A2(n546), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n374), .B(KEYINPUT46), .ZN(n375) );
  NOR2_X1 U437 ( .A1(n556), .A2(n375), .ZN(n377) );
  NAND2_X1 U438 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n387) );
  INV_X1 U440 ( .A(n568), .ZN(n383) );
  XNOR2_X1 U441 ( .A(KEYINPUT45), .B(KEYINPUT117), .ZN(n381) );
  XNOR2_X1 U442 ( .A(KEYINPUT36), .B(n538), .ZN(n576) );
  NAND2_X1 U443 ( .A1(n576), .A2(n556), .ZN(n380) );
  XOR2_X1 U444 ( .A(n381), .B(n380), .Z(n382) );
  NOR2_X1 U445 ( .A1(n383), .A2(n382), .ZN(n384) );
  XNOR2_X1 U446 ( .A(KEYINPUT118), .B(n384), .ZN(n385) );
  NAND2_X1 U447 ( .A1(n385), .A2(n562), .ZN(n386) );
  NOR2_X1 U448 ( .A1(n453), .A2(n543), .ZN(n390) );
  INV_X1 U449 ( .A(KEYINPUT54), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n415) );
  XOR2_X1 U451 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n392) );
  XNOR2_X1 U452 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U454 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n394) );
  XNOR2_X1 U455 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U457 ( .A(n396), .B(n395), .Z(n406) );
  XNOR2_X1 U458 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n397), .B(KEYINPUT85), .ZN(n398) );
  XOR2_X1 U460 ( .A(n398), .B(KEYINPUT84), .Z(n400) );
  XNOR2_X1 U461 ( .A(G113GAT), .B(G134GAT), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n445) );
  XNOR2_X1 U463 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n401), .B(KEYINPUT2), .ZN(n426) );
  XOR2_X1 U465 ( .A(n426), .B(KEYINPUT94), .Z(n403) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U468 ( .A(n445), .B(n404), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n414) );
  XOR2_X1 U470 ( .A(G57GAT), .B(G148GAT), .Z(n408) );
  XNOR2_X1 U471 ( .A(G1GAT), .B(G155GAT), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U473 ( .A(G85GAT), .B(G162GAT), .Z(n410) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(G120GAT), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U476 ( .A(n412), .B(n411), .Z(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n515) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U480 ( .A(n421), .B(n420), .Z(n423) );
  XNOR2_X1 U481 ( .A(G218GAT), .B(G106GAT), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n432) );
  XOR2_X1 U483 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n425) );
  XNOR2_X1 U484 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n430) );
  XOR2_X1 U486 ( .A(n426), .B(KEYINPUT24), .Z(n428) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U489 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n460) );
  NAND2_X1 U491 ( .A1(n561), .A2(n460), .ZN(n434) );
  XOR2_X1 U492 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n450) );
  XOR2_X1 U494 ( .A(G176GAT), .B(G183GAT), .Z(n436) );
  XNOR2_X1 U495 ( .A(G190GAT), .B(G99GAT), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U497 ( .A(n438), .B(n437), .Z(n440) );
  XNOR2_X1 U498 ( .A(G43GAT), .B(G15GAT), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U500 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n442) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n447) );
  XNOR2_X1 U504 ( .A(n445), .B(KEYINPUT20), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  INV_X1 U506 ( .A(n521), .ZN(n527) );
  NAND2_X1 U507 ( .A1(n538), .A2(n557), .ZN(n452) );
  NAND2_X1 U508 ( .A1(n554), .A2(n568), .ZN(n484) );
  INV_X1 U509 ( .A(n453), .ZN(n518) );
  XNOR2_X1 U510 ( .A(n518), .B(KEYINPUT27), .ZN(n462) );
  NAND2_X1 U511 ( .A1(n462), .A2(n515), .ZN(n455) );
  XOR2_X1 U512 ( .A(KEYINPUT28), .B(n460), .Z(n524) );
  NOR2_X1 U513 ( .A1(n542), .A2(n524), .ZN(n529) );
  INV_X1 U514 ( .A(KEYINPUT100), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n529), .B(n456), .ZN(n457) );
  NOR2_X1 U516 ( .A1(n521), .A2(n457), .ZN(n468) );
  NAND2_X1 U517 ( .A1(n521), .A2(n518), .ZN(n458) );
  NAND2_X1 U518 ( .A1(n460), .A2(n458), .ZN(n459) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n459), .Z(n464) );
  NOR2_X1 U520 ( .A1(n460), .A2(n521), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n461), .B(KEYINPUT26), .ZN(n560) );
  NAND2_X1 U522 ( .A1(n462), .A2(n560), .ZN(n463) );
  NAND2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U524 ( .A(KEYINPUT101), .B(n465), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n515), .A2(n466), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n482) );
  NOR2_X1 U527 ( .A1(n556), .A2(n482), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n469), .A2(n576), .ZN(n471) );
  OR2_X1 U529 ( .A1(n484), .A2(n514), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT38), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n473), .B(KEYINPUT107), .ZN(n500) );
  NAND2_X1 U532 ( .A1(n521), .A2(n500), .ZN(n476) );
  XOR2_X1 U533 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n474) );
  XOR2_X1 U534 ( .A(n546), .B(KEYINPUT110), .Z(n532) );
  NAND2_X1 U535 ( .A1(n532), .A2(n557), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(G176GAT), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(G1349GAT) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n486) );
  NOR2_X1 U540 ( .A1(n538), .A2(n573), .ZN(n480) );
  XOR2_X1 U541 ( .A(KEYINPUT16), .B(n480), .Z(n481) );
  NOR2_X1 U542 ( .A1(n482), .A2(n481), .ZN(n483) );
  XOR2_X1 U543 ( .A(KEYINPUT102), .B(n483), .Z(n502) );
  NOR2_X1 U544 ( .A1(n502), .A2(n484), .ZN(n492) );
  NAND2_X1 U545 ( .A1(n492), .A2(n515), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1324GAT) );
  XOR2_X1 U547 ( .A(G8GAT), .B(KEYINPUT103), .Z(n488) );
  NAND2_X1 U548 ( .A1(n492), .A2(n518), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT35), .B(KEYINPUT104), .Z(n490) );
  NAND2_X1 U551 ( .A1(n492), .A2(n521), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U553 ( .A(G15GAT), .B(n491), .ZN(G1326GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n494) );
  NAND2_X1 U555 ( .A1(n492), .A2(n524), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n495), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT108), .B(KEYINPUT39), .Z(n497) );
  NAND2_X1 U559 ( .A1(n500), .A2(n515), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U562 ( .A1(n500), .A2(n518), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U564 ( .A1(n500), .A2(n524), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n504) );
  NAND2_X1 U567 ( .A1(n562), .A2(n532), .ZN(n513) );
  NOR2_X1 U568 ( .A1(n502), .A2(n513), .ZN(n509) );
  NAND2_X1 U569 ( .A1(n509), .A2(n515), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n518), .A2(n509), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n509), .A2(n521), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n507), .B(KEYINPUT112), .ZN(n508) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U578 ( .A1(n509), .A2(n524), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U580 ( .A(G78GAT), .B(n512), .Z(G1335GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n523), .A2(n515), .ZN(n516) );
  XNOR2_X1 U583 ( .A(KEYINPUT114), .B(n516), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT115), .Z(n520) );
  NAND2_X1 U586 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n521), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n543), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(KEYINPUT119), .B(n530), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n554), .A2(n539), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U599 ( .A1(n539), .A2(n532), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n536) );
  NAND2_X1 U602 ( .A1(n539), .A2(n556), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U604 ( .A(G127GAT), .B(n537), .Z(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n544), .A2(n560), .ZN(n552) );
  NOR2_X1 U610 ( .A1(n562), .A2(n552), .ZN(n545) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n546), .A2(n552), .ZN(n548) );
  XNOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n573), .A2(n552), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n376), .A2(n552), .ZN(n553) );
  XOR2_X1 U620 ( .A(G162GAT), .B(n553), .Z(G1347GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n557), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(G183GAT), .B(KEYINPUT123), .Z(n559) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1350GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n575) );
  NOR2_X1 U627 ( .A1(n562), .A2(n575), .ZN(n567) );
  XOR2_X1 U628 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n564) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT124), .B(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  NOR2_X1 U633 ( .A1(n575), .A2(n568), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n570) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n575), .ZN(n574) );
  XOR2_X1 U639 ( .A(G211GAT), .B(n574), .Z(G1354GAT) );
  INV_X1 U640 ( .A(n575), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

