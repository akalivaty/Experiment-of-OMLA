

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(n647), .B(KEYINPUT102), .ZN(n670) );
  AND2_X1 U552 ( .A1(n969), .A2(n750), .ZN(n517) );
  NOR2_X1 U553 ( .A1(n627), .A2(n972), .ZN(n628) );
  INV_X1 U554 ( .A(n613), .ZN(n641) );
  BUF_X1 U555 ( .A(n613), .Z(n657) );
  OR2_X1 U556 ( .A1(n756), .A2(n595), .ZN(n596) );
  XNOR2_X1 U557 ( .A(G543), .B(KEYINPUT0), .ZN(n518) );
  XNOR2_X1 U558 ( .A(G2104), .B(KEYINPUT65), .ZN(n536) );
  OR2_X1 U559 ( .A1(n734), .A2(n517), .ZN(n735) );
  XNOR2_X1 U560 ( .A(n518), .B(KEYINPUT67), .ZN(n567) );
  NOR2_X2 U561 ( .A1(G2105), .A2(n536), .ZN(n876) );
  OR2_X1 U562 ( .A1(n736), .A2(n735), .ZN(n753) );
  XOR2_X1 U563 ( .A(KEYINPUT15), .B(n609), .Z(n967) );
  NOR2_X1 U564 ( .A1(G651), .A2(n567), .ZN(n785) );
  INV_X1 U565 ( .A(G651), .ZN(n525) );
  OR2_X1 U566 ( .A1(n525), .A2(n567), .ZN(n519) );
  XOR2_X2 U567 ( .A(KEYINPUT68), .B(n519), .Z(n789) );
  NAND2_X1 U568 ( .A1(G78), .A2(n789), .ZN(n522) );
  NOR2_X1 U569 ( .A1(G543), .A2(G651), .ZN(n520) );
  XNOR2_X1 U570 ( .A(n520), .B(KEYINPUT64), .ZN(n786) );
  NAND2_X1 U571 ( .A1(G91), .A2(n786), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U573 ( .A(KEYINPUT72), .B(n523), .Z(n531) );
  NAND2_X1 U574 ( .A1(n785), .A2(G53), .ZN(n524) );
  XOR2_X1 U575 ( .A(KEYINPUT73), .B(n524), .Z(n528) );
  NOR2_X1 U576 ( .A1(G543), .A2(n525), .ZN(n526) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n526), .Z(n783) );
  NAND2_X1 U578 ( .A1(n783), .A2(G65), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT74), .B(n529), .Z(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(G299) );
  AND2_X1 U582 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U583 ( .A1(G114), .A2(n879), .ZN(n534) );
  NOR2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  XOR2_X2 U585 ( .A(KEYINPUT17), .B(n532), .Z(n875) );
  NAND2_X1 U586 ( .A1(G138), .A2(n875), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U588 ( .A1(G102), .A2(n876), .ZN(n535) );
  XNOR2_X1 U589 ( .A(n535), .B(KEYINPUT90), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n536), .A2(G2105), .ZN(n537) );
  XOR2_X2 U591 ( .A(KEYINPUT66), .B(n537), .Z(n880) );
  NAND2_X1 U592 ( .A1(G126), .A2(n880), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U594 ( .A1(n541), .A2(n540), .ZN(G164) );
  NAND2_X1 U595 ( .A1(G52), .A2(n785), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G64), .A2(n783), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n549) );
  NAND2_X1 U598 ( .A1(G77), .A2(n789), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G90), .A2(n786), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  XNOR2_X1 U602 ( .A(KEYINPUT70), .B(n547), .ZN(n548) );
  NOR2_X1 U603 ( .A1(n549), .A2(n548), .ZN(G171) );
  NAND2_X1 U604 ( .A1(G89), .A2(n786), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U606 ( .A1(G76), .A2(n789), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U608 ( .A(n553), .B(KEYINPUT5), .ZN(n558) );
  NAND2_X1 U609 ( .A1(G51), .A2(n785), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G63), .A2(n783), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U614 ( .A(n559), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U615 ( .A1(G75), .A2(n789), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G88), .A2(n786), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U618 ( .A1(G62), .A2(n783), .ZN(n562) );
  XNOR2_X1 U619 ( .A(KEYINPUT87), .B(n562), .ZN(n563) );
  NOR2_X1 U620 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n785), .A2(G50), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n566), .A2(n565), .ZN(G303) );
  INV_X1 U623 ( .A(G303), .ZN(G166) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G87), .A2(n567), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G74), .A2(G651), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U628 ( .A1(n783), .A2(n570), .ZN(n573) );
  NAND2_X1 U629 ( .A1(G49), .A2(n785), .ZN(n571) );
  XOR2_X1 U630 ( .A(KEYINPUT85), .B(n571), .Z(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(G288) );
  NAND2_X1 U632 ( .A1(G61), .A2(n783), .ZN(n580) );
  NAND2_X1 U633 ( .A1(n785), .A2(G48), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G86), .A2(n786), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n789), .A2(G73), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT2), .B(n576), .Z(n577) );
  NOR2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U640 ( .A(n581), .B(KEYINPUT86), .ZN(G305) );
  NAND2_X1 U641 ( .A1(n785), .A2(G47), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G85), .A2(n786), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U644 ( .A1(G72), .A2(n789), .ZN(n584) );
  XNOR2_X1 U645 ( .A(KEYINPUT69), .B(n584), .ZN(n585) );
  NOR2_X1 U646 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n783), .A2(G60), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n588), .A2(n587), .ZN(G290) );
  NAND2_X1 U649 ( .A1(G125), .A2(n880), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G101), .A2(n876), .ZN(n589) );
  XOR2_X1 U651 ( .A(KEYINPUT23), .B(n589), .Z(n590) );
  NAND2_X1 U652 ( .A1(n591), .A2(n590), .ZN(n756) );
  INV_X1 U653 ( .A(G40), .ZN(n594) );
  NAND2_X1 U654 ( .A1(n875), .A2(G137), .ZN(n593) );
  NAND2_X1 U655 ( .A1(n879), .A2(G113), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n593), .A2(n592), .ZN(n755) );
  OR2_X1 U657 ( .A1(n594), .A2(n755), .ZN(n595) );
  XNOR2_X1 U658 ( .A(n596), .B(KEYINPUT92), .ZN(n704) );
  XNOR2_X1 U659 ( .A(n704), .B(KEYINPUT95), .ZN(n597) );
  NOR2_X1 U660 ( .A1(G164), .A2(G1384), .ZN(n703) );
  NAND2_X2 U661 ( .A1(n597), .A2(n703), .ZN(n613) );
  NAND2_X1 U662 ( .A1(n641), .A2(G2072), .ZN(n598) );
  XOR2_X1 U663 ( .A(KEYINPUT27), .B(n598), .Z(n600) );
  NAND2_X1 U664 ( .A1(G1956), .A2(n657), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n636) );
  NOR2_X1 U666 ( .A1(G299), .A2(n636), .ZN(n601) );
  XOR2_X1 U667 ( .A(KEYINPUT101), .B(n601), .Z(n635) );
  NAND2_X1 U668 ( .A1(n783), .A2(G66), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G92), .A2(n786), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n603), .A2(n602), .ZN(n608) );
  NAND2_X1 U671 ( .A1(n785), .A2(G54), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G79), .A2(n789), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U674 ( .A(KEYINPUT79), .B(n606), .Z(n607) );
  NOR2_X1 U675 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U676 ( .A1(G2067), .A2(n641), .ZN(n611) );
  NAND2_X1 U677 ( .A1(G1348), .A2(n613), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U679 ( .A(n612), .B(KEYINPUT99), .ZN(n630) );
  OR2_X1 U680 ( .A1(n967), .A2(n630), .ZN(n629) );
  INV_X1 U681 ( .A(G1996), .ZN(n944) );
  NOR2_X1 U682 ( .A1(n613), .A2(n944), .ZN(n614) );
  XOR2_X1 U683 ( .A(n614), .B(KEYINPUT26), .Z(n616) );
  NAND2_X1 U684 ( .A1(n657), .A2(G1341), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n616), .A2(n615), .ZN(n627) );
  NAND2_X1 U686 ( .A1(G81), .A2(n786), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n617), .B(KEYINPUT12), .ZN(n619) );
  NAND2_X1 U688 ( .A1(G68), .A2(n789), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n620), .B(KEYINPUT13), .ZN(n622) );
  NAND2_X1 U691 ( .A1(G43), .A2(n785), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U693 ( .A1(n783), .A2(G56), .ZN(n623) );
  XOR2_X1 U694 ( .A(KEYINPUT14), .B(n623), .Z(n624) );
  NOR2_X1 U695 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U696 ( .A(KEYINPUT75), .B(n626), .ZN(n972) );
  NAND2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U698 ( .A1(n630), .A2(n967), .ZN(n631) );
  NAND2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U700 ( .A(n633), .B(KEYINPUT100), .ZN(n634) );
  NOR2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U702 ( .A1(G299), .A2(n636), .ZN(n637) );
  XOR2_X1 U703 ( .A(KEYINPUT28), .B(n637), .Z(n638) );
  NOR2_X1 U704 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U705 ( .A(n640), .B(KEYINPUT29), .ZN(n646) );
  NOR2_X1 U706 ( .A1(n641), .A2(G1961), .ZN(n642) );
  XOR2_X1 U707 ( .A(KEYINPUT98), .B(n642), .Z(n644) );
  XNOR2_X1 U708 ( .A(G2078), .B(KEYINPUT25), .ZN(n949) );
  NAND2_X1 U709 ( .A1(n641), .A2(n949), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U711 ( .A1(n648), .A2(G171), .ZN(n645) );
  NAND2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U713 ( .A1(G171), .A2(n648), .ZN(n654) );
  NAND2_X1 U714 ( .A1(G8), .A2(n657), .ZN(n649) );
  XNOR2_X1 U715 ( .A(KEYINPUT96), .B(n649), .ZN(n683) );
  NOR2_X1 U716 ( .A1(n683), .A2(G1966), .ZN(n675) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n657), .ZN(n671) );
  NOR2_X1 U718 ( .A1(n675), .A2(n671), .ZN(n650) );
  NAND2_X1 U719 ( .A1(G8), .A2(n650), .ZN(n651) );
  XNOR2_X1 U720 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  NOR2_X1 U721 ( .A1(G168), .A2(n652), .ZN(n653) );
  NOR2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U723 ( .A(KEYINPUT31), .B(n655), .Z(n669) );
  NOR2_X1 U724 ( .A1(n683), .A2(G1971), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT103), .B(n656), .ZN(n660) );
  NOR2_X1 U726 ( .A1(G2090), .A2(n657), .ZN(n658) );
  NOR2_X1 U727 ( .A1(G166), .A2(n658), .ZN(n659) );
  NAND2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n662) );
  AND2_X1 U729 ( .A1(n669), .A2(n662), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n670), .A2(n661), .ZN(n665) );
  INV_X1 U731 ( .A(n662), .ZN(n663) );
  OR2_X1 U732 ( .A1(n663), .A2(G286), .ZN(n664) );
  AND2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n666), .A2(G8), .ZN(n668) );
  XOR2_X1 U735 ( .A(KEYINPUT32), .B(KEYINPUT104), .Z(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(n677) );
  NAND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n673) );
  NAND2_X1 U738 ( .A1(G8), .A2(n671), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X2 U741 ( .A1(n677), .A2(n676), .ZN(n698) );
  INV_X1 U742 ( .A(n698), .ZN(n681) );
  NOR2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n682) );
  NOR2_X1 U744 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n682), .A2(n678), .ZN(n976) );
  INV_X1 U746 ( .A(KEYINPUT33), .ZN(n679) );
  AND2_X1 U747 ( .A1(n976), .A2(n679), .ZN(n680) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n690) );
  AND2_X1 U749 ( .A1(n682), .A2(KEYINPUT33), .ZN(n684) );
  INV_X1 U750 ( .A(n683), .ZN(n699) );
  NAND2_X1 U751 ( .A1(n684), .A2(n699), .ZN(n688) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n980) );
  AND2_X1 U753 ( .A1(n699), .A2(n980), .ZN(n685) );
  NOR2_X1 U754 ( .A1(KEYINPUT33), .A2(n685), .ZN(n686) );
  XNOR2_X1 U755 ( .A(G1981), .B(G305), .ZN(n986) );
  NOR2_X1 U756 ( .A1(n686), .A2(n986), .ZN(n687) );
  AND2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n695) );
  NOR2_X1 U759 ( .A1(G1981), .A2(G305), .ZN(n691) );
  XOR2_X1 U760 ( .A(n691), .B(KEYINPUT24), .Z(n692) );
  XNOR2_X1 U761 ( .A(KEYINPUT97), .B(n692), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n693), .A2(n699), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n702) );
  NAND2_X1 U764 ( .A1(G166), .A2(G8), .ZN(n696) );
  NOR2_X1 U765 ( .A1(G2090), .A2(n696), .ZN(n697) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n700) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n736) );
  NOR2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n750) );
  NAND2_X1 U770 ( .A1(G140), .A2(n875), .ZN(n706) );
  NAND2_X1 U771 ( .A1(G104), .A2(n876), .ZN(n705) );
  NAND2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U773 ( .A(KEYINPUT34), .B(n707), .ZN(n713) );
  NAND2_X1 U774 ( .A1(G116), .A2(n879), .ZN(n709) );
  NAND2_X1 U775 ( .A1(G128), .A2(n880), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U777 ( .A(KEYINPUT35), .B(n710), .ZN(n711) );
  XNOR2_X1 U778 ( .A(KEYINPUT93), .B(n711), .ZN(n712) );
  NOR2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U780 ( .A(KEYINPUT36), .B(n714), .Z(n889) );
  XOR2_X1 U781 ( .A(G2067), .B(KEYINPUT37), .Z(n746) );
  AND2_X1 U782 ( .A1(n889), .A2(n746), .ZN(n921) );
  NAND2_X1 U783 ( .A1(n750), .A2(n921), .ZN(n744) );
  NAND2_X1 U784 ( .A1(G131), .A2(n875), .ZN(n716) );
  NAND2_X1 U785 ( .A1(G95), .A2(n876), .ZN(n715) );
  NAND2_X1 U786 ( .A1(n716), .A2(n715), .ZN(n720) );
  NAND2_X1 U787 ( .A1(G107), .A2(n879), .ZN(n718) );
  NAND2_X1 U788 ( .A1(G119), .A2(n880), .ZN(n717) );
  NAND2_X1 U789 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n868) );
  INV_X1 U791 ( .A(G1991), .ZN(n942) );
  NOR2_X1 U792 ( .A1(n868), .A2(n942), .ZN(n730) );
  NAND2_X1 U793 ( .A1(G117), .A2(n879), .ZN(n722) );
  NAND2_X1 U794 ( .A1(G129), .A2(n880), .ZN(n721) );
  NAND2_X1 U795 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U796 ( .A1(n876), .A2(G105), .ZN(n723) );
  XOR2_X1 U797 ( .A(KEYINPUT38), .B(n723), .Z(n724) );
  NOR2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U799 ( .A(n726), .B(KEYINPUT94), .ZN(n728) );
  NAND2_X1 U800 ( .A1(G141), .A2(n875), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n890) );
  AND2_X1 U802 ( .A1(G1996), .A2(n890), .ZN(n729) );
  NOR2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n923) );
  INV_X1 U804 ( .A(n750), .ZN(n731) );
  NOR2_X1 U805 ( .A1(n923), .A2(n731), .ZN(n740) );
  INV_X1 U806 ( .A(n740), .ZN(n732) );
  NAND2_X1 U807 ( .A1(n744), .A2(n732), .ZN(n734) );
  XOR2_X1 U808 ( .A(G1986), .B(KEYINPUT91), .Z(n733) );
  XNOR2_X1 U809 ( .A(G290), .B(n733), .ZN(n969) );
  AND2_X1 U810 ( .A1(n942), .A2(n868), .ZN(n917) );
  NOR2_X1 U811 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n917), .A2(n737), .ZN(n738) );
  XOR2_X1 U813 ( .A(KEYINPUT105), .B(n738), .Z(n739) );
  NOR2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n890), .ZN(n934) );
  NOR2_X1 U816 ( .A1(n741), .A2(n934), .ZN(n742) );
  XNOR2_X1 U817 ( .A(n742), .B(KEYINPUT106), .ZN(n743) );
  XNOR2_X1 U818 ( .A(n743), .B(KEYINPUT39), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n748) );
  NOR2_X1 U820 ( .A1(n746), .A2(n889), .ZN(n747) );
  XNOR2_X1 U821 ( .A(n747), .B(KEYINPUT107), .ZN(n931) );
  NAND2_X1 U822 ( .A1(n748), .A2(n931), .ZN(n749) );
  XNOR2_X1 U823 ( .A(KEYINPUT108), .B(n749), .ZN(n751) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U826 ( .A(n754), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U827 ( .A(G57), .ZN(G237) );
  INV_X1 U828 ( .A(G132), .ZN(G219) );
  INV_X1 U829 ( .A(G82), .ZN(G220) );
  NOR2_X1 U830 ( .A1(n755), .A2(n756), .ZN(G160) );
  NAND2_X1 U831 ( .A1(G94), .A2(G452), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n757), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n758) );
  XNOR2_X1 U834 ( .A(n758), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U835 ( .A(G223), .ZN(n824) );
  NAND2_X1 U836 ( .A1(n824), .A2(G567), .ZN(n759) );
  XOR2_X1 U837 ( .A(KEYINPUT11), .B(n759), .Z(G234) );
  XOR2_X1 U838 ( .A(G860), .B(KEYINPUT76), .Z(n766) );
  OR2_X1 U839 ( .A1(n766), .A2(n972), .ZN(G153) );
  XNOR2_X1 U840 ( .A(G171), .B(KEYINPUT77), .ZN(G301) );
  NAND2_X1 U841 ( .A1(G868), .A2(G301), .ZN(n760) );
  XNOR2_X1 U842 ( .A(n760), .B(KEYINPUT78), .ZN(n762) );
  INV_X1 U843 ( .A(G868), .ZN(n806) );
  INV_X1 U844 ( .A(n967), .ZN(n769) );
  NAND2_X1 U845 ( .A1(n806), .A2(n769), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U847 ( .A(KEYINPUT80), .B(n763), .ZN(G284) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n765) );
  NOR2_X1 U849 ( .A1(G286), .A2(n806), .ZN(n764) );
  NOR2_X1 U850 ( .A1(n765), .A2(n764), .ZN(G297) );
  NAND2_X1 U851 ( .A1(n766), .A2(G559), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n767), .A2(n967), .ZN(n768) );
  XNOR2_X1 U853 ( .A(n768), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 U854 ( .A1(G559), .A2(n769), .ZN(n770) );
  NAND2_X1 U855 ( .A1(n770), .A2(G868), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n972), .A2(n806), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(G282) );
  XNOR2_X1 U858 ( .A(G2100), .B(KEYINPUT81), .ZN(n781) );
  NAND2_X1 U859 ( .A1(G111), .A2(n879), .ZN(n774) );
  NAND2_X1 U860 ( .A1(G135), .A2(n875), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G123), .A2(n880), .ZN(n775) );
  XNOR2_X1 U863 ( .A(n775), .B(KEYINPUT18), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G99), .A2(n876), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n916) );
  XNOR2_X1 U867 ( .A(n916), .B(G2096), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(G156) );
  NAND2_X1 U869 ( .A1(n967), .A2(G559), .ZN(n803) );
  XNOR2_X1 U870 ( .A(n972), .B(n803), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n782), .A2(G860), .ZN(n796) );
  NAND2_X1 U872 ( .A1(G67), .A2(n783), .ZN(n784) );
  XNOR2_X1 U873 ( .A(n784), .B(KEYINPUT84), .ZN(n794) );
  NAND2_X1 U874 ( .A1(n785), .A2(G55), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G93), .A2(n786), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G80), .A2(n789), .ZN(n790) );
  XNOR2_X1 U878 ( .A(KEYINPUT83), .B(n790), .ZN(n791) );
  NOR2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n805) );
  XOR2_X1 U881 ( .A(n805), .B(KEYINPUT82), .Z(n795) );
  XNOR2_X1 U882 ( .A(n796), .B(n795), .ZN(G145) );
  XNOR2_X1 U883 ( .A(KEYINPUT19), .B(G288), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(n805), .ZN(n800) );
  XNOR2_X1 U885 ( .A(G305), .B(G299), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n798), .B(n972), .ZN(n799) );
  XNOR2_X1 U887 ( .A(n800), .B(n799), .ZN(n802) );
  XNOR2_X1 U888 ( .A(G290), .B(G166), .ZN(n801) );
  XNOR2_X1 U889 ( .A(n802), .B(n801), .ZN(n895) );
  XNOR2_X1 U890 ( .A(n803), .B(n895), .ZN(n804) );
  NAND2_X1 U891 ( .A1(n804), .A2(G868), .ZN(n808) );
  NAND2_X1 U892 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U894 ( .A1(G2084), .A2(G2078), .ZN(n809) );
  XOR2_X1 U895 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U896 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U897 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U898 ( .A1(n812), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U899 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U900 ( .A1(G220), .A2(G219), .ZN(n813) );
  XOR2_X1 U901 ( .A(KEYINPUT22), .B(n813), .Z(n814) );
  NOR2_X1 U902 ( .A1(G218), .A2(n814), .ZN(n815) );
  NAND2_X1 U903 ( .A1(G96), .A2(n815), .ZN(n829) );
  NAND2_X1 U904 ( .A1(G2106), .A2(n829), .ZN(n819) );
  NAND2_X1 U905 ( .A1(G69), .A2(G120), .ZN(n816) );
  NOR2_X1 U906 ( .A1(G237), .A2(n816), .ZN(n817) );
  NAND2_X1 U907 ( .A1(G108), .A2(n817), .ZN(n830) );
  NAND2_X1 U908 ( .A1(G567), .A2(n830), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U910 ( .A(KEYINPUT88), .B(n820), .Z(G319) );
  INV_X1 U911 ( .A(G319), .ZN(n822) );
  NAND2_X1 U912 ( .A1(G661), .A2(G483), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n828) );
  NAND2_X1 U914 ( .A1(n828), .A2(G36), .ZN(n823) );
  XOR2_X1 U915 ( .A(KEYINPUT89), .B(n823), .Z(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n824), .ZN(G217) );
  NAND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n825) );
  XNOR2_X1 U918 ( .A(KEYINPUT111), .B(n825), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n826), .A2(G661), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XOR2_X1 U928 ( .A(G2474), .B(G1956), .Z(n832) );
  XNOR2_X1 U929 ( .A(G1986), .B(G1961), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U931 ( .A(n833), .B(KEYINPUT113), .Z(n835) );
  XNOR2_X1 U932 ( .A(G1996), .B(G1991), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U934 ( .A(G1976), .B(G1966), .Z(n837) );
  XNOR2_X1 U935 ( .A(G1981), .B(G1971), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U937 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U938 ( .A(KEYINPUT41), .B(KEYINPUT114), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(G229) );
  XOR2_X1 U940 ( .A(G2100), .B(KEYINPUT43), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2072), .B(G2678), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(n844), .B(KEYINPUT112), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2090), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2096), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2084), .B(G2078), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(G227) );
  NAND2_X1 U950 ( .A1(G112), .A2(n879), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G136), .A2(n875), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U953 ( .A1(G124), .A2(n880), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G100), .A2(n876), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U957 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U958 ( .A1(G118), .A2(n879), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n858), .B(KEYINPUT116), .ZN(n867) );
  NAND2_X1 U960 ( .A1(G130), .A2(n880), .ZN(n859) );
  XNOR2_X1 U961 ( .A(KEYINPUT115), .B(n859), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G142), .A2(n875), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G106), .A2(n876), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U965 ( .A(KEYINPUT45), .B(n862), .ZN(n863) );
  XNOR2_X1 U966 ( .A(KEYINPUT117), .B(n863), .ZN(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n872) );
  XOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n870) );
  XNOR2_X1 U970 ( .A(n868), .B(KEYINPUT118), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n874) );
  XNOR2_X1 U973 ( .A(G162), .B(n916), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n886) );
  NAND2_X1 U975 ( .A1(G139), .A2(n875), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G103), .A2(n876), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U978 ( .A1(G115), .A2(n879), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G127), .A2(n880), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U981 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n924) );
  XOR2_X1 U983 ( .A(n886), .B(n924), .Z(n888) );
  XNOR2_X1 U984 ( .A(G160), .B(G164), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U986 ( .A(n890), .B(n889), .Z(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U988 ( .A1(G37), .A2(n893), .ZN(n894) );
  XOR2_X1 U989 ( .A(KEYINPUT119), .B(n894), .Z(G395) );
  XOR2_X1 U990 ( .A(n895), .B(n967), .Z(n897) );
  XNOR2_X1 U991 ( .A(G286), .B(G171), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U993 ( .A1(G37), .A2(n898), .ZN(G397) );
  XNOR2_X1 U994 ( .A(G2443), .B(G2427), .ZN(n908) );
  XOR2_X1 U995 ( .A(G2430), .B(KEYINPUT110), .Z(n900) );
  XNOR2_X1 U996 ( .A(G2454), .B(G2435), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U998 ( .A(G2438), .B(KEYINPUT109), .Z(n902) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G2451), .B(G2446), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n909), .A2(G14), .ZN(n915) );
  NAND2_X1 U1006 ( .A1(n915), .A2(G319), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n915), .ZN(G401) );
  XNOR2_X1 U1015 ( .A(G160), .B(G2084), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n930) );
  XNOR2_X1 U1020 ( .A(G2072), .B(n924), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(G164), .B(G2078), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT50), .B(n927), .Z(n928) );
  XNOR2_X1 U1024 ( .A(KEYINPUT121), .B(n928), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n938) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1029 ( .A(KEYINPUT120), .B(n935), .Z(n936) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n936), .Z(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n963) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n963), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(G29), .ZN(n1021) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n958) );
  XNOR2_X1 U1037 ( .A(G25), .B(n942), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1039 ( .A(G32), .B(n944), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n952) );
  XOR2_X1 U1044 ( .A(G27), .B(n949), .Z(n950) );
  XNOR2_X1 U1045 ( .A(KEYINPUT122), .B(n950), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n953), .B(KEYINPUT123), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n963), .B(n962), .ZN(n965) );
  INV_X1 U1055 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n966), .ZN(n1019) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XNOR2_X1 U1059 ( .A(n967), .B(G1348), .ZN(n971) );
  XOR2_X1 U1060 ( .A(G171), .B(G1961), .Z(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(G1341), .B(n972), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n983) );
  NAND2_X1 U1065 ( .A1(G1971), .A2(G303), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(G1956), .B(G299), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1070 ( .A(KEYINPUT124), .B(n981), .Z(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(KEYINPUT125), .B(n984), .ZN(n989) );
  XOR2_X1 U1073 ( .A(G168), .B(G1966), .Z(n985) );
  NOR2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1075 ( .A(KEYINPUT57), .B(n987), .Z(n988) );
  NAND2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n1017) );
  INV_X1 U1078 ( .A(G16), .ZN(n1015) );
  XNOR2_X1 U1079 ( .A(KEYINPUT59), .B(G1348), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(n992), .B(G4), .ZN(n997) );
  XOR2_X1 U1081 ( .A(G1981), .B(KEYINPUT127), .Z(n993) );
  XNOR2_X1 U1082 ( .A(G6), .B(n993), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G20), .B(G1956), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(KEYINPUT126), .B(G1341), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G19), .B(n998), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(KEYINPUT60), .B(n1001), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G21), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G1961), .B(G5), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(G1986), .B(G24), .Z(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

