

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n727), .A2(G1341), .ZN(n520) );
  XOR2_X1 U554 ( .A(KEYINPUT97), .B(n692), .Z(n521) );
  XOR2_X1 U555 ( .A(KEYINPUT83), .B(n802), .Z(n522) );
  NOR2_X1 U556 ( .A1(n927), .A2(n520), .ZN(n685) );
  AND2_X1 U557 ( .A1(n686), .A2(n685), .ZN(n693) );
  NAND2_X1 U558 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U559 ( .A(n708), .B(KEYINPUT29), .ZN(n713) );
  AND2_X1 U560 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n785) );
  NAND2_X1 U562 ( .A1(n803), .A2(n522), .ZN(n804) );
  NOR2_X1 U563 ( .A1(n626), .A2(G651), .ZN(n647) );
  AND2_X1 U564 ( .A1(n527), .A2(G2104), .ZN(n888) );
  NOR2_X1 U565 ( .A1(n531), .A2(n530), .ZN(G160) );
  AND2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U567 ( .A1(n891), .A2(G113), .ZN(n525) );
  INV_X1 U568 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U569 ( .A1(G101), .A2(n888), .ZN(n523) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n523), .Z(n524) );
  NAND2_X1 U571 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XOR2_X2 U573 ( .A(KEYINPUT17), .B(n526), .Z(n887) );
  NAND2_X1 U574 ( .A1(G137), .A2(n887), .ZN(n529) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n527), .ZN(n892) );
  NAND2_X1 U576 ( .A1(G125), .A2(n892), .ZN(n528) );
  NAND2_X1 U577 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U578 ( .A1(G138), .A2(n887), .ZN(n537) );
  AND2_X1 U579 ( .A1(G102), .A2(n888), .ZN(n535) );
  NAND2_X1 U580 ( .A1(G114), .A2(n891), .ZN(n533) );
  NAND2_X1 U581 ( .A1(G126), .A2(n892), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U583 ( .A1(n535), .A2(n534), .ZN(n536) );
  AND2_X1 U584 ( .A1(n537), .A2(n536), .ZN(G164) );
  INV_X1 U585 ( .A(G651), .ZN(n541) );
  NOR2_X1 U586 ( .A1(G543), .A2(n541), .ZN(n538) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n538), .Z(n641) );
  NAND2_X1 U588 ( .A1(G64), .A2(n641), .ZN(n540) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n626) );
  NAND2_X1 U590 ( .A1(G52), .A2(n647), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n547) );
  NOR2_X1 U592 ( .A1(n626), .A2(n541), .ZN(n645) );
  NAND2_X1 U593 ( .A1(G77), .A2(n645), .ZN(n544) );
  NOR2_X1 U594 ( .A1(G543), .A2(G651), .ZN(n542) );
  XOR2_X1 U595 ( .A(KEYINPUT65), .B(n542), .Z(n639) );
  NAND2_X1 U596 ( .A1(G90), .A2(n639), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n545), .Z(n546) );
  NOR2_X1 U599 ( .A1(n547), .A2(n546), .ZN(G171) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  NAND2_X1 U604 ( .A1(n641), .A2(G62), .ZN(n548) );
  XOR2_X1 U605 ( .A(KEYINPUT79), .B(n548), .Z(n550) );
  NAND2_X1 U606 ( .A1(n647), .A2(G50), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U608 ( .A(KEYINPUT80), .B(n551), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G75), .A2(n645), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G88), .A2(n639), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U612 ( .A1(n555), .A2(n554), .ZN(G166) );
  NAND2_X1 U613 ( .A1(n639), .A2(G89), .ZN(n556) );
  XNOR2_X1 U614 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U615 ( .A1(G76), .A2(n645), .ZN(n557) );
  NAND2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U617 ( .A(KEYINPUT5), .B(n559), .Z(n566) );
  NAND2_X1 U618 ( .A1(n641), .A2(G63), .ZN(n560) );
  XOR2_X1 U619 ( .A(KEYINPUT69), .B(n560), .Z(n562) );
  NAND2_X1 U620 ( .A1(n647), .A2(G51), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n564) );
  XOR2_X1 U622 ( .A(KEYINPUT6), .B(KEYINPUT70), .Z(n563) );
  XOR2_X1 U623 ( .A(n564), .B(n563), .Z(n565) );
  NOR2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U625 ( .A(KEYINPUT71), .B(KEYINPUT7), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n568), .B(n567), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U630 ( .A(G223), .ZN(n822) );
  NAND2_X1 U631 ( .A1(n822), .A2(G567), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U633 ( .A1(n641), .A2(G56), .ZN(n571) );
  XNOR2_X1 U634 ( .A(KEYINPUT14), .B(n571), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n639), .A2(G81), .ZN(n572) );
  XNOR2_X1 U636 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G68), .A2(n645), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT13), .B(n575), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT67), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n647), .A2(G43), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n927) );
  INV_X1 U644 ( .A(G860), .ZN(n623) );
  OR2_X1 U645 ( .A1(n927), .A2(n623), .ZN(G153) );
  INV_X1 U646 ( .A(G171), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT68), .ZN(n590) );
  NAND2_X1 U649 ( .A1(G66), .A2(n641), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G92), .A2(n639), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G79), .A2(n645), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G54), .A2(n647), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT15), .B(n588), .Z(n930) );
  OR2_X1 U657 ( .A1(G868), .A2(n930), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U659 ( .A1(G65), .A2(n641), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G53), .A2(n647), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G78), .A2(n645), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G91), .A2(n639), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n931) );
  INV_X1 U666 ( .A(n931), .ZN(G299) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n597), .B(KEYINPUT72), .ZN(n599) );
  INV_X1 U669 ( .A(G868), .ZN(n662) );
  NOR2_X1 U670 ( .A1(n662), .A2(G286), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n623), .A2(G559), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n600), .A2(n930), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U675 ( .A1(G868), .A2(n927), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G868), .A2(n930), .ZN(n602) );
  NOR2_X1 U677 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U678 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U679 ( .A1(G123), .A2(n892), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n891), .A2(G111), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G135), .A2(n887), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G99), .A2(n888), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n1003) );
  XNOR2_X1 U687 ( .A(n1003), .B(G2096), .ZN(n613) );
  INV_X1 U688 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U690 ( .A1(G67), .A2(n641), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G55), .A2(n647), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n616), .B(KEYINPUT75), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G80), .A2(n645), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n639), .A2(G93), .ZN(n619) );
  XOR2_X1 U697 ( .A(KEYINPUT74), .B(n619), .Z(n620) );
  OR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n661) );
  NAND2_X1 U699 ( .A1(G559), .A2(n930), .ZN(n622) );
  XOR2_X1 U700 ( .A(n927), .B(n622), .Z(n659) );
  NAND2_X1 U701 ( .A1(n623), .A2(n659), .ZN(n624) );
  XNOR2_X1 U702 ( .A(n624), .B(KEYINPUT73), .ZN(n625) );
  XOR2_X1 U703 ( .A(n661), .B(n625), .Z(G145) );
  NAND2_X1 U704 ( .A1(G49), .A2(n647), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G87), .A2(n626), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n641), .A2(n629), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G651), .A2(G74), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G60), .A2(n641), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G47), .A2(n647), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G72), .A2(n645), .ZN(n634) );
  XOR2_X1 U714 ( .A(KEYINPUT66), .B(n634), .Z(n635) );
  NOR2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(G85), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U718 ( .A1(n639), .A2(G86), .ZN(n640) );
  XNOR2_X1 U719 ( .A(n640), .B(KEYINPUT76), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G61), .A2(n641), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U722 ( .A(KEYINPUT77), .B(n644), .ZN(n652) );
  NAND2_X1 U723 ( .A1(G73), .A2(n645), .ZN(n646) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n646), .Z(n650) );
  NAND2_X1 U725 ( .A1(n647), .A2(G48), .ZN(n648) );
  XOR2_X1 U726 ( .A(KEYINPUT78), .B(n648), .Z(n649) );
  NOR2_X1 U727 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(G305) );
  XOR2_X1 U729 ( .A(KEYINPUT19), .B(n661), .Z(n654) );
  XNOR2_X1 U730 ( .A(G288), .B(KEYINPUT81), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U732 ( .A(n931), .B(n655), .ZN(n657) );
  XNOR2_X1 U733 ( .A(G290), .B(G166), .ZN(n656) );
  XNOR2_X1 U734 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n658), .B(G305), .ZN(n854) );
  XNOR2_X1 U736 ( .A(n659), .B(n854), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n660), .A2(G868), .ZN(n664) );
  NAND2_X1 U738 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U742 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U744 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U746 ( .A1(G120), .A2(G69), .ZN(n669) );
  NOR2_X1 U747 ( .A1(G237), .A2(n669), .ZN(n670) );
  XNOR2_X1 U748 ( .A(KEYINPUT82), .B(n670), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n671), .A2(G108), .ZN(n828) );
  NAND2_X1 U750 ( .A1(n828), .A2(G567), .ZN(n676) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n672) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n672), .Z(n673) );
  NOR2_X1 U753 ( .A1(G218), .A2(n673), .ZN(n674) );
  NAND2_X1 U754 ( .A1(G96), .A2(n674), .ZN(n829) );
  NAND2_X1 U755 ( .A1(n829), .A2(G2106), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n830) );
  NAND2_X1 U757 ( .A1(G483), .A2(G661), .ZN(n677) );
  NOR2_X1 U758 ( .A1(n830), .A2(n677), .ZN(n827) );
  NAND2_X1 U759 ( .A1(n827), .A2(G36), .ZN(G176) );
  INV_X1 U760 ( .A(G166), .ZN(G303) );
  NAND2_X1 U761 ( .A1(G160), .A2(G40), .ZN(n786) );
  INV_X1 U762 ( .A(n786), .ZN(n678) );
  NAND2_X1 U763 ( .A1(n678), .A2(n785), .ZN(n679) );
  XNOR2_X2 U764 ( .A(n679), .B(KEYINPUT64), .ZN(n727) );
  NOR2_X1 U765 ( .A1(n727), .A2(G2084), .ZN(n680) );
  XOR2_X1 U766 ( .A(KEYINPUT92), .B(n680), .Z(n714) );
  INV_X1 U767 ( .A(n714), .ZN(n681) );
  NAND2_X1 U768 ( .A1(n681), .A2(G8), .ZN(n726) );
  NAND2_X1 U769 ( .A1(n727), .A2(G8), .ZN(n762) );
  NOR2_X1 U770 ( .A1(G1966), .A2(n762), .ZN(n716) );
  INV_X1 U771 ( .A(n716), .ZN(n724) );
  INV_X1 U772 ( .A(G1996), .ZN(n682) );
  NOR2_X1 U773 ( .A1(n727), .A2(n682), .ZN(n684) );
  XNOR2_X1 U774 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n683) );
  XNOR2_X1 U775 ( .A(n684), .B(n683), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n930), .A2(n693), .ZN(n687) );
  XNOR2_X1 U777 ( .A(n687), .B(KEYINPUT96), .ZN(n691) );
  NOR2_X1 U778 ( .A1(G2067), .A2(n727), .ZN(n689) );
  INV_X1 U779 ( .A(n727), .ZN(n709) );
  NOR2_X1 U780 ( .A1(G1348), .A2(n709), .ZN(n688) );
  NOR2_X1 U781 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X1 U783 ( .A1(n930), .A2(n693), .ZN(n700) );
  XOR2_X1 U784 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n695) );
  NAND2_X1 U785 ( .A1(G2072), .A2(n709), .ZN(n694) );
  XNOR2_X1 U786 ( .A(n695), .B(n694), .ZN(n697) );
  INV_X1 U787 ( .A(G1956), .ZN(n840) );
  NOR2_X1 U788 ( .A1(n709), .A2(n840), .ZN(n696) );
  NOR2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n703) );
  NOR2_X1 U790 ( .A1(n703), .A2(n931), .ZN(n699) );
  XOR2_X1 U791 ( .A(KEYINPUT94), .B(KEYINPUT28), .Z(n698) );
  XNOR2_X1 U792 ( .A(n699), .B(n698), .ZN(n702) );
  AND2_X1 U793 ( .A1(n700), .A2(n702), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n521), .A2(n701), .ZN(n707) );
  INV_X1 U795 ( .A(n702), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n703), .A2(n931), .ZN(n704) );
  OR2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U798 ( .A(G2078), .B(KEYINPUT25), .ZN(n987) );
  NAND2_X1 U799 ( .A1(n709), .A2(n987), .ZN(n711) );
  INV_X1 U800 ( .A(G1961), .ZN(n956) );
  NAND2_X1 U801 ( .A1(n727), .A2(n956), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n719) );
  NAND2_X1 U803 ( .A1(n719), .A2(G171), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n735) );
  NAND2_X1 U805 ( .A1(G8), .A2(n714), .ZN(n715) );
  NOR2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U807 ( .A(KEYINPUT30), .B(n717), .Z(n718) );
  NOR2_X1 U808 ( .A1(G168), .A2(n718), .ZN(n721) );
  NOR2_X1 U809 ( .A1(G171), .A2(n719), .ZN(n720) );
  NOR2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U811 ( .A(KEYINPUT31), .B(n722), .Z(n733) );
  NAND2_X1 U812 ( .A1(n735), .A2(n733), .ZN(n723) );
  NAND2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n742) );
  INV_X1 U814 ( .A(G8), .ZN(n732) );
  NOR2_X1 U815 ( .A1(n727), .A2(G2090), .ZN(n729) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n762), .ZN(n728) );
  NOR2_X1 U817 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U818 ( .A1(n730), .A2(G303), .ZN(n731) );
  OR2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n736) );
  AND2_X1 U820 ( .A1(n733), .A2(n736), .ZN(n734) );
  NAND2_X1 U821 ( .A1(n735), .A2(n734), .ZN(n739) );
  INV_X1 U822 ( .A(n736), .ZN(n737) );
  OR2_X1 U823 ( .A1(n737), .A2(G286), .ZN(n738) );
  NAND2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U825 ( .A(n740), .B(KEYINPUT32), .ZN(n741) );
  NAND2_X1 U826 ( .A1(n742), .A2(n741), .ZN(n758) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n743) );
  XOR2_X1 U828 ( .A(KEYINPUT98), .B(n743), .Z(n933) );
  NAND2_X1 U829 ( .A1(n758), .A2(n933), .ZN(n745) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n749) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n936) );
  INV_X1 U833 ( .A(n936), .ZN(n746) );
  OR2_X1 U834 ( .A1(n746), .A2(n762), .ZN(n747) );
  OR2_X1 U835 ( .A1(KEYINPUT99), .A2(n747), .ZN(n748) );
  NOR2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U837 ( .A1(KEYINPUT33), .A2(n750), .ZN(n754) );
  XNOR2_X1 U838 ( .A(n933), .B(KEYINPUT99), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U840 ( .A1(n762), .A2(n752), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n922) );
  AND2_X1 U843 ( .A1(n755), .A2(n922), .ZN(n767) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U845 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n759), .A2(n762), .ZN(n765) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n760) );
  XOR2_X1 U849 ( .A(n760), .B(KEYINPUT24), .Z(n761) );
  NOR2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U851 ( .A(KEYINPUT91), .B(n763), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n805) );
  NAND2_X1 U854 ( .A1(n891), .A2(G107), .ZN(n770) );
  NAND2_X1 U855 ( .A1(G95), .A2(n888), .ZN(n768) );
  XOR2_X1 U856 ( .A(KEYINPUT87), .B(n768), .Z(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G131), .A2(n887), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G119), .A2(n892), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n868) );
  INV_X1 U862 ( .A(G1991), .ZN(n981) );
  NOR2_X1 U863 ( .A1(n868), .A2(n981), .ZN(n784) );
  XOR2_X1 U864 ( .A(KEYINPUT38), .B(KEYINPUT88), .Z(n776) );
  NAND2_X1 U865 ( .A1(G105), .A2(n888), .ZN(n775) );
  XNOR2_X1 U866 ( .A(n776), .B(n775), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G141), .A2(n887), .ZN(n778) );
  NAND2_X1 U868 ( .A1(G117), .A2(n891), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n892), .A2(G129), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n880) );
  AND2_X1 U873 ( .A1(n880), .A2(G1996), .ZN(n783) );
  NOR2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n1005) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n817) );
  INV_X1 U876 ( .A(n817), .ZN(n787) );
  NOR2_X1 U877 ( .A1(n1005), .A2(n787), .ZN(n808) );
  XNOR2_X1 U878 ( .A(KEYINPUT89), .B(n808), .ZN(n800) );
  XNOR2_X1 U879 ( .A(KEYINPUT85), .B(KEYINPUT36), .ZN(n798) );
  NAND2_X1 U880 ( .A1(G140), .A2(n887), .ZN(n789) );
  NAND2_X1 U881 ( .A1(G104), .A2(n888), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U883 ( .A(KEYINPUT34), .B(n790), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G116), .A2(n891), .ZN(n792) );
  NAND2_X1 U885 ( .A1(G128), .A2(n892), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U887 ( .A(n793), .B(KEYINPUT35), .Z(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U889 ( .A(KEYINPUT84), .B(n796), .Z(n797) );
  XNOR2_X1 U890 ( .A(n798), .B(n797), .ZN(n901) );
  XNOR2_X1 U891 ( .A(KEYINPUT37), .B(G2067), .ZN(n813) );
  NOR2_X1 U892 ( .A1(n901), .A2(n813), .ZN(n799) );
  XNOR2_X1 U893 ( .A(KEYINPUT86), .B(n799), .ZN(n1011) );
  NAND2_X1 U894 ( .A1(n817), .A2(n1011), .ZN(n811) );
  NAND2_X1 U895 ( .A1(n800), .A2(n811), .ZN(n801) );
  XOR2_X1 U896 ( .A(KEYINPUT90), .B(n801), .Z(n803) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n944) );
  NAND2_X1 U898 ( .A1(n817), .A2(n944), .ZN(n802) );
  OR2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n819) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n880), .ZN(n1000) );
  AND2_X1 U901 ( .A1(n981), .A2(n868), .ZN(n1007) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n1007), .A2(n806), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n1000), .A2(n809), .ZN(n810) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n810), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n901), .A2(n813), .ZN(n814) );
  XNOR2_X1 U909 ( .A(KEYINPUT100), .B(n814), .ZN(n1013) );
  NAND2_X1 U910 ( .A1(n815), .A2(n1013), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n821) );
  XOR2_X1 U913 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n820) );
  XNOR2_X1 U914 ( .A(n821), .B(n820), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n822), .ZN(G217) );
  INV_X1 U916 ( .A(G661), .ZN(n824) );
  NAND2_X1 U917 ( .A1(G2), .A2(G15), .ZN(n823) );
  NOR2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  XOR2_X1 U919 ( .A(KEYINPUT104), .B(n825), .Z(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G69), .ZN(G235) );
  NOR2_X1 U927 ( .A1(n829), .A2(n828), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  INV_X1 U929 ( .A(n830), .ZN(G319) );
  XOR2_X1 U930 ( .A(G1961), .B(G1966), .Z(n832) );
  XNOR2_X1 U931 ( .A(G1981), .B(G1976), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U933 ( .A(G1971), .B(G1986), .Z(n834) );
  XNOR2_X1 U934 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U937 ( .A(KEYINPUT107), .B(G2474), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U939 ( .A(KEYINPUT41), .B(n839), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(G229) );
  XOR2_X1 U941 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n843) );
  XNOR2_X1 U942 ( .A(G2678), .B(KEYINPUT43), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2090), .Z(n845) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2096), .B(G2100), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U950 ( .A(G2078), .B(G2084), .Z(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U952 ( .A(KEYINPUT115), .B(G286), .Z(n853) );
  XNOR2_X1 U953 ( .A(G171), .B(n930), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n927), .B(n854), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  NOR2_X1 U957 ( .A1(G37), .A2(n857), .ZN(n858) );
  XNOR2_X1 U958 ( .A(KEYINPUT116), .B(n858), .ZN(G397) );
  NAND2_X1 U959 ( .A1(G100), .A2(n888), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G112), .A2(n891), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U962 ( .A(KEYINPUT108), .B(n861), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n892), .A2(G124), .ZN(n862) );
  XOR2_X1 U964 ( .A(KEYINPUT44), .B(n862), .Z(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n887), .A2(G136), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U968 ( .A(KEYINPUT109), .B(n867), .ZN(G162) );
  XNOR2_X1 U969 ( .A(n868), .B(n1003), .ZN(n878) );
  NAND2_X1 U970 ( .A1(G118), .A2(n891), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G130), .A2(n892), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G142), .A2(n887), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G106), .A2(n888), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U976 ( .A(KEYINPUT45), .B(n873), .Z(n874) );
  XNOR2_X1 U977 ( .A(KEYINPUT110), .B(n874), .ZN(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U980 ( .A(n879), .B(G162), .Z(n882) );
  XOR2_X1 U981 ( .A(G160), .B(n880), .Z(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n886) );
  XOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n884) );
  XNOR2_X1 U984 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(n886), .B(n885), .Z(n900) );
  NAND2_X1 U987 ( .A1(G139), .A2(n887), .ZN(n890) );
  NAND2_X1 U988 ( .A1(G103), .A2(n888), .ZN(n889) );
  NAND2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n898) );
  NAND2_X1 U990 ( .A1(G115), .A2(n891), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G127), .A2(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U993 ( .A(KEYINPUT47), .B(n895), .ZN(n896) );
  XNOR2_X1 U994 ( .A(KEYINPUT111), .B(n896), .ZN(n897) );
  NOR2_X1 U995 ( .A1(n898), .A2(n897), .ZN(n1015) );
  XNOR2_X1 U996 ( .A(G164), .B(n1015), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G37), .A2(n903), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(KEYINPUT114), .B(n904), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(G2427), .B(KEYINPUT102), .ZN(n914) );
  XOR2_X1 U1002 ( .A(G2430), .B(G2446), .Z(n906) );
  XNOR2_X1 U1003 ( .A(G2435), .B(G2438), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1005 ( .A(G2454), .B(KEYINPUT103), .Z(n908) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1008 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1009 ( .A(G2451), .B(G2443), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(n915), .A2(G14), .ZN(n921) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G397), .A2(G395), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n921), .ZN(G401) );
  XNOR2_X1 U1021 ( .A(G16), .B(KEYINPUT56), .ZN(n948) );
  XNOR2_X1 U1022 ( .A(G1971), .B(G166), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G168), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(n924), .B(KEYINPUT57), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(G1341), .B(n927), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n946) );
  XNOR2_X1 U1029 ( .A(n930), .B(G1348), .ZN(n942) );
  XNOR2_X1 U1030 ( .A(n931), .B(G1956), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(KEYINPUT123), .ZN(n935) );
  INV_X1 U1032 ( .A(n933), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n940) );
  XOR2_X1 U1035 ( .A(G1961), .B(G171), .Z(n938) );
  XNOR2_X1 U1036 ( .A(KEYINPUT122), .B(n938), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT124), .B(n949), .ZN(n1029) );
  XOR2_X1 U1043 ( .A(G1986), .B(KEYINPUT126), .Z(n950) );
  XNOR2_X1 U1044 ( .A(G24), .B(n950), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G1976), .B(G23), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G1971), .B(G22), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1049 ( .A(KEYINPUT58), .B(n955), .Z(n971) );
  XOR2_X1 U1050 ( .A(G1966), .B(G21), .Z(n958) );
  XNOR2_X1 U1051 ( .A(n956), .B(G5), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n969) );
  XNOR2_X1 U1053 ( .A(G1956), .B(G20), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G1981), .B(G6), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G19), .B(G1341), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT125), .B(n961), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(G1348), .B(KEYINPUT59), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(G4), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(KEYINPUT60), .B(n967), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT127), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT61), .B(n973), .ZN(n975) );
  INV_X1 U1067 ( .A(G16), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n976), .A2(G11), .ZN(n1027) );
  XOR2_X1 U1070 ( .A(G34), .B(KEYINPUT121), .Z(n978) );
  XNOR2_X1 U1071 ( .A(G2084), .B(KEYINPUT54), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n978), .B(n977), .ZN(n996) );
  XNOR2_X1 U1073 ( .A(G2090), .B(G35), .ZN(n993) );
  XOR2_X1 U1074 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n991) );
  XNOR2_X1 U1075 ( .A(G1996), .B(G32), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(G33), .B(G2072), .ZN(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G25), .B(n981), .ZN(n982) );
  NAND2_X1 U1079 ( .A1(n982), .A2(G28), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(G26), .B(G2067), .ZN(n983) );
  NOR2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n989) );
  XOR2_X1 U1083 ( .A(G27), .B(n987), .Z(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(n991), .B(n990), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1087 ( .A(KEYINPUT120), .B(n994), .Z(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(G29), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(n998), .B(KEYINPUT55), .ZN(n1025) );
  XOR2_X1 U1091 ( .A(G2090), .B(G162), .Z(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1093 ( .A(KEYINPUT51), .B(n1001), .Z(n1009) );
  XOR2_X1 U1094 ( .A(G2084), .B(G160), .Z(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT117), .B(n1014), .ZN(n1021) );
  XOR2_X1 U1102 ( .A(G2072), .B(n1015), .Z(n1017) );
  XOR2_X1 U1103 ( .A(G164), .B(G2078), .Z(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(n1018), .B(KEYINPUT118), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(n1019), .B(KEYINPUT50), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(G29), .A2(n1023), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

