//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019;
  INV_X1    g000(.A(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(G227gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT28), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT27), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G183gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT27), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(KEYINPUT27), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(G183gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT67), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n206), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT26), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  AND4_X1   g023(.A1(KEYINPUT68), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT68), .B1(new_n226), .B2(new_n222), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n221), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT27), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n208), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n231), .A2(new_n232), .A3(new_n206), .A4(new_n217), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n237), .A3(new_n220), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n229), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n210), .A2(new_n217), .A3(KEYINPUT64), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(G183gat), .B2(G190gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n241), .A2(new_n242), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT25), .B1(new_n239), .B2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n235), .A2(new_n237), .A3(KEYINPUT25), .A4(new_n220), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n210), .A2(new_n217), .ZN(new_n249));
  NAND4_X1  g048(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n241), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n245), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n248), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OAI22_X1  g053(.A1(new_n218), .A2(new_n234), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(G113gat), .B2(G120gat), .ZN(new_n258));
  AND2_X1   g057(.A1(G113gat), .A2(G120gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n261), .B(new_n256), .C1(new_n259), .C2(new_n258), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n255), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n233), .A2(new_n229), .ZN(new_n267));
  AOI21_X1  g066(.A(G190gat), .B1(new_n212), .B2(new_n215), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n228), .B(new_n267), .C1(new_n268), .C2(new_n206), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n241), .A3(new_n249), .A4(new_n250), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n239), .A2(new_n270), .A3(KEYINPUT25), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n242), .A2(new_n244), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n241), .A2(new_n245), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n238), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n271), .B1(new_n274), .B2(KEYINPUT25), .ZN(new_n275));
  INV_X1    g074(.A(new_n265), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n269), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n205), .B1(new_n266), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n202), .B1(new_n278), .B2(KEYINPUT71), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n278), .B2(KEYINPUT71), .ZN(new_n281));
  INV_X1    g080(.A(new_n205), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n269), .A2(new_n275), .A3(new_n276), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n276), .B1(new_n269), .B2(new_n275), .ZN(new_n284));
  OAI211_X1 g083(.A(KEYINPUT71), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(KEYINPUT72), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n279), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT34), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n278), .A2(KEYINPUT71), .A3(new_n280), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(KEYINPUT72), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT32), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n266), .A2(new_n205), .A3(new_n277), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT70), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n266), .A2(new_n298), .A3(new_n205), .A4(new_n277), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT33), .B1(new_n297), .B2(new_n299), .ZN(new_n301));
  XOR2_X1   g100(.A(G15gat), .B(G43gat), .Z(new_n302));
  XNOR2_X1  g101(.A(G71gat), .B(G99gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n300), .A2(new_n301), .A3(new_n305), .ZN(new_n306));
  AOI221_X4 g105(.A(new_n295), .B1(KEYINPUT33), .B2(new_n304), .C1(new_n297), .C2(new_n299), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n294), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n283), .A2(new_n284), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n298), .B1(new_n309), .B2(new_n205), .ZN(new_n310));
  INV_X1    g109(.A(new_n299), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT32), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT33), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n310), .B2(new_n311), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n314), .A3(new_n304), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n300), .B1(new_n301), .B2(new_n305), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n315), .A2(new_n316), .A3(new_n293), .A4(new_n287), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n308), .A2(new_n317), .A3(KEYINPUT73), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n315), .A2(new_n316), .B1(new_n293), .B2(new_n287), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT36), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n317), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT36), .B1(new_n325), .B2(new_n319), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328));
  INV_X1    g127(.A(G50gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G22gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G141gat), .ZN(new_n335));
  INV_X1    g134(.A(G148gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338));
  AND2_X1   g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT2), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT76), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G155gat), .B(G162gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .A4(new_n343), .ZN(new_n351));
  INV_X1    g150(.A(new_n349), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n342), .A2(KEYINPUT75), .A3(KEYINPUT2), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n348), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n345), .A2(new_n351), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  INV_X1    g157(.A(G211gat), .ZN(new_n359));
  INV_X1    g158(.A(G218gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G211gat), .A2(G218gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n363), .B1(new_n366), .B2(new_n364), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n358), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT83), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT3), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(G197gat), .A2(G204gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n362), .B(new_n361), .C1(new_n375), .C2(new_n365), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT29), .B1(new_n376), .B2(new_n367), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT83), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n357), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n368), .A2(new_n369), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n357), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n383), .B2(new_n358), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n334), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n345), .A2(new_n351), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n356), .A2(new_n352), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n386), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n380), .B1(new_n388), .B2(KEYINPUT29), .ZN(new_n389));
  INV_X1    g188(.A(new_n357), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n370), .A2(KEYINPUT82), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n382), .B1(new_n377), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n394), .A3(new_n333), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n385), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n397), .B1(new_n385), .B2(new_n395), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n332), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n389), .A2(new_n394), .A3(new_n333), .ZN(new_n401));
  INV_X1    g200(.A(new_n378), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n382), .B1(new_n377), .B2(KEYINPUT83), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n390), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n333), .B1(new_n404), .B2(new_n389), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n396), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n395), .A3(new_n397), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n331), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n386), .A2(new_n265), .A3(new_n387), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n265), .B1(new_n386), .B2(new_n387), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n417));
  AND4_X1   g216(.A1(KEYINPUT4), .A2(new_n386), .A3(new_n265), .A4(new_n387), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT4), .B1(new_n357), .B2(new_n265), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n276), .B1(new_n357), .B2(new_n382), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n413), .B1(new_n422), .B2(new_n383), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n417), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n418), .B2(new_n419), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n386), .A2(new_n265), .A3(new_n387), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n357), .A2(KEYINPUT4), .A3(new_n265), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(KEYINPUT77), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n433), .B(new_n412), .C1(new_n421), .C2(new_n388), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT78), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n434), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT78), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n426), .A4(new_n431), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n424), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT0), .ZN(new_n441));
  XNOR2_X1  g240(.A(G57gat), .B(G85gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n443), .B(KEYINPUT84), .Z(new_n444));
  OAI21_X1  g243(.A(new_n411), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n435), .A2(new_n438), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n424), .A2(new_n443), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT79), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT79), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G8gat), .B(G36gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(G64gat), .B(G92gat), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n453), .B(new_n454), .Z(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(G226gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(new_n204), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n255), .B2(new_n358), .ZN(new_n459));
  INV_X1    g258(.A(new_n458), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n269), .B2(new_n275), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n381), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n255), .A2(new_n458), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT74), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(KEYINPUT74), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n463), .B1(new_n468), .B2(new_n381), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n456), .B1(new_n469), .B2(KEYINPUT37), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n459), .A2(new_n380), .A3(new_n461), .ZN(new_n471));
  INV_X1    g270(.A(new_n459), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n461), .A2(KEYINPUT74), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n465), .B(new_n460), .C1(new_n269), .C2(new_n275), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n471), .B1(new_n475), .B2(new_n380), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT38), .B1(new_n470), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n463), .B(new_n455), .C1(new_n468), .C2(new_n381), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n475), .A2(new_n381), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n477), .B1(new_n462), .B2(new_n380), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT38), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n483), .B(new_n456), .C1(KEYINPUT37), .C2(new_n469), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n443), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n439), .A2(new_n411), .A3(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n452), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n456), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n490));
  OR3_X1    g289(.A1(new_n469), .A2(KEYINPUT30), .A3(new_n456), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n439), .A2(new_n444), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n422), .A2(new_n383), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(new_n426), .A3(new_n431), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n413), .ZN(new_n497));
  XOR2_X1   g296(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n498));
  OAI21_X1  g297(.A(new_n444), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT39), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n414), .A2(new_n415), .A3(new_n413), .ZN(new_n501));
  AOI211_X1 g300(.A(new_n500), .B(new_n501), .C1(new_n496), .C2(new_n413), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n494), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT40), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n494), .B(new_n505), .C1(new_n499), .C2(new_n502), .ZN(new_n506));
  AND4_X1   g305(.A1(new_n492), .A2(new_n493), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n410), .B1(new_n488), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n492), .ZN(new_n509));
  INV_X1    g308(.A(new_n487), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n411), .B1(new_n439), .B2(new_n486), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n450), .B2(new_n451), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n512), .B2(KEYINPUT80), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT80), .ZN(new_n514));
  AOI211_X1 g313(.A(new_n514), .B(new_n511), .C1(new_n450), .C2(new_n451), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n509), .B(new_n409), .C1(new_n513), .C2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n327), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n318), .A2(new_n321), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n400), .A2(new_n520), .A3(new_n408), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n491), .B2(new_n490), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n452), .B2(new_n487), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n325), .A2(new_n319), .A3(new_n409), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n509), .B(new_n525), .C1(new_n513), .C2(new_n515), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n526), .B2(KEYINPUT35), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n518), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G183gat), .B(G211gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT97), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n532));
  INV_X1    g331(.A(G155gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n531), .B(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G57gat), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT95), .B1(new_n537), .B2(G64gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT95), .ZN(new_n539));
  INV_X1    g338(.A(G64gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n540), .A3(G57gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(G64gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n543), .A2(KEYINPUT96), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(KEYINPUT96), .ZN(new_n545));
  NAND2_X1  g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT9), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT94), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n547), .B1(new_n550), .B2(new_n546), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n550), .B2(new_n546), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n540), .A2(G57gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT9), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n553), .A2(new_n542), .B1(KEYINPUT94), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G231gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(new_n204), .ZN(new_n559));
  OR3_X1    g358(.A1(new_n557), .A2(KEYINPUT21), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n557), .B2(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G127gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n557), .A2(KEYINPUT21), .ZN(new_n565));
  XNOR2_X1  g364(.A(G15gat), .B(G22gat), .ZN(new_n566));
  INV_X1    g365(.A(G1gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT16), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(G1gat), .B2(new_n566), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G8gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n564), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n564), .A2(new_n573), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n536), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n574), .A3(new_n535), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT98), .Z(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G36gat), .ZN(new_n587));
  AND2_X1   g386(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G29gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n329), .B2(G43gat), .ZN(new_n595));
  INV_X1    g394(.A(G43gat), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT88), .B1(new_n596), .B2(G50gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n329), .A3(G43gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n600));
  AND4_X1   g399(.A1(new_n595), .A2(new_n597), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n593), .B1(new_n601), .B2(KEYINPUT15), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT15), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n596), .A2(G50gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n329), .A2(G43gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT87), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT87), .B1(new_n604), .B2(new_n605), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n608), .A2(new_n609), .A3(new_n593), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT7), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  INV_X1    g416(.A(G85gat), .ZN(new_n618));
  INV_X1    g417(.A(G92gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(KEYINPUT8), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G99gat), .B(G106gat), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(new_n623), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n614), .A2(new_n624), .B1(KEYINPUT41), .B2(new_n581), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT17), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n626), .A3(new_n612), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT90), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n611), .A2(KEYINPUT90), .A3(new_n626), .A4(new_n612), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n621), .B(new_n622), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n614), .B2(new_n626), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n625), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G190gat), .B(G218gat), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n586), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n585), .A3(new_n637), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n544), .A2(new_n545), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n548), .A2(new_n546), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n556), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n624), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n633), .B1(new_n549), .B2(new_n556), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n557), .A2(KEYINPUT10), .A3(new_n624), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n647), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n646), .B1(new_n652), .B2(new_n653), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  AOI21_X1  g461(.A(new_n645), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n662), .ZN(new_n665));
  NOR4_X1   g464(.A1(new_n657), .A2(KEYINPUT99), .A3(new_n658), .A4(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n657), .B2(new_n658), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n580), .A2(new_n644), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G113gat), .B(G141gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G197gat), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT11), .B(G169gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT12), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n571), .B1(new_n613), .B2(KEYINPUT17), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n631), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(G229gat), .A2(G233gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n572), .A2(new_n613), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n680), .A2(KEYINPUT18), .A3(new_n681), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n631), .B2(new_n679), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT92), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n686), .A2(new_n687), .A3(KEYINPUT18), .A4(new_n681), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n681), .B(KEYINPUT13), .Z(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n572), .A2(new_n613), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n683), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n686), .A2(new_n681), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n678), .B1(new_n689), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n689), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n678), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT93), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI211_X1 g499(.A(new_n693), .B(new_n677), .C1(new_n694), .C2(new_n695), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT93), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n689), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n697), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n672), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n529), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n513), .A2(new_n515), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n492), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT16), .B(G8gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT42), .Z(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(G8gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT100), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1325gat));
  INV_X1    g515(.A(new_n706), .ZN(new_n717));
  INV_X1    g516(.A(new_n327), .ZN(new_n718));
  OAI21_X1  g517(.A(G15gat), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n519), .A2(G15gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n717), .B2(new_n720), .ZN(G1326gat));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n409), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT101), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT43), .B(G22gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1327gat));
  AOI21_X1  g524(.A(new_n644), .B1(new_n518), .B2(new_n528), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n704), .A2(new_n580), .A3(new_n670), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n726), .A2(new_n591), .A3(new_n707), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT45), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n730), .B(new_n643), .C1(new_n517), .C2(new_n527), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n731), .A2(KEYINPUT102), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(KEYINPUT102), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n735), .B(new_n643), .C1(new_n517), .C2(new_n527), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(KEYINPUT44), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n733), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n738), .A2(new_n707), .A3(new_n727), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n729), .B1(new_n739), .B2(new_n591), .ZN(G1328gat));
  NAND3_X1  g539(.A1(new_n529), .A2(new_n643), .A3(new_n727), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n492), .A2(new_n587), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT46), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n734), .A2(KEYINPUT44), .A3(new_n736), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n731), .A2(KEYINPUT102), .A3(new_n732), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n745), .A2(new_n492), .A3(new_n746), .A4(new_n727), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G36gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT104), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n744), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1329gat));
  NAND4_X1  g552(.A1(new_n745), .A2(new_n327), .A3(new_n746), .A4(new_n727), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n596), .B1(new_n754), .B2(KEYINPUT106), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n738), .A2(new_n756), .A3(new_n327), .A4(new_n727), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n322), .A2(new_n596), .ZN(new_n760));
  OR3_X1    g559(.A1(new_n741), .A2(KEYINPUT105), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT105), .B1(new_n741), .B2(new_n760), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n754), .A2(G43gat), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n761), .A2(new_n762), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n759), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(G1330gat));
  NOR2_X1   g567(.A1(new_n410), .A2(new_n329), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n745), .A2(new_n746), .A3(new_n727), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n329), .B1(new_n741), .B2(new_n410), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g572(.A1(new_n704), .A2(new_n580), .A3(new_n644), .A4(new_n670), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n528), .B2(new_n518), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n707), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G57gat), .ZN(G1332gat));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n492), .B1(new_n778), .B2(new_n540), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT107), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n540), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1333gat));
  NAND2_X1  g582(.A1(new_n775), .A2(new_n327), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n519), .A2(G71gat), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n784), .A2(G71gat), .B1(new_n775), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g586(.A1(new_n775), .A2(new_n409), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G78gat), .ZN(G1335gat));
  INV_X1    g588(.A(new_n697), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n701), .A2(new_n702), .A3(new_n689), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n702), .B1(new_n701), .B2(new_n689), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(new_n580), .A3(new_n671), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n738), .A2(new_n707), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n580), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n726), .A2(KEYINPUT51), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT51), .B1(new_n726), .B2(new_n796), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n670), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n707), .A2(new_n618), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n795), .A2(new_n618), .B1(new_n799), .B2(new_n800), .ZN(G1336gat));
  NAND4_X1  g600(.A1(new_n745), .A2(new_n492), .A3(new_n746), .A4(new_n794), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G92gat), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n492), .A2(new_n619), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT52), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n803), .B(new_n807), .C1(new_n799), .C2(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1337gat));
  NAND4_X1  g608(.A1(new_n745), .A2(new_n327), .A3(new_n746), .A4(new_n794), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G99gat), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n519), .A2(G99gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n799), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT108), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT108), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n811), .B(new_n815), .C1(new_n799), .C2(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1338gat));
  NAND4_X1  g616(.A1(new_n745), .A2(new_n409), .A3(new_n746), .A4(new_n794), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G106gat), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n410), .A2(G106gat), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n670), .B(new_n820), .C1(new_n797), .C2(new_n798), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(KEYINPUT109), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT53), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n819), .B(new_n821), .C1(KEYINPUT109), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(G1339gat));
  NAND2_X1  g626(.A1(new_n322), .A2(new_n410), .ZN(new_n828));
  INV_X1    g627(.A(new_n580), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n657), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n655), .A2(new_n656), .A3(new_n647), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g632(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n834));
  AOI21_X1  g633(.A(new_n662), .B1(new_n657), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n836), .A2(new_n837), .B1(new_n663), .B2(new_n666), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n793), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n686), .B2(new_n681), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n683), .A2(new_n692), .A3(new_n691), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n686), .A2(new_n841), .A3(new_n681), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n676), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n670), .B(new_n846), .C1(new_n791), .C2(new_n792), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n643), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n791), .B2(new_n792), .ZN(new_n849));
  INV_X1    g648(.A(new_n838), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n836), .A2(new_n837), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n643), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n829), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n672), .A2(new_n793), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n828), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n513), .A2(new_n515), .A3(new_n492), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(G113gat), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n858), .A2(new_n859), .A3(new_n704), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n850), .A2(new_n851), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n847), .B1(new_n704), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n853), .B1(new_n862), .B2(new_n644), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n855), .B1(new_n863), .B2(new_n580), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n707), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n865), .A2(new_n509), .A3(new_n525), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n793), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n860), .B1(new_n867), .B2(new_n859), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n858), .A2(new_n869), .A3(new_n671), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n670), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n869), .ZN(G1341gat));
  NAND3_X1  g671(.A1(new_n866), .A2(new_n563), .A3(new_n580), .ZN(new_n873));
  OAI21_X1  g672(.A(G127gat), .B1(new_n858), .B2(new_n829), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT112), .Z(G1342gat));
  NOR2_X1   g675(.A1(new_n644), .A2(new_n492), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT113), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(G134gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n865), .A2(new_n525), .A3(new_n879), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n881));
  OAI21_X1  g680(.A(G134gat), .B1(new_n858), .B2(new_n644), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G1343gat));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n410), .B1(new_n854), .B2(new_n855), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT114), .B1(new_n886), .B2(KEYINPUT57), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n864), .A2(new_n409), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n892));
  INV_X1    g691(.A(new_n832), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(new_n657), .A3(new_n830), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n657), .A2(new_n834), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n665), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n892), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n835), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT116), .A4(new_n837), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n837), .A3(new_n898), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n838), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n793), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n643), .B1(new_n903), .B2(new_n847), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n829), .B1(new_n904), .B2(new_n853), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n410), .B1(new_n905), .B2(new_n855), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT57), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n887), .A2(new_n891), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n718), .A2(new_n857), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n704), .A2(new_n335), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n327), .A2(new_n410), .ZN(new_n913));
  AND4_X1   g712(.A1(new_n707), .A2(new_n864), .A3(new_n509), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G141gat), .B1(new_n914), .B2(new_n793), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n885), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT58), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n885), .B(new_n918), .C1(new_n912), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n908), .A2(new_n670), .A3(new_n910), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n336), .A2(KEYINPUT59), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n909), .A2(new_n671), .ZN(new_n924));
  AOI211_X1 g723(.A(new_n890), .B(new_n410), .C1(new_n854), .C2(new_n855), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n900), .A2(new_n901), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n850), .A3(new_n899), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n847), .B1(new_n927), .B2(new_n704), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n853), .B1(new_n928), .B2(new_n644), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n855), .B1(new_n929), .B2(new_n580), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT57), .B1(new_n930), .B2(new_n409), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n924), .B1(new_n925), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G148gat), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n922), .A2(new_n923), .B1(new_n933), .B2(KEYINPUT59), .ZN(new_n934));
  INV_X1    g733(.A(new_n914), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n935), .A2(G148gat), .A3(new_n671), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n921), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n936), .ZN(new_n938));
  INV_X1    g737(.A(new_n923), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT57), .B1(new_n864), .B2(new_n409), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n940), .A2(new_n889), .B1(new_n906), .B2(KEYINPUT57), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n909), .B1(new_n941), .B2(new_n887), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n939), .B1(new_n942), .B2(new_n670), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n944), .B1(new_n932), .B2(G148gat), .ZN(new_n945));
  OAI211_X1 g744(.A(KEYINPUT118), .B(new_n938), .C1(new_n943), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n937), .A2(new_n946), .ZN(G1345gat));
  NOR2_X1   g746(.A1(new_n935), .A2(new_n829), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n948), .A2(KEYINPUT119), .ZN(new_n949));
  AOI21_X1  g748(.A(G155gat), .B1(new_n948), .B2(KEYINPUT119), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n829), .A2(new_n533), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n949), .A2(new_n950), .B1(new_n942), .B2(new_n951), .ZN(G1346gat));
  NAND2_X1  g751(.A1(new_n942), .A2(new_n643), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT120), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n942), .A2(new_n955), .A3(new_n643), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n954), .A2(G162gat), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n878), .A2(G162gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n865), .A2(new_n913), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1347gat));
  NOR2_X1   g759(.A1(new_n707), .A2(new_n509), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n856), .A2(new_n961), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n962), .A2(new_n223), .A3(new_n704), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n961), .A2(new_n525), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n864), .A2(new_n793), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n963), .B1(new_n223), .B2(new_n965), .ZN(G1348gat));
  OAI21_X1  g765(.A(G176gat), .B1(new_n962), .B2(new_n671), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n864), .A2(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n670), .A2(new_n224), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(G1349gat));
  OAI21_X1  g769(.A(KEYINPUT121), .B1(new_n962), .B2(new_n829), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G183gat), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n962), .A2(KEYINPUT121), .A3(new_n829), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n580), .A2(new_n216), .ZN(new_n974));
  OAI22_X1  g773(.A1(new_n972), .A2(new_n973), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g775(.A1(new_n856), .A2(new_n643), .A3(new_n961), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n217), .B1(new_n978), .B2(KEYINPUT61), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n979), .B1(new_n977), .B2(new_n980), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n643), .A2(new_n217), .ZN(new_n983));
  OAI22_X1  g782(.A1(new_n981), .A2(new_n982), .B1(new_n968), .B2(new_n983), .ZN(G1351gat));
  NOR2_X1   g783(.A1(new_n925), .A2(new_n931), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT124), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n961), .A2(new_n718), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n989), .B1(new_n925), .B2(new_n931), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n986), .A2(new_n793), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(KEYINPUT125), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n990), .A2(new_n988), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT125), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n993), .A2(new_n994), .A3(new_n793), .A4(new_n986), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n992), .A2(new_n995), .A3(G197gat), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n886), .A2(new_n988), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n997), .A2(KEYINPUT123), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(KEYINPUT123), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(G197gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n1000), .A2(new_n1001), .A3(new_n793), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n996), .A2(new_n1002), .ZN(G1352gat));
  NAND2_X1  g802(.A1(new_n993), .A2(new_n986), .ZN(new_n1004));
  OAI21_X1  g803(.A(G204gat), .B1(new_n1004), .B2(new_n671), .ZN(new_n1005));
  AOI21_X1  g804(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n1006));
  NAND4_X1  g805(.A1(new_n886), .A2(new_n670), .A3(new_n988), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g806(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1005), .A2(new_n1009), .ZN(G1353gat));
  NAND4_X1  g809(.A1(new_n998), .A2(new_n359), .A3(new_n999), .A4(new_n580), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1011), .B(KEYINPUT127), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n988), .A2(new_n580), .ZN(new_n1013));
  OAI21_X1  g812(.A(G211gat), .B1(new_n985), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g813(.A1(new_n1014), .A2(KEYINPUT63), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1014), .A2(KEYINPUT63), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(G1354gat));
  NOR3_X1   g816(.A1(new_n1004), .A2(new_n360), .A3(new_n644), .ZN(new_n1018));
  AOI21_X1  g817(.A(G218gat), .B1(new_n1000), .B2(new_n643), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n1018), .A2(new_n1019), .ZN(G1355gat));
endmodule


