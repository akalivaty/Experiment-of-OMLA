//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n461));
  AND2_X1   g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G125), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n465), .A2(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g050(.A(KEYINPUT65), .B(G2105), .C1(new_n475), .C2(new_n462), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n469), .A2(new_n465), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n470), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(new_n463), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n465), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(new_n465), .A3(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n469), .A2(KEYINPUT66), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n491), .A2(new_n465), .A3(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n463), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n490), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT67), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  INV_X1    g082(.A(G75), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(new_n502), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n503), .A2(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n502), .B1(new_n511), .B2(new_n512), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n517), .B1(new_n514), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n510), .B1(new_n518), .B2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(G51), .B2(new_n515), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT5), .B1(new_n504), .B2(G543), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n503), .A2(KEYINPUT69), .A3(new_n505), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n528), .A2(G63), .A3(G651), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n513), .A2(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n524), .A2(new_n530), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(new_n528), .A2(new_n529), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n513), .A2(G90), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n515), .A2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n538), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n534), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n513), .A2(G81), .B1(new_n515), .B2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(new_n512), .ZN(new_n556));
  NOR2_X1   g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n511), .A2(new_n512), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n560), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n503), .B2(new_n505), .ZN(new_n565));
  AND2_X1   g140(.A1(G78), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n513), .A2(G91), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT70), .ZN(G299));
  AOI22_X1  g145(.A1(new_n513), .A2(G87), .B1(new_n515), .B2(G49), .ZN(new_n571));
  AOI21_X1  g146(.A(G74), .B1(new_n528), .B2(new_n529), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n537), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g150(.A(KEYINPUT71), .B(new_n571), .C1(new_n572), .C2(new_n537), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n513), .A2(G86), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n515), .A2(new_n581), .A3(G48), .ZN(new_n582));
  OAI211_X1 g157(.A(G48), .B(G543), .C1(new_n556), .C2(new_n557), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT73), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n506), .B2(G61), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n537), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n513), .A2(KEYINPUT72), .A3(G86), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(G305));
  AND2_X1   g167(.A1(new_n535), .A2(G60), .ZN(new_n593));
  AND2_X1   g168(.A1(G72), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n513), .A2(G85), .B1(new_n515), .B2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(new_n515), .A2(G54), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n537), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT74), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n513), .A2(G92), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT10), .Z(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G321));
  XNOR2_X1  g183(.A(G321), .B(KEYINPUT75), .ZN(G284));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G860), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n605), .B1(G559), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT76), .ZN(G148));
  NAND2_X1  g191(.A1(new_n549), .A2(new_n606), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n605), .A2(G559), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n617), .B1(new_n619), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n463), .A2(new_n471), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n479), .A2(G123), .ZN(new_n628));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(G135), .B2(new_n470), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(G156));
  XOR2_X1   g209(.A(KEYINPUT15), .B(G2435), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2430), .Z(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT78), .B(KEYINPUT14), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(G14), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n646), .ZN(G401));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT79), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NOR2_X1   g231(.A1(G2072), .A2(G2078), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n655), .B(new_n656), .C1(new_n442), .C2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(KEYINPUT80), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n442), .A2(new_n657), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(KEYINPUT17), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n662), .B(new_n654), .C1(new_n660), .C2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n655), .A2(new_n660), .A3(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n659), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  AOI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n670), .C2(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT81), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(G229));
  MUX2_X1   g262(.A(G6), .B(G305), .S(G16), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT32), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  MUX2_X1   g265(.A(G23), .B(new_n573), .S(G16), .Z(new_n691));
  XOR2_X1   g266(.A(KEYINPUT33), .B(G1976), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT83), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT82), .B(KEYINPUT34), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n694), .A2(new_n702), .A3(new_n700), .ZN(new_n705));
  MUX2_X1   g280(.A(G24), .B(G290), .S(G16), .Z(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(G1986), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(G1986), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n479), .A2(G119), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n470), .A2(G131), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n465), .A2(G107), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G25), .B(new_n713), .S(G29), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT35), .B(G1991), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n707), .A2(new_n708), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n704), .A2(new_n705), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT36), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n704), .A2(new_n721), .A3(new_n705), .A4(new_n718), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G32), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n470), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n471), .A2(G105), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT26), .Z(new_n730));
  INV_X1    g305(.A(G129), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n486), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n725), .B1(new_n734), .B2(new_n724), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT27), .B(G1996), .Z(new_n736));
  NAND2_X1  g311(.A1(G160), .A2(G29), .ZN(new_n737));
  INV_X1    g312(.A(G34), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT24), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(KEYINPUT24), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(KEYINPUT87), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(KEYINPUT87), .B2(new_n740), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G2084), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n735), .A2(new_n736), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n695), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n695), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT92), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n745), .B1(new_n748), .B2(G1961), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT93), .Z(new_n750));
  NAND2_X1  g325(.A1(G168), .A2(G16), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n751), .B(KEYINPUT88), .C1(G16), .C2(G21), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(KEYINPUT88), .B2(new_n751), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT89), .B(G1966), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G19), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n550), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1341), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT90), .ZN(new_n761));
  INV_X1    g336(.A(G28), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n762), .B2(KEYINPUT30), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(KEYINPUT30), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n632), .A2(G29), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n768), .B1(new_n767), .B2(new_n766), .C1(new_n735), .C2(new_n736), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n724), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n724), .ZN(new_n772));
  INV_X1    g347(.A(G2090), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n769), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n775), .B1(new_n744), .B2(new_n743), .C1(new_n770), .C2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(G115), .A2(G2104), .ZN(new_n777));
  INV_X1    g352(.A(G127), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n469), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n465), .B1(new_n779), .B2(KEYINPUT86), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(KEYINPUT86), .B2(new_n779), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n470), .A2(G139), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT25), .Z(new_n784));
  NAND3_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G33), .B(new_n785), .S(G29), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2072), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n724), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n479), .A2(G128), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n470), .A2(G140), .ZN(new_n792));
  OR2_X1    g367(.A1(G104), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(new_n724), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT85), .B(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G27), .A2(G29), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G164), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2078), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n776), .A2(new_n787), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n695), .A2(G20), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT95), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT23), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n611), .B2(new_n695), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1956), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n695), .A2(G4), .ZN(new_n809));
  INV_X1    g384(.A(new_n605), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n695), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1348), .ZN(new_n812));
  AOI211_X1 g387(.A(new_n808), .B(new_n812), .C1(G1961), .C2(new_n748), .ZN(new_n813));
  AND4_X1   g388(.A1(new_n750), .A2(new_n759), .A3(new_n803), .A4(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n723), .A2(KEYINPUT96), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(KEYINPUT96), .B1(new_n723), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(G311));
  NAND2_X1  g392(.A1(new_n723), .A2(new_n814), .ZN(G150));
  XNOR2_X1  g393(.A(KEYINPUT98), .B(G93), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n513), .A2(new_n819), .B1(new_n515), .B2(G55), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  INV_X1    g397(.A(G67), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n534), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n537), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n821), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT100), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n828), .A2(KEYINPUT100), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(new_n614), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n810), .A2(G559), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT38), .Z(new_n836));
  NOR3_X1   g411(.A1(new_n830), .A2(new_n831), .A3(new_n550), .ZN(new_n837));
  OR3_X1    g412(.A1(new_n828), .A2(KEYINPUT99), .A3(new_n549), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT99), .B1(new_n828), .B2(new_n549), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n836), .B(new_n841), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n614), .B1(new_n843), .B2(KEYINPUT39), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n834), .B1(new_n844), .B2(new_n845), .ZN(G145));
  OAI21_X1  g421(.A(KEYINPUT66), .B1(new_n469), .B2(new_n492), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n463), .A2(new_n495), .A3(new_n494), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n499), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n488), .A2(new_n489), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n479), .B2(G126), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n795), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n734), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n785), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n479), .A2(G130), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n470), .A2(G142), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n465), .A2(G118), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n856), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(new_n623), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n713), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT102), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n862), .B(KEYINPUT102), .Z(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n855), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n632), .B(new_n484), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT101), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G160), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n866), .A2(new_n869), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n870), .A2(new_n871), .A3(G37), .ZN(new_n872));
  XNOR2_X1  g447(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(G395));
  XNOR2_X1  g449(.A(new_n841), .B(new_n619), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n810), .A2(G299), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n611), .A2(new_n605), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT104), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(KEYINPUT105), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n876), .A2(new_n877), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n875), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n884), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(G290), .B(G305), .Z(new_n889));
  XOR2_X1   g464(.A(G303), .B(new_n573), .Z(new_n890));
  XOR2_X1   g465(.A(new_n889), .B(new_n890), .Z(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT42), .Z(new_n892));
  AND2_X1   g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n888), .A2(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(G868), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(G868), .B2(new_n832), .ZN(G295));
  OAI21_X1  g471(.A(new_n895), .B1(G868), .B2(new_n832), .ZN(G331));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n898));
  OAI21_X1  g473(.A(G171), .B1(new_n837), .B2(new_n840), .ZN(new_n899));
  INV_X1    g474(.A(new_n831), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n549), .A3(new_n829), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n901), .A2(G301), .A3(new_n838), .A4(new_n839), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n902), .A3(G168), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(G168), .B1(new_n899), .B2(new_n902), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n878), .A2(new_n879), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  OAI22_X1  g483(.A1(new_n904), .A2(new_n905), .B1(new_n908), .B2(new_n881), .ZN(new_n909));
  INV_X1    g484(.A(new_n905), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n878), .A3(new_n903), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n912), .B2(new_n891), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(KEYINPUT106), .ZN(new_n914));
  INV_X1    g489(.A(new_n891), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n882), .B1(new_n904), .B2(new_n905), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n910), .A2(new_n917), .A3(new_n878), .A4(new_n903), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n911), .A2(KEYINPUT106), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n916), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n891), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .A4(new_n919), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n898), .B1(new_n921), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n926), .A3(new_n919), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n919), .A2(new_n925), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n929), .A2(KEYINPUT43), .B1(new_n930), .B2(new_n913), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n898), .B2(new_n931), .ZN(G397));
  INV_X1    g507(.A(KEYINPUT126), .ZN(new_n933));
  NOR2_X1   g508(.A1(G290), .A2(G1986), .ZN(new_n934));
  AOI21_X1  g509(.A(G1384), .B1(new_n849), .B2(new_n851), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT108), .B(G40), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n476), .A2(new_n466), .A3(new_n472), .A4(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(G1986), .A3(G290), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT109), .Z(new_n945));
  XNOR2_X1  g520(.A(new_n795), .B(G2067), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT110), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n733), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n941), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT111), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n713), .A2(new_n716), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n716), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n941), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n945), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(G164), .B2(G1384), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n935), .A2(KEYINPUT112), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n940), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(new_n936), .B2(KEYINPUT50), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n957), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n563), .A2(new_n567), .A3(KEYINPUT57), .A4(new_n568), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT118), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT116), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n563), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n559), .A2(new_n562), .A3(KEYINPUT116), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(new_n567), .A3(new_n568), .A4(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT117), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT57), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n971), .B2(new_n973), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n967), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n940), .B1(KEYINPUT45), .B2(new_n935), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT56), .B(G2072), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n938), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n965), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT119), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT112), .B1(new_n852), .B2(new_n982), .ZN(new_n983));
  AOI211_X1 g558(.A(new_n959), .B(G1384), .C1(new_n849), .C2(new_n851), .ZN(new_n984));
  NOR4_X1   g559(.A1(new_n983), .A2(new_n984), .A3(G2067), .A4(new_n940), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n960), .A2(new_n958), .A3(new_n961), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n935), .A2(new_n958), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n963), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1348), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n981), .B1(new_n991), .B2(new_n605), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n966), .B(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n971), .A2(new_n973), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT117), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT50), .B1(new_n983), .B2(new_n984), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n940), .B1(new_n958), .B2(new_n935), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1956), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n979), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n992), .A2(new_n1003), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n991), .A2(new_n981), .A3(new_n605), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n980), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT61), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n976), .B1(new_n965), .B2(new_n979), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n980), .A3(KEYINPUT61), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n977), .A2(new_n948), .A3(new_n938), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT120), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n977), .A2(new_n938), .A3(new_n1015), .A4(new_n948), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n960), .A2(new_n963), .A3(new_n961), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT58), .B(G1341), .Z(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1012), .B1(new_n1020), .B2(new_n550), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1020), .A2(new_n1012), .A3(new_n550), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1010), .B(new_n1011), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n989), .A2(new_n990), .ZN(new_n1024));
  INV_X1    g599(.A(new_n985), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT60), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n810), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n991), .A2(KEYINPUT60), .A3(new_n605), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1028), .A2(new_n1029), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1006), .B1(new_n1023), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n937), .B1(new_n983), .B2(new_n984), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n1034));
  INV_X1    g609(.A(G2078), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n977), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1036), .A2(KEYINPUT53), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1035), .A3(new_n977), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT121), .ZN(new_n1039));
  INV_X1    g614(.A(G1961), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1037), .A2(new_n1039), .B1(new_n1040), .B2(new_n989), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n977), .A2(new_n1035), .A3(new_n938), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(G301), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n989), .A2(new_n1040), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n935), .A2(KEYINPUT45), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n472), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n472), .A2(new_n1051), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n464), .A2(new_n465), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1035), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n938), .A2(new_n1050), .A3(new_n1052), .A4(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1049), .A2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1047), .A2(G301), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1032), .B1(new_n1048), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1033), .A2(new_n977), .ZN(new_n1061));
  INV_X1    g636(.A(G1966), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n986), .A2(new_n744), .A3(new_n963), .A4(new_n988), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(G168), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G8), .ZN(new_n1066));
  AOI21_X1  g641(.A(G168), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT51), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1065), .A2(new_n1069), .A3(G8), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n999), .A2(new_n773), .A3(new_n1000), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1050), .A2(new_n963), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n935), .A2(KEYINPUT45), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n698), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  AND2_X1   g652(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1078));
  NOR2_X1   g653(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(G303), .B2(G8), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(G303), .B(G8), .C1(KEYINPUT113), .C2(KEYINPUT55), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1077), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G8), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n983), .A2(new_n984), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n963), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT49), .ZN(new_n1090));
  INV_X1    g665(.A(G1981), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n589), .A2(new_n537), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n581), .B1(new_n515), .B2(G48), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n583), .A2(KEYINPUT73), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n578), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n582), .A2(new_n584), .B1(G86), .B2(new_n513), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT115), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1091), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n590), .A2(new_n591), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1101), .A2(new_n586), .A3(G1981), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1090), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n590), .B1(new_n1098), .B2(KEYINPUT115), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1105));
  OAI21_X1  g680(.A(G1981), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n587), .A2(new_n1091), .A3(new_n590), .A4(new_n591), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT49), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1089), .A2(new_n1103), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1976), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n575), .A2(new_n1110), .A3(new_n576), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n573), .A2(new_n1110), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1089), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1017), .A2(G8), .A3(new_n1114), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT52), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1109), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(G1971), .B1(new_n977), .B2(new_n938), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n987), .B1(new_n1088), .B2(new_n958), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n940), .A2(G2090), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G303), .A2(G8), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(new_n1079), .ZN(new_n1124));
  OAI21_X1  g699(.A(G8), .B1(new_n1124), .B2(new_n1081), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1122), .A2(KEYINPUT114), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n986), .A2(new_n988), .A3(new_n1121), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1075), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1087), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1086), .B(new_n1118), .C1(new_n1126), .C2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1041), .A2(G301), .A3(new_n1047), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1049), .B(new_n1057), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1032), .B1(new_n1134), .B2(G171), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1132), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1031), .A2(new_n1060), .A3(new_n1071), .A4(new_n1136), .ZN(new_n1137));
  AOI211_X1 g712(.A(G1976), .B(G288), .C1(new_n1103), .C2(new_n1108), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1089), .B1(new_n1138), .B2(new_n1102), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1140));
  AOI21_X1  g715(.A(G286), .B1(new_n1122), .B2(new_n1085), .ZN(new_n1141));
  AND4_X1   g716(.A1(G8), .A2(new_n1118), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1109), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G286), .A2(KEYINPUT63), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1086), .A2(G8), .A3(new_n1140), .A4(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT114), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1129), .A2(new_n1130), .A3(new_n1127), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1145), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1144), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1137), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1068), .A2(new_n1154), .A3(new_n1070), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1132), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(new_n1156), .A3(new_n1048), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1155), .A2(new_n1156), .A3(KEYINPUT125), .A4(new_n1048), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1071), .A2(KEYINPUT62), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1153), .A2(KEYINPUT124), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1137), .A2(new_n1164), .A3(new_n1152), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n956), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n952), .A2(new_n954), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(G2067), .B2(new_n795), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1168), .A2(new_n941), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n941), .A2(new_n948), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT46), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n734), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n941), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT47), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n952), .A2(new_n955), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n942), .B(KEYINPUT48), .Z(new_n1177));
  OAI21_X1  g752(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1169), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n933), .B1(new_n1166), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1165), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1164), .B1(new_n1137), .B2(new_n1152), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1159), .A2(new_n1161), .A3(new_n1160), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OAI211_X1 g760(.A(KEYINPUT126), .B(new_n1179), .C1(new_n1185), .C2(new_n956), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1181), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(G319), .ZN(new_n1189));
  NOR3_X1   g763(.A1(G401), .A2(G227), .A3(new_n1189), .ZN(new_n1190));
  OR2_X1    g764(.A1(new_n1190), .A2(KEYINPUT127), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1190), .A2(KEYINPUT127), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n1191), .B(new_n1192), .C1(new_n685), .C2(new_n686), .ZN(new_n1193));
  OR2_X1    g767(.A1(new_n1193), .A2(new_n872), .ZN(new_n1194));
  NOR2_X1   g768(.A1(new_n931), .A2(new_n1194), .ZN(G308));
  OR2_X1    g769(.A1(new_n931), .A2(new_n1194), .ZN(G225));
endmodule


