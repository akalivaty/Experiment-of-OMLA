//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT81), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  OAI21_X1  g003(.A(G221), .B1(new_n189), .B2(G902), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT64), .A2(G143), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(G143), .ZN(new_n193));
  OAI21_X1  g007(.A(G146), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n194), .A2(new_n195), .A3(G128), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT64), .A2(G143), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n196), .A3(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n199), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(new_n197), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n203), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n198), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G107), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n210), .A2(G107), .ZN(new_n213));
  OAI21_X1  g027(.A(G101), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G104), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n219), .A4(new_n211), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n209), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT84), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n209), .A2(KEYINPUT84), .A3(new_n221), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n196), .A2(G143), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n192), .A2(new_n193), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n196), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G128), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n227), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n204), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(new_n231), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n233), .A2(new_n198), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n226), .B1(new_n238), .B2(new_n221), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(G137), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT11), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n240), .B(new_n245), .C1(new_n241), .C2(G137), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n243), .A2(new_n249), .A3(new_n244), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n239), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT12), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n239), .A2(KEYINPUT12), .A3(new_n251), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT10), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n229), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n208), .A2(new_n258), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT83), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n220), .A2(new_n263), .A3(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n215), .A2(new_n218), .A3(new_n211), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n264), .B(new_n266), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n226), .A2(new_n257), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n251), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n238), .A2(KEYINPUT68), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n233), .A2(new_n271), .A3(new_n198), .A4(new_n237), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT10), .A3(new_n221), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n256), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(G110), .B(G140), .Z(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT82), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G227), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n278), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n275), .A2(new_n281), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT85), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n268), .A2(new_n274), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n251), .ZN(new_n287));
  AOI211_X1 g101(.A(KEYINPUT85), .B(new_n269), .C1(new_n268), .C2(new_n274), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(G469), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT86), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n254), .B2(new_n255), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n254), .A2(new_n292), .A3(new_n255), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n284), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n275), .B1(new_n287), .B2(new_n288), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n282), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G469), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n291), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(G469), .A2(G902), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n191), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT96), .ZN(new_n304));
  XNOR2_X1  g118(.A(G116), .B(G122), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n307), .A2(new_n217), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n308), .A2(KEYINPUT95), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n199), .A2(G143), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n228), .B2(new_n199), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(G134), .ZN(new_n312));
  INV_X1    g126(.A(G116), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT14), .A3(G122), .ZN(new_n314));
  INV_X1    g128(.A(new_n305), .ZN(new_n315));
  OAI211_X1 g129(.A(G107), .B(new_n314), .C1(new_n315), .C2(KEYINPUT14), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n308), .A2(KEYINPUT95), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n309), .A2(new_n312), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT13), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n207), .A2(new_n319), .A3(G128), .ZN(new_n320));
  OAI211_X1 g134(.A(G134), .B(new_n320), .C1(new_n311), .C2(new_n319), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n307), .A2(new_n217), .ZN(new_n322));
  OAI221_X1 g136(.A(new_n321), .B1(G134), .B2(new_n311), .C1(new_n308), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G217), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n189), .A2(new_n325), .A3(G953), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n318), .A2(new_n323), .A3(new_n326), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G902), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT15), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G478), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n332), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  XNOR2_X1  g152(.A(G125), .B(G140), .ZN(new_n339));
  MUX2_X1   g153(.A(new_n338), .B(new_n339), .S(KEYINPUT16), .Z(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(G146), .ZN(new_n341));
  INV_X1    g155(.A(G237), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n279), .A3(G214), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n228), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(G143), .B2(new_n343), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(new_n249), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT17), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n249), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n341), .B(new_n347), .C1(new_n348), .C2(KEYINPUT17), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(KEYINPUT18), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT18), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n345), .B1(new_n351), .B2(new_n249), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT90), .B1(new_n339), .B2(new_n196), .ZN(new_n353));
  INV_X1    g167(.A(new_n339), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(G146), .B2(new_n354), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n339), .A2(KEYINPUT90), .A3(new_n196), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n350), .B(new_n352), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(G113), .B(G122), .Z(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT91), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(new_n210), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n358), .A2(new_n361), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n331), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT93), .B(G475), .Z(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n340), .A2(new_n196), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n339), .B(KEYINPUT19), .Z(new_n369));
  OAI211_X1 g183(.A(new_n348), .B(new_n368), .C1(G146), .C2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n370), .A2(new_n357), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n371), .A2(new_n361), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n362), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n374));
  NOR2_X1   g188(.A1(G475), .A2(G902), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT92), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n374), .B1(new_n373), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n367), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n336), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G214), .B1(G237), .B2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(G234), .A2(G237), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n385), .A2(G952), .A3(new_n279), .ZN(new_n386));
  XOR2_X1   g200(.A(KEYINPUT21), .B(G898), .Z(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n385), .A2(G902), .A3(G953), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT87), .B1(new_n262), .B2(new_n337), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n392), .B(G125), .C1(new_n260), .C2(new_n261), .ZN(new_n393));
  AOI221_X4 g207(.A(KEYINPUT67), .B1(new_n230), .B2(G128), .C1(new_n204), .C2(new_n234), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n236), .B1(new_n235), .B2(new_n231), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n337), .A3(new_n198), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G224), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G953), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT7), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(G116), .B(G119), .Z(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT2), .B(G113), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n267), .A2(new_n406), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n409));
  INV_X1    g223(.A(G119), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(G116), .ZN(new_n411));
  OAI211_X1 g225(.A(G113), .B(new_n411), .C1(new_n404), .C2(new_n409), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n221), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  XOR2_X1   g227(.A(G110), .B(G122), .Z(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n403), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n401), .A2(KEYINPUT88), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n391), .A2(new_n393), .A3(new_n397), .A4(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT7), .B1(new_n401), .B2(KEYINPUT88), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n412), .A2(new_n408), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(new_n221), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n414), .B(KEYINPUT8), .ZN(new_n423));
  OAI22_X1  g237(.A1(new_n419), .A2(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n331), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n398), .B(new_n400), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n407), .A2(new_n413), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n414), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n414), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n428), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT89), .B(new_n331), .C1(new_n417), .C2(new_n424), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G210), .B1(G237), .B2(G902), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n427), .A2(new_n437), .A3(new_n434), .A4(new_n435), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n384), .B(new_n390), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n303), .A2(new_n304), .A3(new_n382), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n296), .A2(new_n298), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n300), .A3(new_n331), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n302), .A3(new_n290), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n445), .A2(new_n441), .A3(new_n382), .A4(new_n190), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT96), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n262), .A2(new_n251), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT69), .ZN(new_n451));
  INV_X1    g265(.A(new_n244), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n241), .A2(G137), .ZN(new_n453));
  OAI21_X1  g267(.A(G131), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n250), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n451), .B1(new_n273), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n250), .A2(new_n454), .ZN(new_n457));
  AOI211_X1 g271(.A(KEYINPUT69), .B(new_n457), .C1(new_n270), .C2(new_n272), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT30), .B(new_n450), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n406), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT66), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n457), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n238), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n450), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n449), .A2(new_n406), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n456), .B2(new_n458), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(G101), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n342), .A2(new_n279), .A3(G210), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(KEYINPUT72), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT72), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n271), .B1(new_n396), .B2(new_n198), .ZN(new_n478));
  INV_X1    g292(.A(new_n272), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n455), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT69), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n273), .A2(new_n451), .A3(new_n455), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n459), .A2(new_n466), .B1(new_n483), .B2(new_n468), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n477), .B1(new_n484), .B2(new_n474), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n476), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT73), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT28), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n464), .A2(new_n406), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n469), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT28), .B1(new_n468), .B2(new_n480), .ZN(new_n492));
  OR3_X1    g306(.A1(new_n491), .A2(new_n475), .A3(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT74), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n483), .A2(new_n495), .A3(new_n468), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n450), .B1(new_n456), .B2(new_n458), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n406), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n469), .A2(KEYINPUT74), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n492), .B1(new_n500), .B2(KEYINPUT28), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n475), .A2(new_n488), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n493), .A2(new_n476), .A3(new_n485), .A4(new_n488), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT73), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n494), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G472), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT32), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT71), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT31), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n449), .B1(new_n238), .B2(new_n462), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n406), .B1(new_n511), .B2(KEYINPUT30), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n449), .B1(new_n481), .B2(new_n482), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(KEYINPUT30), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n469), .A2(new_n474), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT70), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n475), .B1(new_n483), .B2(new_n468), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n467), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n510), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n475), .B1(new_n491), .B2(new_n492), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n467), .A3(new_n510), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n509), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n517), .A2(new_n467), .A3(new_n518), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n518), .B1(new_n517), .B2(new_n467), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT31), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n521), .A2(new_n522), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT71), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G472), .A2(G902), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n508), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  AOI211_X1 g347(.A(KEYINPUT32), .B(new_n533), .C1(new_n524), .C2(new_n529), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n507), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT75), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT75), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n537), .B(new_n507), .C1(new_n532), .C2(new_n534), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT78), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT25), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT76), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n410), .B2(G128), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n199), .A2(KEYINPUT76), .A3(G119), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n542), .A2(new_n543), .B1(new_n410), .B2(G128), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT24), .B(G110), .Z(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT77), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n410), .B2(G128), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n410), .A2(G128), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(G110), .ZN(new_n553));
  OAI221_X1 g367(.A(new_n368), .B1(G146), .B2(new_n354), .C1(new_n547), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n544), .A2(new_n545), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  INV_X1    g370(.A(new_n552), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n554), .B1(new_n341), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT22), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G137), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n559), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n539), .B(new_n540), .C1(new_n564), .C2(G902), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n563), .B(new_n331), .C1(KEYINPUT78), .C2(KEYINPUT25), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n565), .B(new_n566), .C1(new_n539), .C2(new_n540), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n325), .B1(G234), .B2(new_n331), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(G902), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT79), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT80), .Z(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n448), .A2(new_n536), .A3(new_n538), .A4(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  NOR3_X1   g391(.A1(new_n520), .A2(new_n509), .A3(new_n523), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT71), .B1(new_n527), .B2(new_n528), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n331), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n580), .A2(G472), .B1(new_n531), .B2(new_n530), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n574), .A2(new_n191), .ZN(new_n582));
  INV_X1    g396(.A(new_n441), .ZN(new_n583));
  INV_X1    g397(.A(new_n381), .ZN(new_n584));
  AOI21_X1  g398(.A(G478), .B1(new_n330), .B2(new_n331), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT97), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n586), .A2(KEYINPUT97), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n330), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n328), .A2(KEYINPUT97), .A3(new_n586), .A4(new_n329), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n585), .B1(new_n591), .B2(G478), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n583), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n581), .A2(new_n445), .A3(new_n582), .A4(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT34), .B(G104), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G6));
  NAND3_X1  g412(.A1(new_n581), .A2(new_n445), .A3(new_n582), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n441), .A2(new_n336), .A3(new_n584), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G107), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT98), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n601), .B(new_n603), .ZN(G9));
  INV_X1    g418(.A(new_n562), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(KEYINPUT36), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n559), .B(new_n606), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n567), .A2(new_n568), .B1(new_n571), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n442), .A2(new_n447), .A3(new_n581), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT37), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n556), .ZN(G12));
  INV_X1    g426(.A(new_n303), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n384), .B1(new_n439), .B2(new_n440), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G900), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n389), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n386), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n381), .A2(new_n335), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR4_X1   g436(.A1(new_n613), .A2(new_n608), .A3(new_n615), .A4(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n536), .A3(new_n538), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G128), .ZN(G30));
  XOR2_X1   g439(.A(new_n619), .B(KEYINPUT39), .Z(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n303), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n608), .B1(new_n628), .B2(KEYINPUT40), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(KEYINPUT40), .B2(new_n628), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n532), .A2(new_n534), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n500), .A2(new_n475), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT99), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n516), .A2(new_n519), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n331), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n439), .A2(new_n440), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT38), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n584), .A2(new_n335), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n640), .A2(new_n383), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n630), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n228), .ZN(G45));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n584), .A2(new_n592), .A3(new_n620), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n645), .B1(new_n647), .B2(new_n615), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n614), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n649), .A2(new_n303), .A3(new_n609), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n536), .A2(new_n538), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G146), .ZN(G48));
  INV_X1    g466(.A(new_n295), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n293), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n654), .A2(new_n284), .B1(new_n297), .B2(new_n282), .ZN(new_n655));
  OAI21_X1  g469(.A(G469), .B1(new_n655), .B2(G902), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n190), .A3(new_n444), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n656), .A2(KEYINPUT101), .A3(new_n190), .A4(new_n444), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n536), .A2(new_n538), .A3(new_n575), .A4(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n595), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT41), .B(G113), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G15));
  NOR2_X1   g480(.A1(new_n662), .A2(new_n600), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n313), .ZN(G18));
  INV_X1    g482(.A(new_n390), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n614), .A2(new_n659), .A3(new_n669), .A4(new_n660), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n608), .A2(new_n336), .A3(new_n381), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n536), .A2(new_n538), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G119), .ZN(G21));
  NAND2_X1  g487(.A1(new_n500), .A2(KEYINPUT28), .ZN(new_n674));
  INV_X1    g488(.A(new_n492), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n474), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT102), .B1(new_n676), .B2(new_n520), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n527), .B(new_n678), .C1(new_n474), .C2(new_n501), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n677), .A2(new_n679), .A3(new_n522), .ZN(new_n680));
  AOI22_X1  g494(.A1(G472), .A2(new_n580), .B1(new_n680), .B2(new_n531), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n681), .A2(new_n575), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n670), .A3(new_n641), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  AND4_X1   g498(.A1(new_n614), .A2(new_n659), .A3(new_n646), .A4(new_n660), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n681), .B2(new_n609), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n580), .A2(G472), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n680), .A2(new_n531), .ZN(new_n689));
  AND4_X1   g503(.A1(new_n686), .A2(new_n688), .A3(new_n609), .A4(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n685), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G125), .ZN(G27));
  NAND3_X1  g506(.A1(new_n439), .A2(new_n383), .A3(new_n440), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n646), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n613), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n535), .A3(new_n575), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT42), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n613), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n536), .A2(new_n538), .A3(new_n575), .A4(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n647), .A2(KEYINPUT42), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n700), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n249), .ZN(G33));
  AND4_X1   g521(.A1(new_n536), .A2(new_n538), .A3(new_n575), .A4(new_n702), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n621), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT105), .B1(new_n703), .B2(new_n622), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G134), .ZN(G36));
  NAND2_X1  g527(.A1(new_n283), .A2(new_n289), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT45), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT46), .B1(new_n716), .B2(new_n302), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n300), .B2(new_n299), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n716), .A2(KEYINPUT46), .A3(new_n302), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n191), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n627), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n592), .A2(new_n381), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT43), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n724), .B1(new_n592), .B2(new_n381), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  OR3_X1    g541(.A1(new_n581), .A2(new_n727), .A3(new_n608), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n721), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n701), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n728), .A2(new_n729), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n733), .A2(KEYINPUT106), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(KEYINPUT106), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n731), .B(new_n732), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G137), .ZN(G39));
  XNOR2_X1  g551(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n720), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n720), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n697), .B1(new_n536), .B2(new_n538), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n574), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G140), .ZN(G42));
  INV_X1    g559(.A(new_n638), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n656), .A2(new_n444), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n722), .B1(new_n747), .B2(KEYINPUT49), .ZN(new_n748));
  AOI211_X1 g562(.A(new_n384), .B(new_n748), .C1(KEYINPUT49), .C2(new_n747), .ZN(new_n749));
  INV_X1    g563(.A(new_n640), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n746), .A2(new_n749), .A3(new_n582), .A4(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n661), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n701), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n746), .A3(new_n575), .A4(new_n386), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT113), .ZN(new_n755));
  INV_X1    g569(.A(new_n592), .ZN(new_n756));
  OR3_X1    g570(.A1(new_n755), .A2(new_n381), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n727), .A2(new_n618), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n690), .B2(new_n687), .ZN(new_n760));
  XOR2_X1   g574(.A(new_n760), .B(KEYINPUT112), .Z(new_n761));
  NAND2_X1  g575(.A1(new_n682), .A2(new_n758), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n747), .A2(new_n190), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n732), .B(new_n763), .C1(new_n742), .C2(new_n764), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n762), .A2(new_n383), .A3(new_n640), .A4(new_n752), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT50), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n757), .A2(new_n761), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n768), .B(new_n771), .Z(new_n772));
  NOR2_X1   g586(.A1(new_n755), .A2(new_n594), .ZN(new_n773));
  INV_X1    g587(.A(G952), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n762), .A2(new_n615), .A3(new_n752), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n773), .A2(new_n774), .A3(G953), .A4(new_n775), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n776), .A2(KEYINPUT115), .B1(new_n769), .B2(new_n770), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n778));
  INV_X1    g592(.A(new_n651), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n691), .A2(new_n624), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n691), .A2(new_n624), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n779), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n641), .A2(new_n614), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n190), .A2(new_n608), .A3(new_n445), .A4(new_n619), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n785), .B1(new_n786), .B2(KEYINPUT111), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n303), .A2(new_n608), .A3(new_n619), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n638), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT52), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n651), .A2(new_n691), .A3(new_n791), .A4(new_n624), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n784), .A2(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n593), .B1(new_n687), .B2(new_n690), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n536), .A2(new_n538), .A3(new_n671), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n620), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n706), .B1(new_n702), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n683), .B1(new_n662), .B2(new_n663), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n672), .B1(new_n662), .B2(new_n600), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n584), .B2(new_n336), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n381), .A2(KEYINPUT108), .A3(new_n335), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT109), .B1(new_n807), .B2(new_n441), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n807), .A2(KEYINPUT109), .A3(new_n441), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n599), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n610), .A2(new_n596), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n576), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n800), .A2(new_n712), .A3(new_n803), .A4(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n778), .B1(new_n796), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n802), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n682), .A2(new_n641), .A3(new_n670), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n536), .A2(new_n538), .A3(new_n575), .A4(new_n661), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n817), .B2(new_n595), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n709), .B1(new_n708), .B2(new_n621), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n703), .A2(KEYINPUT105), .A3(new_n622), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n815), .B(new_n818), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n797), .A2(new_n798), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n619), .A3(new_n702), .ZN(new_n823));
  INV_X1    g637(.A(new_n706), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n812), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n795), .B(new_n794), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(KEYINPUT53), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n814), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT54), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n795), .A2(new_n794), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n691), .A2(new_n624), .A3(new_n782), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n782), .B1(new_n691), .B2(new_n624), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n651), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n832), .B1(new_n835), .B2(new_n792), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n778), .B1(new_n826), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n795), .B(KEYINPUT52), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n813), .A2(new_n838), .A3(KEYINPUT53), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n831), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n777), .A2(new_n830), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n776), .A2(KEYINPUT115), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n535), .A2(new_n575), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n759), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n772), .A2(new_n841), .A3(new_n842), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(G952), .A2(G953), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n751), .B1(new_n847), .B2(new_n848), .ZN(G75));
  OAI21_X1  g663(.A(KEYINPUT53), .B1(new_n796), .B2(new_n813), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n826), .A2(new_n778), .A3(new_n827), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n331), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT56), .B1(new_n853), .B2(G210), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n433), .A2(new_n431), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(new_n428), .Z(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT55), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n854), .B(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n279), .A2(G952), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT117), .Z(new_n860));
  AND2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(G51));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT54), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n840), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n852), .A2(KEYINPUT118), .A3(new_n831), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n302), .B(KEYINPUT57), .Z(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n443), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n716), .B(KEYINPUT119), .Z(new_n869));
  AND2_X1   g683(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n859), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(KEYINPUT120), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n870), .B1(new_n867), .B2(new_n443), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(new_n859), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(G54));
  NAND3_X1  g692(.A1(new_n853), .A2(KEYINPUT58), .A3(G475), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(new_n373), .Z(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n859), .ZN(G60));
  NAND2_X1  g695(.A1(new_n589), .A2(new_n590), .ZN(new_n882));
  XNOR2_X1  g696(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n883));
  NAND2_X1  g697(.A1(G478), .A2(G902), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n864), .A2(new_n882), .A3(new_n865), .A4(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n887), .A2(KEYINPUT122), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(KEYINPUT122), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n885), .B1(new_n830), .B2(new_n840), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n860), .B1(new_n890), .B2(new_n882), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(G63));
  XNOR2_X1  g706(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n325), .A2(new_n331), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n850), .A2(new_n851), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n564), .ZN(new_n897));
  INV_X1    g711(.A(new_n607), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n897), .B(new_n860), .C1(new_n898), .C2(new_n896), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g714(.A(G953), .B1(new_n388), .B2(new_n399), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n803), .A2(new_n812), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n902), .A2(KEYINPUT124), .A3(new_n279), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT124), .B1(new_n902), .B2(new_n279), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n855), .B1(G898), .B2(new_n279), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(G69));
  OAI21_X1  g721(.A(new_n459), .B1(KEYINPUT30), .B2(new_n511), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT125), .Z(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n369), .ZN(new_n910));
  NAND2_X1  g724(.A1(G900), .A2(G953), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n744), .A2(new_n736), .ZN(new_n912));
  INV_X1    g726(.A(new_n712), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n843), .A2(new_n614), .A3(new_n641), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n824), .B1(new_n721), .B2(new_n914), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n912), .A2(new_n913), .A3(new_n835), .A4(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n910), .B(new_n911), .C1(new_n917), .C2(G953), .ZN(new_n918));
  NAND2_X1  g732(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n784), .A2(new_n643), .A3(new_n919), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n920), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n921));
  INV_X1    g735(.A(new_n912), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n708), .B(new_n627), .C1(new_n593), .C2(new_n807), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n920), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(new_n279), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n918), .B1(new_n926), .B2(new_n910), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n279), .B1(G227), .B2(G900), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n918), .B2(KEYINPUT127), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n927), .B(new_n929), .Z(G72));
  NAND2_X1  g744(.A1(G472), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT63), .Z(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n925), .B2(new_n902), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n474), .A3(new_n470), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n917), .B2(new_n902), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n475), .A3(new_n484), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n486), .A2(new_n634), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n829), .A2(new_n932), .A3(new_n937), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n873), .A2(new_n934), .A3(new_n936), .A4(new_n938), .ZN(G57));
endmodule


