

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U558 ( .A1(G2104), .A2(n541), .ZN(n887) );
  AND2_X2 U559 ( .A1(n541), .A2(G2104), .ZN(n884) );
  NOR2_X1 U560 ( .A1(G651), .A2(n547), .ZN(n798) );
  AND2_X1 U561 ( .A1(n691), .A2(n952), .ZN(n525) );
  NOR2_X1 U562 ( .A1(n706), .A2(KEYINPUT33), .ZN(n526) );
  XNOR2_X1 U563 ( .A(KEYINPUT32), .B(KEYINPUT99), .ZN(n678) );
  XNOR2_X1 U564 ( .A(n679), .B(n678), .ZN(n686) );
  NOR2_X1 U565 ( .A1(n686), .A2(n685), .ZN(n699) );
  INV_X1 U566 ( .A(KEYINPUT101), .ZN(n695) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n792) );
  INV_X1 U568 ( .A(G651), .ZN(n527) );
  NOR2_X1 U569 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U570 ( .A(n528), .B(KEYINPUT66), .Z(n529) );
  XNOR2_X1 U571 ( .A(KEYINPUT1), .B(n529), .ZN(n796) );
  XOR2_X1 U572 ( .A(KEYINPUT0), .B(G543), .Z(n547) );
  NAND2_X1 U573 ( .A1(G87), .A2(n547), .ZN(n531) );
  NAND2_X1 U574 ( .A1(G74), .A2(G651), .ZN(n530) );
  NAND2_X1 U575 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U576 ( .A1(n796), .A2(n532), .ZN(n534) );
  NAND2_X1 U577 ( .A1(n798), .A2(G49), .ZN(n533) );
  NAND2_X1 U578 ( .A1(n534), .A2(n533), .ZN(G288) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U580 ( .A1(G113), .A2(n889), .ZN(n535) );
  XNOR2_X1 U581 ( .A(n535), .B(KEYINPUT64), .ZN(n538) );
  INV_X1 U582 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U583 ( .A1(G101), .A2(n884), .ZN(n536) );
  XOR2_X1 U584 ( .A(KEYINPUT23), .B(n536), .Z(n537) );
  NAND2_X1 U585 ( .A1(n538), .A2(n537), .ZN(n545) );
  XNOR2_X1 U586 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n540) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  XNOR2_X2 U588 ( .A(n540), .B(n539), .ZN(n883) );
  NAND2_X1 U589 ( .A1(G137), .A2(n883), .ZN(n543) );
  NAND2_X1 U590 ( .A1(G125), .A2(n887), .ZN(n542) );
  NAND2_X1 U591 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U592 ( .A1(n545), .A2(n544), .ZN(G160) );
  NAND2_X1 U593 ( .A1(n792), .A2(G90), .ZN(n546) );
  XOR2_X1 U594 ( .A(KEYINPUT69), .B(n546), .Z(n549) );
  INV_X1 U595 ( .A(n547), .ZN(n631) );
  AND2_X1 U596 ( .A1(n631), .A2(G651), .ZN(n793) );
  NAND2_X1 U597 ( .A1(n793), .A2(G77), .ZN(n548) );
  NAND2_X1 U598 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U599 ( .A(n550), .B(KEYINPUT9), .ZN(n552) );
  NAND2_X1 U600 ( .A1(G52), .A2(n798), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U602 ( .A1(n796), .A2(G64), .ZN(n553) );
  XOR2_X1 U603 ( .A(KEYINPUT68), .B(n553), .Z(n554) );
  NOR2_X1 U604 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U605 ( .A(KEYINPUT70), .B(n556), .Z(G301) );
  INV_X1 U606 ( .A(G301), .ZN(G171) );
  NAND2_X1 U607 ( .A1(n792), .A2(G89), .ZN(n557) );
  XNOR2_X1 U608 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U609 ( .A1(G76), .A2(n793), .ZN(n558) );
  NAND2_X1 U610 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U611 ( .A(KEYINPUT5), .B(n560), .ZN(n567) );
  XNOR2_X1 U612 ( .A(KEYINPUT6), .B(KEYINPUT78), .ZN(n565) );
  NAND2_X1 U613 ( .A1(n798), .A2(G51), .ZN(n563) );
  NAND2_X1 U614 ( .A1(G63), .A2(n796), .ZN(n561) );
  XOR2_X1 U615 ( .A(KEYINPUT77), .B(n561), .Z(n562) );
  NAND2_X1 U616 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U617 ( .A(n565), .B(n564), .Z(n566) );
  NAND2_X1 U618 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U619 ( .A(KEYINPUT7), .B(n568), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G88), .A2(n792), .ZN(n570) );
  NAND2_X1 U622 ( .A1(G75), .A2(n793), .ZN(n569) );
  NAND2_X1 U623 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U624 ( .A1(n798), .A2(G50), .ZN(n572) );
  NAND2_X1 U625 ( .A1(G62), .A2(n796), .ZN(n571) );
  NAND2_X1 U626 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U627 ( .A1(n574), .A2(n573), .ZN(G166) );
  INV_X1 U628 ( .A(G166), .ZN(G303) );
  NAND2_X1 U629 ( .A1(n798), .A2(G48), .ZN(n576) );
  NAND2_X1 U630 ( .A1(G61), .A2(n796), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U632 ( .A1(n793), .A2(G73), .ZN(n577) );
  XOR2_X1 U633 ( .A(KEYINPUT2), .B(n577), .Z(n578) );
  NOR2_X1 U634 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U635 ( .A1(n792), .A2(G86), .ZN(n580) );
  NAND2_X1 U636 ( .A1(n581), .A2(n580), .ZN(G305) );
  NAND2_X1 U637 ( .A1(G85), .A2(n792), .ZN(n583) );
  NAND2_X1 U638 ( .A1(G72), .A2(n793), .ZN(n582) );
  NAND2_X1 U639 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U640 ( .A1(G60), .A2(n796), .ZN(n584) );
  XNOR2_X1 U641 ( .A(KEYINPUT67), .B(n584), .ZN(n585) );
  NOR2_X1 U642 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U643 ( .A1(n798), .A2(G47), .ZN(n587) );
  NAND2_X1 U644 ( .A1(n588), .A2(n587), .ZN(G290) );
  NOR2_X1 U645 ( .A1(G1976), .A2(G288), .ZN(n955) );
  INV_X1 U646 ( .A(G1384), .ZN(n589) );
  AND2_X1 U647 ( .A1(G40), .A2(n589), .ZN(n590) );
  NAND2_X1 U648 ( .A1(G160), .A2(n590), .ZN(n599) );
  NAND2_X1 U649 ( .A1(G126), .A2(n887), .ZN(n591) );
  XOR2_X1 U650 ( .A(KEYINPUT92), .B(n591), .Z(n593) );
  AND2_X1 U651 ( .A1(G114), .A2(n889), .ZN(n592) );
  NOR2_X1 U652 ( .A1(n593), .A2(n592), .ZN(n598) );
  NAND2_X1 U653 ( .A1(G138), .A2(n883), .ZN(n595) );
  NAND2_X1 U654 ( .A1(G102), .A2(n884), .ZN(n594) );
  NAND2_X1 U655 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U656 ( .A(n596), .B(KEYINPUT93), .ZN(n597) );
  AND2_X1 U657 ( .A1(n598), .A2(n597), .ZN(G164) );
  NOR2_X1 U658 ( .A1(n599), .A2(G164), .ZN(n643) );
  INV_X1 U659 ( .A(n643), .ZN(n659) );
  NAND2_X1 U660 ( .A1(G8), .A2(n659), .ZN(n706) );
  INV_X1 U661 ( .A(n706), .ZN(n692) );
  NAND2_X1 U662 ( .A1(n955), .A2(n692), .ZN(n600) );
  NAND2_X1 U663 ( .A1(n600), .A2(KEYINPUT33), .ZN(n694) );
  INV_X1 U664 ( .A(n659), .ZN(n645) );
  XOR2_X1 U665 ( .A(G2078), .B(KEYINPUT25), .Z(n1008) );
  NAND2_X1 U666 ( .A1(n645), .A2(n1008), .ZN(n602) );
  NAND2_X1 U667 ( .A1(G1961), .A2(n659), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U669 ( .A(KEYINPUT96), .B(n603), .Z(n665) );
  NAND2_X1 U670 ( .A1(n665), .A2(G171), .ZN(n658) );
  NAND2_X1 U671 ( .A1(G91), .A2(n792), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G78), .A2(n793), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U674 ( .A(n606), .B(KEYINPUT71), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G53), .A2(n798), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U677 ( .A1(n796), .A2(G65), .ZN(n609) );
  XOR2_X1 U678 ( .A(KEYINPUT72), .B(n609), .Z(n610) );
  NOR2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n958) );
  NAND2_X1 U680 ( .A1(n643), .A2(G2072), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n612), .B(KEYINPUT27), .ZN(n614) );
  INV_X1 U682 ( .A(G1956), .ZN(n957) );
  NOR2_X1 U683 ( .A1(n957), .A2(n645), .ZN(n613) );
  NOR2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n616) );
  NOR2_X1 U685 ( .A1(n958), .A2(n616), .ZN(n615) );
  XOR2_X1 U686 ( .A(n615), .B(KEYINPUT28), .Z(n655) );
  NAND2_X1 U687 ( .A1(n958), .A2(n616), .ZN(n653) );
  AND2_X1 U688 ( .A1(n798), .A2(G54), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G66), .A2(n796), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G92), .A2(n792), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G79), .A2(n793), .ZN(n617) );
  AND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U695 ( .A(KEYINPUT15), .B(n623), .ZN(n965) );
  NAND2_X1 U696 ( .A1(G1341), .A2(n659), .ZN(n624) );
  XNOR2_X1 U697 ( .A(KEYINPUT97), .B(n624), .ZN(n640) );
  NAND2_X1 U698 ( .A1(G1996), .A2(n643), .ZN(n625) );
  XNOR2_X1 U699 ( .A(KEYINPUT26), .B(n625), .ZN(n638) );
  NAND2_X1 U700 ( .A1(G56), .A2(n796), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(KEYINPUT14), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G43), .A2(n798), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n637) );
  NAND2_X1 U704 ( .A1(n792), .A2(G81), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n629), .B(KEYINPUT12), .ZN(n633) );
  AND2_X1 U706 ( .A1(G68), .A2(G651), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U709 ( .A(KEYINPUT13), .B(n634), .Z(n635) );
  XNOR2_X1 U710 ( .A(KEYINPUT74), .B(n635), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n902) );
  NAND2_X1 U712 ( .A1(n638), .A2(n902), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n642) );
  INV_X1 U714 ( .A(n642), .ZN(n641) );
  NAND2_X1 U715 ( .A1(n965), .A2(n641), .ZN(n651) );
  INV_X1 U716 ( .A(n965), .ZN(n789) );
  NAND2_X1 U717 ( .A1(n789), .A2(n642), .ZN(n649) );
  AND2_X1 U718 ( .A1(n643), .A2(G2067), .ZN(n644) );
  XOR2_X1 U719 ( .A(n644), .B(KEYINPUT98), .Z(n647) );
  NAND2_X1 U720 ( .A1(n659), .A2(G1348), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U724 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U726 ( .A(n656), .B(KEYINPUT29), .Z(n657) );
  NAND2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n670) );
  INV_X1 U728 ( .A(KEYINPUT30), .ZN(n663) );
  NOR2_X1 U729 ( .A1(G1966), .A2(n706), .ZN(n683) );
  NOR2_X1 U730 ( .A1(G2084), .A2(n659), .ZN(n681) );
  INV_X1 U731 ( .A(n681), .ZN(n660) );
  NAND2_X1 U732 ( .A1(G8), .A2(n660), .ZN(n661) );
  NOR2_X1 U733 ( .A1(n683), .A2(n661), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(n664) );
  NOR2_X1 U735 ( .A1(G168), .A2(n664), .ZN(n667) );
  NOR2_X1 U736 ( .A1(n665), .A2(G171), .ZN(n666) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U738 ( .A(KEYINPUT31), .B(n668), .Z(n669) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n680) );
  NAND2_X1 U740 ( .A1(n680), .A2(G286), .ZN(n677) );
  INV_X1 U741 ( .A(G8), .ZN(n675) );
  NOR2_X1 U742 ( .A1(G1971), .A2(n706), .ZN(n672) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n659), .ZN(n671) );
  NOR2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n673), .A2(G303), .ZN(n674) );
  OR2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n676) );
  AND2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U748 ( .A1(G8), .A2(n681), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n680), .A2(n682), .ZN(n684) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  INV_X1 U751 ( .A(n955), .ZN(n689) );
  NOR2_X1 U752 ( .A1(G1971), .A2(G303), .ZN(n687) );
  XOR2_X1 U753 ( .A(n687), .B(KEYINPUT100), .Z(n688) );
  NAND2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n690) );
  OR2_X1 U755 ( .A1(n699), .A2(n690), .ZN(n691) );
  NAND2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n952) );
  NAND2_X1 U757 ( .A1(n525), .A2(n526), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n696) );
  XNOR2_X1 U759 ( .A(n696), .B(n695), .ZN(n697) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n949) );
  NAND2_X1 U761 ( .A1(n697), .A2(n949), .ZN(n698) );
  XNOR2_X1 U762 ( .A(n698), .B(KEYINPUT102), .ZN(n710) );
  INV_X1 U763 ( .A(n699), .ZN(n702) );
  NOR2_X1 U764 ( .A1(G2090), .A2(G303), .ZN(n700) );
  NAND2_X1 U765 ( .A1(G8), .A2(n700), .ZN(n701) );
  NAND2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U767 ( .A1(n703), .A2(n706), .ZN(n708) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XOR2_X1 U769 ( .A(n704), .B(KEYINPUT24), .Z(n705) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n739) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n712) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n711) );
  NOR2_X1 U775 ( .A1(n712), .A2(n711), .ZN(n753) );
  NAND2_X1 U776 ( .A1(G140), .A2(n883), .ZN(n714) );
  NAND2_X1 U777 ( .A1(G104), .A2(n884), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U779 ( .A(KEYINPUT34), .B(n715), .ZN(n720) );
  NAND2_X1 U780 ( .A1(G128), .A2(n887), .ZN(n717) );
  NAND2_X1 U781 ( .A1(G116), .A2(n889), .ZN(n716) );
  NAND2_X1 U782 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U783 ( .A(n718), .B(KEYINPUT35), .Z(n719) );
  NOR2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U785 ( .A(KEYINPUT36), .B(n721), .Z(n722) );
  XOR2_X1 U786 ( .A(KEYINPUT94), .B(n722), .Z(n898) );
  XNOR2_X1 U787 ( .A(KEYINPUT37), .B(G2067), .ZN(n751) );
  NOR2_X1 U788 ( .A1(n898), .A2(n751), .ZN(n930) );
  NAND2_X1 U789 ( .A1(n753), .A2(n930), .ZN(n749) );
  NAND2_X1 U790 ( .A1(G131), .A2(n883), .ZN(n724) );
  NAND2_X1 U791 ( .A1(G95), .A2(n884), .ZN(n723) );
  NAND2_X1 U792 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U793 ( .A1(G119), .A2(n887), .ZN(n726) );
  NAND2_X1 U794 ( .A1(G107), .A2(n889), .ZN(n725) );
  NAND2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n867) );
  XNOR2_X1 U797 ( .A(KEYINPUT95), .B(G1991), .ZN(n1007) );
  NOR2_X1 U798 ( .A1(n867), .A2(n1007), .ZN(n737) );
  NAND2_X1 U799 ( .A1(G141), .A2(n883), .ZN(n730) );
  NAND2_X1 U800 ( .A1(G129), .A2(n887), .ZN(n729) );
  NAND2_X1 U801 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U802 ( .A1(n884), .A2(G105), .ZN(n731) );
  XOR2_X1 U803 ( .A(KEYINPUT38), .B(n731), .Z(n732) );
  NOR2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U805 ( .A1(n889), .A2(G117), .ZN(n734) );
  NAND2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n895) );
  AND2_X1 U807 ( .A1(G1996), .A2(n895), .ZN(n736) );
  OR2_X1 U808 ( .A1(n737), .A2(n736), .ZN(n935) );
  NAND2_X1 U809 ( .A1(n935), .A2(n753), .ZN(n742) );
  AND2_X1 U810 ( .A1(n749), .A2(n742), .ZN(n738) );
  AND2_X1 U811 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U812 ( .A(G1986), .B(G290), .ZN(n963) );
  NAND2_X1 U813 ( .A1(n963), .A2(n753), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n756) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n895), .ZN(n932) );
  INV_X1 U816 ( .A(n742), .ZN(n746) );
  NAND2_X1 U817 ( .A1(n1007), .A2(n867), .ZN(n743) );
  XNOR2_X1 U818 ( .A(n743), .B(KEYINPUT103), .ZN(n934) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n744) );
  NOR2_X1 U820 ( .A1(n934), .A2(n744), .ZN(n745) );
  NOR2_X1 U821 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U822 ( .A1(n932), .A2(n747), .ZN(n748) );
  XNOR2_X1 U823 ( .A(n748), .B(KEYINPUT39), .ZN(n750) );
  NAND2_X1 U824 ( .A1(n750), .A2(n749), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n898), .A2(n751), .ZN(n927) );
  NAND2_X1 U826 ( .A1(n752), .A2(n927), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n758) );
  XNOR2_X1 U829 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n757) );
  XNOR2_X1 U830 ( .A(n758), .B(n757), .ZN(G329) );
  AND2_X1 U831 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U832 ( .A(G132), .ZN(G219) );
  INV_X1 U833 ( .A(G82), .ZN(G220) );
  INV_X1 U834 ( .A(G57), .ZN(G237) );
  INV_X1 U835 ( .A(G120), .ZN(G236) );
  NAND2_X1 U836 ( .A1(G7), .A2(G661), .ZN(n760) );
  XOR2_X1 U837 ( .A(n760), .B(KEYINPUT10), .Z(n832) );
  NAND2_X1 U838 ( .A1(n832), .A2(G567), .ZN(n761) );
  XOR2_X1 U839 ( .A(KEYINPUT11), .B(n761), .Z(G234) );
  INV_X1 U840 ( .A(G860), .ZN(n791) );
  INV_X1 U841 ( .A(n902), .ZN(n968) );
  NOR2_X1 U842 ( .A1(n791), .A2(n968), .ZN(n762) );
  XNOR2_X1 U843 ( .A(n762), .B(KEYINPUT75), .ZN(G153) );
  INV_X1 U844 ( .A(G868), .ZN(n772) );
  NOR2_X1 U845 ( .A1(n772), .A2(G171), .ZN(n763) );
  XOR2_X1 U846 ( .A(n763), .B(KEYINPUT76), .Z(n765) );
  NAND2_X1 U847 ( .A1(n772), .A2(n965), .ZN(n764) );
  NAND2_X1 U848 ( .A1(n765), .A2(n764), .ZN(G284) );
  XNOR2_X1 U849 ( .A(n958), .B(KEYINPUT73), .ZN(G299) );
  NOR2_X1 U850 ( .A1(G286), .A2(n772), .ZN(n766) );
  XOR2_X1 U851 ( .A(KEYINPUT79), .B(n766), .Z(n768) );
  NOR2_X1 U852 ( .A1(G868), .A2(G299), .ZN(n767) );
  NOR2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U854 ( .A(KEYINPUT80), .B(n769), .ZN(G297) );
  NAND2_X1 U855 ( .A1(n791), .A2(G559), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n770), .A2(n789), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U858 ( .A1(n965), .A2(n772), .ZN(n773) );
  XNOR2_X1 U859 ( .A(n773), .B(KEYINPUT81), .ZN(n774) );
  NOR2_X1 U860 ( .A1(G559), .A2(n774), .ZN(n776) );
  NOR2_X1 U861 ( .A1(G868), .A2(n968), .ZN(n775) );
  NOR2_X1 U862 ( .A1(n776), .A2(n775), .ZN(G282) );
  XNOR2_X1 U863 ( .A(G2100), .B(KEYINPUT85), .ZN(n788) );
  NAND2_X1 U864 ( .A1(G123), .A2(n887), .ZN(n777) );
  XNOR2_X1 U865 ( .A(n777), .B(KEYINPUT82), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(KEYINPUT18), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G135), .A2(n883), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U869 ( .A(n781), .B(KEYINPUT83), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G99), .A2(n884), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n889), .A2(G111), .ZN(n784) );
  XOR2_X1 U873 ( .A(KEYINPUT84), .B(n784), .Z(n785) );
  NOR2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n941) );
  XNOR2_X1 U875 ( .A(n941), .B(G2096), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(G156) );
  NAND2_X1 U877 ( .A1(G559), .A2(n789), .ZN(n790) );
  XOR2_X1 U878 ( .A(n790), .B(n968), .Z(n810) );
  NAND2_X1 U879 ( .A1(n791), .A2(n810), .ZN(n803) );
  NAND2_X1 U880 ( .A1(G93), .A2(n792), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G80), .A2(n793), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n802) );
  NAND2_X1 U883 ( .A1(G67), .A2(n796), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(KEYINPUT86), .ZN(n800) );
  NAND2_X1 U885 ( .A1(G55), .A2(n798), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n812) );
  XOR2_X1 U888 ( .A(n803), .B(n812), .Z(G145) );
  XNOR2_X1 U889 ( .A(n812), .B(G290), .ZN(n804) );
  XNOR2_X1 U890 ( .A(n804), .B(G299), .ZN(n805) );
  XNOR2_X1 U891 ( .A(KEYINPUT19), .B(n805), .ZN(n807) );
  XNOR2_X1 U892 ( .A(G288), .B(KEYINPUT87), .ZN(n806) );
  XNOR2_X1 U893 ( .A(n807), .B(n806), .ZN(n808) );
  XOR2_X1 U894 ( .A(n808), .B(G166), .Z(n809) );
  XNOR2_X1 U895 ( .A(n809), .B(G305), .ZN(n901) );
  XNOR2_X1 U896 ( .A(n810), .B(n901), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n811), .A2(G868), .ZN(n814) );
  OR2_X1 U898 ( .A1(G868), .A2(n812), .ZN(n813) );
  NAND2_X1 U899 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U900 ( .A1(G2078), .A2(G2084), .ZN(n816) );
  XOR2_X1 U901 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n815) );
  XNOR2_X1 U902 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U907 ( .A1(G236), .A2(G237), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G69), .A2(n820), .ZN(n821) );
  XNOR2_X1 U909 ( .A(KEYINPUT89), .B(n821), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n822), .A2(G108), .ZN(n838) );
  NAND2_X1 U911 ( .A1(G567), .A2(n838), .ZN(n827) );
  NOR2_X1 U912 ( .A1(G220), .A2(G219), .ZN(n823) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U914 ( .A1(G218), .A2(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(G96), .A2(n825), .ZN(n839) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n839), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U918 ( .A(KEYINPUT90), .B(n828), .ZN(n837) );
  NAND2_X1 U919 ( .A1(G661), .A2(G483), .ZN(n829) );
  XOR2_X1 U920 ( .A(KEYINPUT91), .B(n829), .Z(n830) );
  NOR2_X1 U921 ( .A1(n837), .A2(n830), .ZN(n834) );
  NAND2_X1 U922 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(n832), .A2(G2106), .ZN(n831) );
  XNOR2_X1 U924 ( .A(n831), .B(KEYINPUT106), .ZN(G217) );
  INV_X1 U925 ( .A(n832), .ZN(G223) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U927 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U930 ( .A(KEYINPUT107), .B(n836), .Z(G188) );
  INV_X1 U931 ( .A(n837), .ZN(G319) );
  INV_X1 U933 ( .A(G108), .ZN(G238) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  NOR2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  XOR2_X1 U937 ( .A(G2100), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U938 ( .A(G2072), .B(KEYINPUT42), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U940 ( .A(n842), .B(G2678), .Z(n844) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2090), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U943 ( .A(KEYINPUT108), .B(G2096), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(G227) );
  XNOR2_X1 U947 ( .A(G1981), .B(n957), .ZN(n850) );
  XNOR2_X1 U948 ( .A(G1966), .B(G1961), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n851), .B(KEYINPUT41), .Z(n853) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U953 ( .A(G2474), .B(G1976), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1971), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G100), .A2(n884), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G112), .A2(n889), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U960 ( .A(KEYINPUT110), .B(n860), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G124), .A2(n887), .ZN(n861) );
  XOR2_X1 U962 ( .A(KEYINPUT44), .B(n861), .Z(n862) );
  XNOR2_X1 U963 ( .A(n862), .B(KEYINPUT109), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G136), .A2(n883), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U966 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n869) );
  XNOR2_X1 U968 ( .A(n867), .B(KEYINPUT112), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n878) );
  NAND2_X1 U970 ( .A1(G130), .A2(n887), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G118), .A2(n889), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G142), .A2(n883), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G106), .A2(n884), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U976 ( .A(n874), .B(KEYINPUT45), .Z(n875) );
  NOR2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(n878), .B(n877), .Z(n879) );
  XOR2_X1 U979 ( .A(n879), .B(n941), .Z(n881) );
  XNOR2_X1 U980 ( .A(G164), .B(G160), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U982 ( .A(n882), .B(G162), .Z(n897) );
  NAND2_X1 U983 ( .A1(G139), .A2(n883), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G103), .A2(n884), .ZN(n885) );
  NAND2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U986 ( .A1(n887), .A2(G127), .ZN(n888) );
  XOR2_X1 U987 ( .A(KEYINPUT111), .B(n888), .Z(n891) );
  NAND2_X1 U988 ( .A1(n889), .A2(G115), .ZN(n890) );
  NAND2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U990 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n923) );
  XOR2_X1 U992 ( .A(n895), .B(n923), .Z(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U995 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U996 ( .A(n901), .B(G286), .Z(n904) );
  XOR2_X1 U997 ( .A(n965), .B(n902), .Z(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U999 ( .A(n905), .B(G301), .Z(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U1001 ( .A(G2430), .B(G2451), .Z(n908) );
  XNOR2_X1 U1002 ( .A(G2446), .B(G2427), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n915) );
  XOR2_X1 U1004 ( .A(G2438), .B(G2435), .Z(n910) );
  XNOR2_X1 U1005 ( .A(G2443), .B(KEYINPUT105), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1007 ( .A(n911), .B(G2454), .Z(n913) );
  XNOR2_X1 U1008 ( .A(G1341), .B(G1348), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1011 ( .A1(n916), .A2(G14), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(n922), .A2(G319), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  INV_X1 U1020 ( .A(n922), .ZN(G401) );
  INV_X1 U1021 ( .A(KEYINPUT55), .ZN(n1027) );
  XOR2_X1 U1022 ( .A(G2072), .B(n923), .Z(n925) );
  XOR2_X1 U1023 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n926), .B(KEYINPUT50), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n944) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n933), .Z(n940) );
  OR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(G2084), .B(G160), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(KEYINPUT113), .B(n936), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT114), .B(n945), .ZN(n946) );
  XOR2_X1 U1039 ( .A(KEYINPUT52), .B(n946), .Z(n947) );
  NAND2_X1 U1040 ( .A1(n1027), .A2(n947), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1042 ( .A(KEYINPUT56), .B(G16), .ZN(n977) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G168), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT57), .B(n951), .ZN(n975) );
  XOR2_X1 U1046 ( .A(G303), .B(G1971), .Z(n953) );
  NAND2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1049 ( .A(KEYINPUT118), .B(n956), .Z(n960) );
  XNOR2_X1 U1050 ( .A(n958), .B(n957), .ZN(n959) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(n961), .B(KEYINPUT119), .ZN(n962) );
  NOR2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1054 ( .A(KEYINPUT120), .B(n964), .Z(n967) );
  XNOR2_X1 U1055 ( .A(n965), .B(G1348), .ZN(n966) );
  NOR2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n972) );
  XNOR2_X1 U1057 ( .A(n968), .B(G1341), .ZN(n970) );
  XOR2_X1 U1058 ( .A(G171), .B(G1961), .Z(n969) );
  NOR2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1060 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(KEYINPUT121), .B(n973), .ZN(n974) );
  NAND2_X1 U1062 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1063 ( .A1(n977), .A2(n976), .ZN(n1006) );
  XOR2_X1 U1064 ( .A(G16), .B(KEYINPUT122), .Z(n1004) );
  XOR2_X1 U1065 ( .A(G1961), .B(G5), .Z(n989) );
  XNOR2_X1 U1066 ( .A(KEYINPUT59), .B(G1348), .ZN(n978) );
  XNOR2_X1 U1067 ( .A(n978), .B(G4), .ZN(n983) );
  XNOR2_X1 U1068 ( .A(KEYINPUT123), .B(G20), .ZN(n979) );
  XOR2_X1 U1069 ( .A(n979), .B(G1956), .Z(n981) );
  XNOR2_X1 U1070 ( .A(G6), .B(G1981), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(KEYINPUT124), .B(G1341), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(G19), .B(n984), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(KEYINPUT60), .B(n987), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G21), .B(G1966), .ZN(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(KEYINPUT125), .B(n992), .ZN(n1000) );
  XOR2_X1 U1081 ( .A(G1986), .B(G24), .Z(n996) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G22), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G23), .B(G1976), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(KEYINPUT126), .B(n997), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(KEYINPUT58), .B(n998), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(n1002), .B(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1033) );
  XOR2_X1 U1093 ( .A(G2090), .B(G35), .Z(n1022) );
  XOR2_X1 U1094 ( .A(n1007), .B(G25), .Z(n1010) );
  XNOR2_X1 U1095 ( .A(G27), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1018) );
  XOR2_X1 U1097 ( .A(G32), .B(G1996), .Z(n1011) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(G28), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(G2067), .B(G26), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G2072), .B(G33), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1014), .B(KEYINPUT115), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(n1019), .B(KEYINPUT53), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(n1020), .B(KEYINPUT116), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(G34), .B(G2084), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(KEYINPUT54), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1111 ( .A(n1027), .B(n1026), .Z(n1029) );
  INV_X1 U1112 ( .A(G29), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(G11), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT117), .B(n1031), .Z(n1032) );
  NOR2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1117 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1036), .ZN(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
endmodule

