//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT75), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n203), .A3(new_n207), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(KEYINPUT75), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G183gat), .ZN(new_n221));
  INV_X1    g020(.A(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n226), .B1(KEYINPUT23), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT66), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n227), .A2(new_n234), .A3(KEYINPUT23), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n225), .B(new_n228), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n236), .A2(KEYINPUT67), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT67), .B1(new_n236), .B2(new_n237), .ZN(new_n239));
  OAI211_X1 g038(.A(KEYINPUT25), .B(new_n228), .C1(new_n233), .C2(new_n235), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n220), .A2(KEYINPUT68), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n224), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(new_n218), .B2(new_n219), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n238), .A2(new_n239), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n248), .B1(new_n227), .B2(new_n249), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n250), .A2(KEYINPUT70), .B1(new_n249), .B2(new_n227), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(KEYINPUT70), .B2(new_n250), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253));
  OR3_X1    g052(.A1(new_n253), .A2(new_n221), .A3(KEYINPUT27), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT27), .B1(new_n253), .B2(new_n221), .ZN(new_n255));
  NOR2_X1   g054(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT27), .B(G183gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n222), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n259), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n252), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G226gat), .A2(G233gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n263), .B(KEYINPUT76), .Z(new_n264));
  NOR3_X1   g063(.A1(new_n247), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(KEYINPUT29), .ZN(new_n266));
  INV_X1    g065(.A(new_n239), .ZN(new_n267));
  INV_X1    g066(.A(new_n246), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n236), .A2(KEYINPUT67), .A3(new_n237), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n266), .B1(new_n270), .B2(new_n261), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n217), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n264), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n261), .A3(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n247), .A2(new_n262), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n216), .B(new_n274), .C1(new_n275), .C2(new_n266), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT77), .ZN(new_n279));
  XNOR2_X1  g078(.A(G8gat), .B(G36gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(KEYINPUT30), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT78), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n277), .A2(KEYINPUT78), .A3(KEYINPUT30), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT79), .B1(new_n277), .B2(new_n282), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT79), .ZN(new_n290));
  AOI211_X1 g089(.A(new_n290), .B(new_n281), .C1(new_n272), .C2(new_n276), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n277), .A2(new_n282), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n287), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT74), .B(G71gat), .ZN(new_n296));
  INV_X1    g095(.A(G99gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G15gat), .B(G43gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G127gat), .ZN(new_n301));
  INV_X1    g100(.A(G134gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G127gat), .A2(G134gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G113gat), .B(G120gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n303), .B(new_n304), .C1(new_n305), .C2(KEYINPUT1), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n303), .A2(new_n304), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n307), .B(new_n308), .C1(new_n305), .C2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(G120gat), .ZN(new_n312));
  INV_X1    g111(.A(G120gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G113gat), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT71), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n306), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT73), .ZN(new_n317));
  OR2_X1    g116(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n318));
  NAND2_X1  g117(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n318), .A2(new_n319), .B1(new_n303), .B2(new_n304), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n309), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT71), .B1(new_n312), .B2(new_n314), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n306), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(new_n247), .B2(new_n262), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n323), .A2(new_n324), .A3(new_n306), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n324), .B1(new_n323), .B2(new_n306), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n270), .A2(new_n330), .A3(new_n261), .ZN(new_n331));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT64), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT65), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n327), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n300), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(KEYINPUT32), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n336), .B(KEYINPUT32), .C1(new_n337), .C2(new_n300), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n331), .ZN(new_n343));
  INV_X1    g142(.A(new_n333), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n335), .A2(KEYINPUT34), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n345), .A2(KEYINPUT34), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(G141gat), .B(G148gat), .Z(new_n350));
  INV_X1    g149(.A(G155gat), .ZN(new_n351));
  INV_X1    g150(.A(G162gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(KEYINPUT2), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n350), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G141gat), .B(G148gat), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n354), .B(new_n353), .C1(new_n358), .C2(KEYINPUT2), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n216), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n357), .A2(new_n359), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n211), .B2(new_n213), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G228gat), .ZN(new_n369));
  INV_X1    g168(.A(G233gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G22gat), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n357), .A2(new_n359), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n214), .A2(new_n362), .A3(new_n215), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n360), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n364), .A2(new_n371), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n373), .B(new_n374), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT83), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT31), .B(G50gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT82), .ZN(new_n382));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n378), .A2(new_n377), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n371), .B1(new_n364), .B2(new_n367), .ZN(new_n386));
  OAI21_X1  g185(.A(G22gat), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n380), .A2(new_n384), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n389));
  AND4_X1   g188(.A1(new_n389), .A2(new_n387), .A3(new_n379), .A4(new_n384), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n340), .A2(new_n347), .A3(new_n341), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n349), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394));
  INV_X1    g193(.A(G85gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT0), .B(G57gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n316), .A2(new_n365), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n323), .A2(new_n306), .B1(new_n359), .B2(new_n357), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT5), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n365), .B1(new_n317), .B2(new_n325), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n406), .B2(KEYINPUT4), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n316), .A2(new_n361), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n360), .B1(new_n357), .B2(new_n359), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT4), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n375), .A2(new_n306), .A3(new_n323), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n405), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT4), .B1(new_n326), .B2(new_n375), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n316), .A3(new_n361), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n375), .A2(KEYINPUT4), .A3(new_n306), .A4(new_n323), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n401), .A2(KEYINPUT5), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n414), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT6), .B(new_n399), .C1(new_n413), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT81), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n316), .A2(new_n365), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n411), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n424), .B1(new_n426), .B2(new_n401), .ZN(new_n427));
  OAI211_X1 g226(.A(KEYINPUT4), .B(new_n375), .C1(new_n328), .C2(new_n329), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n400), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n402), .B1(new_n416), .B2(KEYINPUT4), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n416), .A2(new_n417), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(new_n419), .C1(KEYINPUT4), .C2(new_n406), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n398), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT81), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT6), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n423), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n431), .A2(new_n433), .A3(new_n398), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT80), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n440), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n434), .B1(new_n442), .B2(KEYINPUT80), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n437), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n295), .A2(new_n393), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT35), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n202), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n441), .ZN(new_n448));
  INV_X1    g247(.A(new_n437), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n450), .A2(new_n287), .A3(new_n292), .A4(new_n294), .ZN(new_n451));
  OAI211_X1 g250(.A(KEYINPUT86), .B(KEYINPUT35), .C1(new_n451), .C2(new_n393), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n442), .A2(new_n434), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n446), .B1(new_n437), .B2(new_n453), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n295), .A2(new_n393), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n447), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n437), .A2(new_n453), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n281), .B1(new_n272), .B2(new_n276), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT79), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n272), .A2(KEYINPUT37), .A3(new_n276), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT37), .B1(new_n272), .B2(new_n276), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n461), .A2(new_n462), .A3(new_n282), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n463), .A2(KEYINPUT38), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(KEYINPUT38), .B2(new_n465), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n458), .B(new_n460), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n414), .A2(new_n418), .ZN(new_n469));
  OR3_X1    g268(.A1(new_n469), .A2(KEYINPUT39), .A3(new_n400), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n400), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT39), .B1(new_n426), .B2(new_n401), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n470), .B(new_n398), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT40), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n434), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n295), .B(new_n475), .C1(new_n474), .C2(new_n473), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n468), .A2(new_n476), .A3(new_n391), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n391), .B(KEYINPUT84), .Z(new_n478));
  INV_X1    g277(.A(KEYINPUT36), .ZN(new_n479));
  INV_X1    g278(.A(new_n349), .ZN(new_n480));
  INV_X1    g279(.A(new_n392), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n349), .A2(KEYINPUT36), .A3(new_n392), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n478), .A2(new_n451), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n457), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT98), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n488));
  INV_X1    g287(.A(G92gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n395), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n491));
  NAND2_X1  g290(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n491), .A2(G85gat), .A3(G92gat), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494));
  AOI22_X1  g293(.A1(KEYINPUT8), .A2(new_n494), .B1(new_n395), .B2(new_n489), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G99gat), .B(G106gat), .Z(new_n497));
  OAI21_X1  g296(.A(new_n487), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n493), .A2(new_n495), .ZN(new_n499));
  INV_X1    g298(.A(new_n497), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n499), .A2(KEYINPUT98), .A3(new_n500), .A4(new_n490), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n498), .A2(new_n501), .B1(new_n497), .B2(new_n496), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(G29gat), .A2(G36gat), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(KEYINPUT14), .Z(new_n505));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(G29gat), .B2(G36gat), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n505), .A2(new_n507), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n504), .B(KEYINPUT14), .ZN(new_n512));
  INV_X1    g311(.A(new_n510), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT15), .B(new_n506), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n511), .A2(new_n514), .A3(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(G232gat), .A2(G233gat), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n502), .A2(new_n515), .B1(KEYINPUT41), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G190gat), .B(G218gat), .Z(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT99), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n523), .ZN(new_n526));
  XNOR2_X1  g325(.A(G134gat), .B(G162gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT96), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n520), .A2(KEYINPUT41), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n528), .B(new_n529), .Z(new_n530));
  AND4_X1   g329(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n530), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n525), .A2(new_n530), .B1(new_n524), .B2(new_n526), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(G57gat), .B2(G64gat), .ZN(new_n536));
  INV_X1    g335(.A(G71gat), .ZN(new_n537));
  INV_X1    g336(.A(G78gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT9), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G57gat), .ZN(new_n545));
  INV_X1    g344(.A(G64gat), .ZN(new_n546));
  OR3_X1    g345(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT92), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n545), .B2(KEYINPUT92), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT93), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n544), .A2(new_n547), .A3(new_n551), .A4(new_n548), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n542), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G127gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G155gat), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n558));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n557), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(G1gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT16), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n564), .B2(G1gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT88), .ZN(new_n568));
  INV_X1    g367(.A(G8gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n569), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n563), .A2(new_n565), .A3(new_n571), .A4(new_n566), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n553), .A2(KEYINPUT21), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT95), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n561), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G120gat), .B(G148gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G230gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(new_n370), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n498), .A2(new_n501), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT100), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n496), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n499), .A2(KEYINPUT100), .A3(new_n490), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(new_n588), .A3(new_n497), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n553), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n502), .A2(new_n553), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n584), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT101), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n595), .B(new_n584), .C1(new_n591), .C2(new_n592), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n590), .B(new_n598), .C1(new_n502), .C2(new_n553), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n502), .A2(KEYINPUT10), .A3(new_n553), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n584), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n582), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n601), .ZN(new_n603));
  INV_X1    g402(.A(new_n582), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n596), .A4(new_n594), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n534), .A2(new_n579), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n570), .A2(new_n572), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n517), .A2(new_n609), .A3(new_n518), .ZN(new_n610));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n515), .A2(new_n570), .A3(new_n572), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT18), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT89), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n610), .A2(KEYINPUT18), .A3(new_n611), .A4(new_n612), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n618), .A2(KEYINPUT90), .ZN(new_n619));
  INV_X1    g418(.A(new_n515), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n612), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n611), .B(KEYINPUT13), .Z(new_n623));
  AOI22_X1  g422(.A1(new_n618), .A2(KEYINPUT90), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n613), .A2(KEYINPUT89), .A3(new_n614), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n617), .A2(new_n619), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G197gat), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT11), .B(G169gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT91), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n631), .B1(new_n615), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n613), .A2(KEYINPUT91), .A3(new_n614), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n634), .A2(new_n619), .A3(new_n624), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n608), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n486), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n444), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G1gat), .ZN(G1324gat));
  INV_X1    g444(.A(new_n295), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n647), .B2(new_n569), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  MUX2_X1   g449(.A(KEYINPUT42), .B(new_n648), .S(new_n650), .Z(G1325gat));
  NAND2_X1  g450(.A1(new_n482), .A2(new_n483), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n641), .A2(G15gat), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n480), .A2(new_n481), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n654), .B1(G15gat), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT103), .ZN(G1326gat));
  INV_X1    g458(.A(new_n478), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n640), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT43), .B(G22gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  AOI21_X1  g462(.A(new_n534), .B1(new_n457), .B2(new_n485), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n579), .A2(new_n638), .A3(new_n606), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n643), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n666), .A2(G29gat), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT45), .Z(new_n669));
  INV_X1    g468(.A(new_n665), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT35), .B1(new_n451), .B2(new_n393), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n455), .B1(new_n671), .B2(new_n202), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n672), .A2(new_n452), .B1(new_n477), .B2(new_n484), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT44), .B1(new_n673), .B2(new_n534), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n664), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n670), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(KEYINPUT104), .A3(new_n643), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(G29gat), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT104), .B1(new_n677), .B2(new_n643), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n669), .B1(new_n679), .B2(new_n680), .ZN(G1328gat));
  NOR3_X1   g480(.A1(new_n666), .A2(G36gat), .A3(new_n646), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT46), .ZN(new_n683));
  INV_X1    g482(.A(new_n677), .ZN(new_n684));
  OAI21_X1  g483(.A(G36gat), .B1(new_n684), .B2(new_n646), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(G1329gat));
  INV_X1    g485(.A(new_n666), .ZN(new_n687));
  INV_X1    g486(.A(G43gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n655), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n684), .A2(new_n652), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT47), .B(new_n689), .C1(new_n690), .C2(new_n688), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1330gat));
  OAI21_X1  g494(.A(G50gat), .B1(new_n684), .B2(new_n660), .ZN(new_n696));
  INV_X1    g495(.A(G50gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n687), .A2(new_n697), .A3(new_n478), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n391), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n697), .B1(new_n677), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(KEYINPUT48), .ZN(new_n702));
  OAI22_X1  g501(.A1(new_n699), .A2(KEYINPUT48), .B1(new_n701), .B2(new_n702), .ZN(G1331gat));
  INV_X1    g502(.A(new_n579), .ZN(new_n704));
  NOR4_X1   g503(.A1(new_n704), .A2(new_n637), .A3(new_n533), .A4(new_n607), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n486), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n667), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT105), .B(G57gat), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1332gat));
  INV_X1    g508(.A(new_n706), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n646), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT106), .Z(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1333gat));
  OAI21_X1  g514(.A(new_n537), .B1(new_n706), .B2(new_n656), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n653), .A2(G71gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n706), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g518(.A1(new_n706), .A2(new_n660), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n538), .ZN(G1335gat));
  NOR2_X1   g520(.A1(new_n579), .A2(new_n637), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n606), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n674), .B2(new_n676), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725), .B2(new_n667), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n486), .A2(new_n533), .A3(new_n722), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n664), .A2(KEYINPUT51), .A3(new_n722), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n607), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n395), .A3(new_n643), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n726), .A2(new_n732), .ZN(G1336gat));
  NOR2_X1   g532(.A1(new_n646), .A2(G92gat), .ZN(new_n734));
  AND4_X1   g533(.A1(KEYINPUT51), .A2(new_n486), .A3(new_n533), .A4(new_n722), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT51), .B1(new_n664), .B2(new_n722), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n606), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n489), .B1(new_n724), .B2(new_n295), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n295), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n740), .A2(KEYINPUT107), .A3(G92gat), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT52), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(G92gat), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n743), .A2(KEYINPUT108), .A3(new_n744), .A4(new_n737), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n737), .A2(new_n744), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(new_n738), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n742), .A2(new_n749), .ZN(G1337gat));
  OAI21_X1  g549(.A(G99gat), .B1(new_n725), .B2(new_n652), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n731), .A2(new_n297), .A3(new_n655), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1338gat));
  INV_X1    g552(.A(G106gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n724), .B2(new_n478), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n607), .A2(G106gat), .A3(new_n391), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT109), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n729), .B2(new_n730), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT53), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n723), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n664), .A2(new_n675), .ZN(new_n761));
  AOI211_X1 g560(.A(KEYINPUT44), .B(new_n534), .C1(new_n457), .C2(new_n485), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n700), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT53), .B1(new_n763), .B2(G106gat), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n729), .A2(new_n730), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n756), .ZN(new_n767));
  INV_X1    g566(.A(new_n756), .ZN(new_n768));
  AOI211_X1 g567(.A(KEYINPUT110), .B(new_n768), .C1(new_n729), .C2(new_n730), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n764), .B(KEYINPUT111), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n756), .B1(new_n735), .B2(new_n736), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT110), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n766), .A2(new_n765), .A3(new_n756), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT111), .B1(new_n775), .B2(new_n764), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n759), .B1(new_n771), .B2(new_n776), .ZN(G1339gat));
  OR2_X1    g576(.A1(new_n608), .A2(new_n637), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n599), .A2(new_n584), .A3(new_n600), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n603), .A2(KEYINPUT54), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n604), .B1(new_n601), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n780), .A2(KEYINPUT55), .A3(new_n782), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n605), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n610), .A2(new_n612), .ZN(new_n788));
  INV_X1    g587(.A(new_n611), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(KEYINPUT112), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n622), .B2(new_n623), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT112), .B1(new_n788), .B2(new_n789), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n630), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT113), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n795), .B(new_n630), .C1(new_n791), .C2(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n636), .ZN(new_n798));
  NOR4_X1   g597(.A1(new_n787), .A2(new_n798), .A3(new_n531), .A4(new_n532), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n606), .A3(new_n636), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n787), .B2(new_n638), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n533), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n800), .B(KEYINPUT114), .C1(new_n787), .C2(new_n638), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n799), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n778), .B1(new_n805), .B2(new_n579), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(new_n643), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n646), .A3(new_n655), .A4(new_n660), .ZN(new_n808));
  OAI21_X1  g607(.A(G113gat), .B1(new_n808), .B2(new_n638), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n807), .A2(new_n646), .A3(new_n391), .A4(new_n655), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n637), .A2(new_n311), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(G1340gat));
  OAI21_X1  g611(.A(G120gat), .B1(new_n808), .B2(new_n607), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n606), .A2(new_n313), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n810), .B2(new_n814), .ZN(G1341gat));
  NOR3_X1   g614(.A1(new_n808), .A2(new_n301), .A3(new_n704), .ZN(new_n816));
  INV_X1    g615(.A(new_n810), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n579), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(KEYINPUT115), .ZN(new_n819));
  AOI21_X1  g618(.A(G127gat), .B1(new_n818), .B2(KEYINPUT115), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(G1342gat));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n302), .A3(new_n533), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n823));
  OAI21_X1  g622(.A(G134gat), .B1(new_n808), .B2(new_n534), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(KEYINPUT56), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(G1343gat));
  NOR3_X1   g625(.A1(new_n667), .A2(new_n653), .A3(new_n295), .ZN(new_n827));
  XOR2_X1   g626(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n806), .B2(new_n700), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n786), .A2(new_n605), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT55), .B1(new_n780), .B2(new_n782), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT117), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n785), .A2(new_n834), .A3(new_n605), .A4(new_n786), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n637), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n533), .B1(new_n836), .B2(new_n800), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n704), .B1(new_n837), .B2(new_n799), .ZN(new_n838));
  AOI211_X1 g637(.A(new_n830), .B(new_n660), .C1(new_n838), .C2(new_n778), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n637), .B(new_n827), .C1(new_n829), .C2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT58), .B1(new_n840), .B2(G141gat), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n653), .A2(new_n391), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n806), .A2(new_n643), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT119), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n638), .A2(G141gat), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n806), .A2(new_n846), .A3(new_n643), .A4(new_n842), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n844), .A2(new_n646), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n841), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n840), .A2(G141gat), .ZN(new_n854));
  INV_X1    g653(.A(new_n845), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n843), .A2(new_n295), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n853), .B1(new_n858), .B2(KEYINPUT58), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n840), .B2(G141gat), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n860), .A2(KEYINPUT118), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n852), .B1(new_n859), .B2(new_n862), .ZN(G1344gat));
  AND3_X1   g662(.A1(new_n844), .A2(new_n646), .A3(new_n847), .ZN(new_n864));
  INV_X1    g663(.A(G148gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n865), .A3(new_n606), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n606), .B(new_n827), .C1(new_n829), .C2(new_n839), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n865), .A2(KEYINPUT59), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n867), .A2(KEYINPUT121), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT121), .B1(new_n867), .B2(new_n868), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n838), .A2(new_n778), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n478), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(KEYINPUT122), .A3(new_n830), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n806), .A2(new_n700), .A3(new_n828), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT122), .B1(new_n874), .B2(new_n830), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n606), .B(new_n827), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n872), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n866), .B1(new_n871), .B2(new_n880), .ZN(G1345gat));
  AOI21_X1  g680(.A(G155gat), .B1(new_n864), .B2(new_n579), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n829), .A2(new_n839), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(new_n827), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n704), .A2(new_n351), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1346gat));
  AOI21_X1  g685(.A(G162gat), .B1(new_n864), .B2(new_n533), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n534), .A2(new_n352), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n884), .B2(new_n888), .ZN(G1347gat));
  NAND3_X1  g688(.A1(new_n806), .A2(KEYINPUT123), .A3(new_n667), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT123), .B1(new_n806), .B2(new_n667), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n646), .A2(new_n393), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n229), .A3(new_n637), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n667), .A2(new_n295), .A3(new_n655), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n897), .A2(KEYINPUT124), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(KEYINPUT124), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n898), .A2(new_n899), .A3(new_n478), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n806), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n638), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n896), .A2(new_n902), .ZN(G1348gat));
  NOR3_X1   g702(.A1(new_n901), .A2(new_n230), .A3(new_n607), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n895), .A2(new_n606), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n230), .ZN(G1349gat));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(KEYINPUT60), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n579), .A2(new_n258), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n894), .B(new_n909), .C1(new_n891), .C2(new_n892), .ZN(new_n910));
  OAI21_X1  g709(.A(G183gat), .B1(new_n901), .B2(new_n704), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n907), .A2(KEYINPUT60), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n912), .B(new_n913), .ZN(G1350gat));
  NAND3_X1  g713(.A1(new_n895), .A2(new_n222), .A3(new_n533), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n533), .A3(new_n806), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n916), .A2(G190gat), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT126), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n916), .A2(KEYINPUT126), .A3(new_n918), .A4(G190gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n915), .B1(new_n919), .B2(new_n921), .ZN(G1351gat));
  OR2_X1    g721(.A1(new_n877), .A2(new_n878), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n653), .A2(new_n643), .A3(new_n646), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n637), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(G197gat), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n842), .A2(new_n295), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT127), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n893), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(G197gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n930), .A3(new_n637), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n926), .A2(new_n931), .ZN(G1352gat));
  NOR2_X1   g731(.A1(new_n607), .A2(G204gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n893), .A2(new_n928), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n606), .B(new_n924), .C1(new_n877), .C2(new_n878), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G204gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n929), .A2(new_n205), .A3(new_n579), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n579), .B(new_n924), .C1(new_n877), .C2(new_n878), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(G1354gat));
  AND2_X1   g743(.A1(new_n923), .A2(new_n924), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n534), .A2(new_n206), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n893), .A2(new_n533), .A3(new_n928), .ZN(new_n947));
  AOI22_X1  g746(.A1(new_n945), .A2(new_n946), .B1(new_n206), .B2(new_n947), .ZN(G1355gat));
endmodule


