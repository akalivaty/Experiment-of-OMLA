//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n596,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1243, new_n1244;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT68), .B1(new_n467), .B2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AOI211_X1 g045(.A(new_n469), .B(new_n470), .C1(new_n465), .C2(new_n466), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n475));
  OAI211_X1 g050(.A(G101), .B(new_n470), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n474), .A2(new_n475), .A3(new_n461), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n479), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n461), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n478), .A2(new_n482), .A3(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n477), .B1(new_n483), .B2(G137), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n472), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n488));
  OR2_X1    g063(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(KEYINPUT3), .A3(new_n473), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n490), .A2(new_n470), .A3(new_n480), .A4(new_n481), .ZN(new_n491));
  INV_X1    g066(.A(G136), .ZN(new_n492));
  INV_X1    g067(.A(G124), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n490), .A2(G2105), .A3(new_n480), .A4(new_n481), .ZN(new_n494));
  OAI221_X1 g069(.A(new_n488), .B1(new_n491), .B2(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  NOR2_X1   g071(.A1(new_n470), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n500), .A2(new_n502), .A3(new_n503), .A4(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G126), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n494), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n462), .A2(new_n464), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(new_n470), .A3(G138), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n470), .A2(G138), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n490), .A2(new_n480), .A3(new_n481), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n513), .B2(KEYINPUT4), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n507), .A2(new_n514), .ZN(G164));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n523), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT7), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n533), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(KEYINPUT6), .A2(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(KEYINPUT6), .A2(G651), .ZN(new_n537));
  OAI211_X1 g112(.A(G51), .B(G543), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(G89), .B1(new_n536), .B2(new_n537), .ZN(new_n541));
  NAND2_X1  g116(.A1(G63), .A2(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(new_n520), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  INV_X1    g121(.A(KEYINPUT6), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(new_n522), .ZN(new_n548));
  NAND2_X1  g123(.A1(KEYINPUT6), .A2(G651), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n518), .A2(new_n519), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n517), .B1(new_n548), .B2(new_n549), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n550), .A2(G90), .B1(new_n551), .B2(G52), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n518), .B2(new_n519), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n552), .A2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n525), .A2(new_n560), .B1(new_n527), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n520), .A2(G56), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n522), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g143(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n569));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  OAI211_X1 g147(.A(G53), .B(G543), .C1(new_n536), .C2(new_n537), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n551), .A2(G53), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n575), .A2(new_n577), .B1(G91), .B2(new_n550), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  INV_X1    g154(.A(new_n519), .ZN(new_n580));
  NOR2_X1   g155(.A1(KEYINPUT5), .A2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(G65), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G78), .A2(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT74), .B1(new_n584), .B2(G651), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  AOI211_X1 g161(.A(new_n586), .B(new_n522), .C1(new_n582), .C2(new_n583), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n578), .B(new_n579), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n586), .B1(new_n590), .B2(new_n522), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n584), .A2(KEYINPUT74), .A3(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n579), .B1(new_n593), .B2(new_n578), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n589), .A2(new_n594), .ZN(G299));
  INV_X1    g170(.A(KEYINPUT76), .ZN(new_n596));
  XNOR2_X1  g171(.A(G166), .B(new_n596), .ZN(G303));
  NAND2_X1  g172(.A1(new_n550), .A2(G87), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n551), .A2(G49), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(G288));
  AND2_X1   g176(.A1(new_n520), .A2(G61), .ZN(new_n602));
  NAND2_X1  g177(.A1(G73), .A2(G543), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT77), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n550), .A2(G86), .B1(new_n551), .B2(G48), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G305));
  AOI22_X1  g182(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n522), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  INV_X1    g185(.A(G47), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n525), .A2(new_n610), .B1(new_n527), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n550), .A2(G92), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT10), .Z(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n580), .A2(new_n581), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n621), .A2(G651), .B1(G54), .B2(new_n551), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n615), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n615), .B1(new_n624), .B2(G868), .ZN(G321));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NOR2_X1   g202(.A1(G286), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G299), .B(KEYINPUT78), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n627), .ZN(G297));
  AOI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(new_n627), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n624), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n624), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g212(.A1(new_n478), .A2(new_n482), .A3(new_n470), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G123), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT79), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(G111), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G2105), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n483), .A2(G135), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT80), .B(G2096), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(G2105), .B1(new_n489), .B2(new_n473), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n648), .A2(new_n462), .A3(new_n464), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT13), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n647), .A2(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(KEYINPUT81), .B(KEYINPUT14), .Z(new_n654));
  XOR2_X1   g229(.A(KEYINPUT15), .B(G2435), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2438), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  AOI21_X1  g232(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n656), .B2(new_n657), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G401));
  XNOR2_X1  g244(.A(G2084), .B(G2090), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(KEYINPUT17), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n673), .B1(new_n674), .B2(new_n671), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT82), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n677), .A2(new_n670), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n671), .A2(new_n670), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n679), .C1(new_n674), .C2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G2100), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT83), .B(G2096), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n687));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1956), .B(G2474), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1961), .B(G1966), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n691), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n691), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n695), .A2(KEYINPUT20), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(KEYINPUT20), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n692), .B1(new_n689), .B2(new_n693), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT85), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(G229));
  NAND2_X1  g280(.A1(new_n566), .A2(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G16), .B2(G19), .ZN(new_n707));
  INV_X1    g282(.A(G1341), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT30), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G28), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n710), .B2(G28), .ZN(new_n713));
  AND2_X1   g288(.A1(KEYINPUT31), .A2(G11), .ZN(new_n714));
  NOR2_X1   g289(.A1(KEYINPUT31), .A2(G11), .ZN(new_n715));
  OAI22_X1  g290(.A1(new_n711), .A2(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n707), .B2(new_n708), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G5), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G171), .B2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(G21), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G168), .B2(new_n718), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n720), .A2(G1961), .B1(new_n722), .B2(G1966), .ZN(new_n723));
  NAND2_X1  g298(.A1(G115), .A2(G2104), .ZN(new_n724));
  INV_X1    g299(.A(G127), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n508), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G2105), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  INV_X1    g304(.A(G139), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n727), .B(new_n729), .C1(new_n730), .C2(new_n491), .ZN(new_n731));
  MUX2_X1   g306(.A(G33), .B(new_n731), .S(G29), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G2072), .ZN(new_n733));
  AND4_X1   g308(.A1(new_n709), .A2(new_n717), .A3(new_n723), .A4(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n718), .A2(G4), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n623), .B2(G16), .ZN(new_n736));
  INV_X1    g311(.A(G1348), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n732), .A2(G2072), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n712), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n712), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT29), .B(G2090), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n742), .B(new_n743), .Z(new_n744));
  AOI22_X1  g319(.A1(new_n737), .A2(new_n736), .B1(new_n645), .B2(G29), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n734), .A2(new_n740), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n712), .A2(G26), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  INV_X1    g323(.A(G140), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n491), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G116), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G2105), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n638), .B2(G128), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n748), .B1(new_n757), .B2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n712), .B1(KEYINPUT24), .B2(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(KEYINPUT24), .B2(G34), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n485), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2078), .ZN(new_n766));
  NAND2_X1  g341(.A1(G164), .A2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G27), .B2(G29), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n765), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n722), .A2(G1966), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT93), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n769), .B(new_n771), .C1(new_n766), .C2(new_n768), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n746), .A2(new_n760), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n718), .A2(G20), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT23), .ZN(new_n775));
  INV_X1    g350(.A(G299), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n718), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  OR2_X1    g353(.A1(G29), .A2(G32), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n648), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n638), .A2(G129), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT90), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT26), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n780), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g364(.A(KEYINPUT92), .B(new_n779), .C1(new_n789), .C2(new_n712), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n787), .A2(new_n788), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n791), .A2(new_n792), .A3(G29), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT27), .B(G1996), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n778), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n763), .A2(new_n764), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G1961), .B2(new_n720), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(KEYINPUT94), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n796), .B1(new_n790), .B2(new_n793), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n804), .A2(new_n805), .A3(new_n801), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n773), .B(new_n797), .C1(new_n803), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n718), .A2(G23), .ZN(new_n808));
  INV_X1    g383(.A(G288), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n718), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT33), .B(G1976), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT86), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n523), .A2(new_n529), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G16), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n718), .A2(G22), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n816), .ZN(new_n818));
  AOI211_X1 g393(.A(KEYINPUT86), .B(new_n818), .C1(new_n814), .C2(G16), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n812), .B1(new_n820), .B2(G1971), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT34), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n605), .A2(G16), .A3(new_n606), .ZN(new_n823));
  OR2_X1    g398(.A1(G6), .A2(G16), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT32), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n823), .A2(new_n827), .A3(new_n824), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G1981), .ZN(new_n830));
  INV_X1    g405(.A(G1981), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n826), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G1971), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n817), .B2(new_n819), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n821), .A2(new_n822), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n483), .A2(G131), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n638), .A2(G119), .ZN(new_n838));
  OR2_X1    g413(.A1(G95), .A2(G2105), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n839), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G29), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G25), .B2(G29), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G1991), .Z(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n718), .A2(G24), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n613), .B2(new_n718), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G1986), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n846), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n836), .A2(KEYINPUT87), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT87), .B1(new_n836), .B2(new_n851), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT88), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n810), .B(new_n811), .Z(new_n855));
  NAND3_X1  g430(.A1(new_n815), .A2(new_n813), .A3(new_n816), .ZN(new_n856));
  NOR2_X1   g431(.A1(G166), .A2(new_n718), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT86), .B1(new_n857), .B2(new_n818), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n858), .A3(G1971), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n835), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n830), .A2(new_n832), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n854), .B(KEYINPUT34), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n821), .A2(new_n833), .A3(new_n835), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n854), .B1(new_n864), .B2(KEYINPUT34), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n852), .A2(new_n853), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT36), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n868));
  OAI221_X1 g443(.A(new_n868), .B1(new_n865), .B2(new_n863), .C1(new_n852), .C2(new_n853), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n807), .B1(new_n867), .B2(new_n869), .ZN(G311));
  NOR2_X1   g445(.A1(G311), .A2(KEYINPUT95), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n872));
  AOI211_X1 g447(.A(new_n872), .B(new_n807), .C1(new_n869), .C2(new_n867), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(G150));
  NAND2_X1  g449(.A1(new_n624), .A2(G559), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT97), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT38), .ZN(new_n877));
  INV_X1    g452(.A(G67), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n518), .B2(new_n519), .ZN(new_n879));
  NAND2_X1  g454(.A1(G80), .A2(G543), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(KEYINPUT96), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n883), .B(new_n880), .C1(new_n619), .C2(new_n878), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n884), .A3(G651), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n550), .A2(G93), .B1(new_n551), .B2(G55), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n563), .A2(new_n564), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(G651), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n550), .A2(G81), .B1(new_n551), .B2(G43), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n885), .A2(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n877), .B(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(KEYINPUT39), .ZN(new_n896));
  INV_X1    g471(.A(G860), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(KEYINPUT39), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n887), .A2(G860), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(KEYINPUT37), .Z(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(G145));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n903));
  OR2_X1    g478(.A1(G106), .A2(G2105), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n904), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n905));
  INV_X1    g480(.A(G130), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n494), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(G142), .B2(new_n483), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n650), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n909), .A2(new_n841), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n841), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(KEYINPUT101), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(KEYINPUT101), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n499), .A2(new_n504), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(new_n638), .B2(G126), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n513), .A2(KEYINPUT4), .ZN(new_n918));
  INV_X1    g493(.A(new_n511), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT98), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT98), .B1(new_n507), .B2(new_n514), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n752), .A2(new_n756), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n731), .A2(KEYINPUT99), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n731), .A2(KEYINPUT100), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n926), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n757), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n791), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n791), .A3(new_n930), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n924), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n933), .ZN(new_n935));
  INV_X1    g510(.A(new_n924), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n935), .A2(new_n931), .A3(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n914), .B(new_n915), .C1(new_n934), .C2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n485), .B(new_n495), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n645), .B(new_n939), .Z(new_n940));
  OAI21_X1  g515(.A(new_n936), .B1(new_n935), .B2(new_n931), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n932), .A2(new_n924), .A3(new_n933), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n913), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G37), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n940), .B1(new_n938), .B2(new_n943), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n903), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n949), .A2(KEYINPUT40), .A3(new_n945), .A4(new_n944), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(G395));
  NAND2_X1  g526(.A1(new_n887), .A2(new_n627), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n634), .B(new_n894), .Z(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT102), .B1(new_n589), .B2(new_n594), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n578), .B1(new_n585), .B2(new_n587), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT75), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n588), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(new_n624), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(G299), .A2(new_n959), .A3(new_n623), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n953), .B1(new_n955), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT41), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(KEYINPUT41), .A3(new_n962), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n955), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n961), .A2(new_n962), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n954), .A2(KEYINPUT103), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n964), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n613), .B(G305), .ZN(new_n972));
  XNOR2_X1  g547(.A(G166), .B(G288), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n972), .B(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT42), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n971), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n952), .B1(new_n976), .B2(new_n627), .ZN(G295));
  OAI21_X1  g552(.A(new_n952), .B1(new_n976), .B2(new_n627), .ZN(G331));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n974), .B(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n524), .A2(G52), .A3(G543), .ZN(new_n984));
  INV_X1    g559(.A(G90), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n525), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n520), .A2(G64), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n522), .B1(new_n987), .B2(new_n555), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n619), .B1(new_n542), .B2(new_n541), .ZN(new_n989));
  OAI22_X1  g564(.A1(new_n986), .A2(new_n988), .B1(new_n989), .B2(new_n539), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n552), .A2(new_n540), .A3(new_n544), .A4(new_n557), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n892), .A2(new_n992), .A3(new_n893), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n887), .A2(new_n891), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n566), .A2(new_n885), .A3(new_n886), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n994), .A2(new_n995), .B1(new_n990), .B2(new_n991), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n983), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n994), .A2(new_n995), .A3(new_n990), .A4(new_n991), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT104), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n997), .A2(new_n961), .A3(new_n962), .A4(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT106), .ZN(new_n1001));
  INV_X1    g576(.A(new_n996), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n998), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n966), .A2(new_n967), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n982), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n997), .A2(new_n999), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n966), .A2(new_n967), .A3(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n963), .A2(new_n1003), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n974), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n945), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n980), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n982), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n969), .A2(KEYINPUT106), .A3(new_n999), .A4(new_n997), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1000), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n966), .A2(new_n967), .A3(new_n1003), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(KEYINPUT107), .A3(new_n945), .A4(new_n1009), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n979), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n982), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1010), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(KEYINPUT43), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT44), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1018), .A2(new_n979), .A3(new_n945), .A4(new_n1009), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT43), .B1(new_n1010), .B2(new_n1021), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n1029), .ZN(G397));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n922), .A2(new_n923), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT45), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT108), .B(G40), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n472), .A2(new_n484), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G1996), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT46), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1036), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT109), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n925), .A2(new_n759), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n757), .A2(G2067), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n791), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1038), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(G1996), .B1(new_n787), .B2(new_n788), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1037), .A2(new_n791), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(KEYINPUT110), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT110), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(new_n841), .B(new_n845), .Z(new_n1058));
  NAND2_X1  g633(.A1(new_n1043), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G290), .A2(G1986), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1039), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT48), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1049), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT110), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n845), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(KEYINPUT126), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1054), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1044), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT127), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(KEYINPUT127), .A3(new_n1044), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1064), .B1(new_n1076), .B2(new_n1043), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n917), .A2(new_n920), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(KEYINPUT113), .A3(new_n1079), .A4(new_n1031), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1079), .B(new_n1031), .C1(new_n507), .C2(new_n514), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n472), .A2(new_n484), .A3(new_n1034), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1031), .B1(new_n507), .B2(new_n514), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(KEYINPUT50), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n764), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1033), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1033), .A2(G1384), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1078), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1091), .A3(new_n1035), .ZN(new_n1092));
  INV_X1    g667(.A(G1966), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1088), .A2(G168), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G8), .ZN(new_n1096));
  AND2_X1   g671(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(G8), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(G8), .A3(G286), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1098), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1105));
  NAND2_X1  g680(.A1(G303), .A2(G8), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1085), .B1(new_n1033), .B2(new_n1086), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n922), .A2(new_n923), .A3(new_n1090), .ZN(new_n1113));
  AOI21_X1  g688(.A(G1971), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1086), .A2(KEYINPUT50), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1115), .A2(new_n1035), .A3(new_n1081), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(G2090), .ZN(new_n1117));
  OAI21_X1  g692(.A(G8), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1111), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G2090), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1084), .A2(new_n1120), .A3(new_n1087), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1114), .B2(KEYINPUT112), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n1123), .B(G1971), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1124));
  OAI211_X1 g699(.A(G8), .B(new_n1110), .C1(new_n1122), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G8), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1086), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1035), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n809), .A2(G1976), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT52), .ZN(new_n1131));
  INV_X1    g706(.A(G1976), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(G288), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1128), .A2(new_n1129), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G305), .A2(G1981), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n831), .B1(new_n605), .B2(new_n606), .ZN(new_n1136));
  NOR2_X1   g711(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1137));
  OR3_X1    g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1137), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n1128), .A3(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1131), .A2(new_n1134), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1142));
  INV_X1    g717(.A(G1961), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1113), .A2(new_n766), .A3(new_n1035), .A4(new_n1089), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1142), .A2(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(G2078), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1112), .A2(new_n1091), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(G301), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  AND4_X1   g724(.A1(new_n1119), .A2(new_n1125), .A3(new_n1141), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1098), .A2(new_n1101), .A3(new_n1151), .A4(new_n1103), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1105), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1126), .B(G286), .C1(new_n1088), .C2(new_n1094), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1125), .A2(new_n1119), .A3(new_n1141), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(G8), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1111), .ZN(new_n1159));
  AND4_X1   g734(.A1(KEYINPUT63), .A2(new_n1102), .A3(G8), .A4(G168), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1159), .A2(new_n1125), .A3(new_n1141), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1125), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1140), .A2(new_n1132), .A3(new_n809), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1135), .B(KEYINPUT115), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1163), .A2(new_n1141), .B1(new_n1128), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1153), .A2(new_n1162), .A3(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT56), .B(G2072), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1112), .A2(new_n1113), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(G1956), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1116), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n957), .A2(KEYINPUT116), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT57), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT118), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1175), .B1(new_n1172), .B2(new_n1170), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT118), .ZN(new_n1181));
  AOI21_X1  g756(.A(G1348), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT117), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1035), .A2(new_n1127), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT117), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1185));
  AOI21_X1  g760(.A(G2067), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n624), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1179), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1175), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1189), .A2(KEYINPUT61), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1179), .A2(new_n1191), .A3(new_n1181), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT122), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1179), .A2(new_n1191), .A3(new_n1181), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1177), .A2(new_n1189), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1196), .A2(KEYINPUT121), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(KEYINPUT121), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1200));
  OAI211_X1 g775(.A(new_n1193), .B(new_n1195), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  NOR4_X1   g776(.A1(new_n1182), .A2(new_n1186), .A3(KEYINPUT60), .A4(new_n623), .ZN(new_n1202));
  OR3_X1    g777(.A1(new_n1182), .A2(new_n1186), .A3(new_n624), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1187), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1202), .B1(new_n1204), .B2(KEYINPUT60), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT59), .ZN(new_n1206));
  XNOR2_X1  g781(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(G1341), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1184), .A2(new_n1185), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(G1996), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1112), .A2(new_n1210), .A3(new_n1113), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT120), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1206), .B1(new_n1214), .B2(new_n566), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1216));
  AOI21_X1  g791(.A(KEYINPUT120), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1217));
  OAI211_X1 g792(.A(new_n1206), .B(new_n566), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1205), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1190), .B1(new_n1201), .B2(new_n1220), .ZN(new_n1221));
  AND3_X1   g796(.A1(new_n1125), .A2(new_n1119), .A3(new_n1141), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1223));
  XNOR2_X1  g798(.A(G301), .B(KEYINPUT54), .ZN(new_n1224));
  INV_X1    g799(.A(new_n467), .ZN(new_n1225));
  AND2_X1   g800(.A1(new_n1225), .A2(KEYINPUT125), .ZN(new_n1226));
  OAI21_X1  g801(.A(G2105), .B1(new_n1225), .B2(KEYINPUT125), .ZN(new_n1227));
  OAI211_X1 g802(.A(G40), .B(new_n1147), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g803(.A(new_n484), .B(KEYINPUT124), .ZN(new_n1229));
  AOI211_X1 g804(.A(new_n1228), .B(new_n1229), .C1(new_n936), .C2(new_n1090), .ZN(new_n1230));
  AND2_X1   g805(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1231));
  INV_X1    g806(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1224), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  AOI22_X1  g808(.A1(new_n1223), .A2(new_n1224), .B1(new_n1233), .B2(new_n1146), .ZN(new_n1234));
  AND3_X1   g809(.A1(new_n1222), .A2(new_n1104), .A3(new_n1234), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1168), .B1(new_n1221), .B2(new_n1235), .ZN(new_n1236));
  AND2_X1   g811(.A1(G290), .A2(G1986), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1039), .B1(new_n1060), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1057), .A2(new_n1059), .A3(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g814(.A(new_n1239), .B(KEYINPUT111), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1077), .B1(new_n1236), .B2(new_n1240), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g816(.A1(new_n685), .A2(G319), .A3(new_n668), .ZN(new_n1243));
  NOR2_X1   g817(.A1(G229), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g818(.A(new_n1027), .B(new_n1244), .C1(new_n947), .C2(new_n946), .ZN(G225));
  INV_X1    g819(.A(G225), .ZN(G308));
endmodule


