

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U325 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U326 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U327 ( .A(n452), .B(KEYINPUT84), .Z(n293) );
  XNOR2_X1 U328 ( .A(n420), .B(n419), .ZN(n448) );
  XNOR2_X1 U329 ( .A(n421), .B(n357), .ZN(n358) );
  XNOR2_X1 U330 ( .A(n359), .B(n358), .ZN(n360) );
  NOR2_X1 U331 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U332 ( .A(n437), .B(KEYINPUT124), .ZN(n438) );
  XNOR2_X1 U333 ( .A(n481), .B(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U334 ( .A(n439), .B(n438), .ZN(n459) );
  XNOR2_X1 U335 ( .A(KEYINPUT37), .B(n497), .ZN(n527) );
  XNOR2_X1 U336 ( .A(n460), .B(G176GAT), .ZN(n461) );
  XNOR2_X1 U337 ( .A(n462), .B(n461), .ZN(G1349GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n295) );
  XNOR2_X1 U339 ( .A(KEYINPUT32), .B(KEYINPUT69), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U341 ( .A(G148GAT), .B(G106GAT), .Z(n327) );
  XOR2_X1 U342 ( .A(n296), .B(n327), .Z(n299) );
  XOR2_X1 U343 ( .A(G85GAT), .B(G99GAT), .Z(n356) );
  XOR2_X1 U344 ( .A(G57GAT), .B(G71GAT), .Z(n297) );
  XNOR2_X1 U345 ( .A(KEYINPUT13), .B(n297), .ZN(n387) );
  XOR2_X1 U346 ( .A(n356), .B(n387), .Z(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n309) );
  XOR2_X1 U348 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n301) );
  XNOR2_X1 U349 ( .A(G120GAT), .B(G78GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n307) );
  XOR2_X1 U351 ( .A(G176GAT), .B(G204GAT), .Z(n303) );
  XNOR2_X1 U352 ( .A(G92GAT), .B(G64GAT), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n303), .B(n302), .ZN(n336) );
  XOR2_X1 U354 ( .A(n336), .B(KEYINPUT70), .Z(n305) );
  NAND2_X1 U355 ( .A1(G230GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U357 ( .A(n307), .B(n306), .Z(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n579) );
  XOR2_X1 U359 ( .A(KEYINPUT41), .B(n579), .Z(n559) );
  INV_X1 U360 ( .A(n559), .ZN(n544) );
  XOR2_X1 U361 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n311) );
  XNOR2_X1 U362 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U364 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n313) );
  XNOR2_X1 U365 ( .A(G211GAT), .B(KEYINPUT24), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U367 ( .A(n315), .B(n314), .Z(n326) );
  XOR2_X1 U368 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n317) );
  XNOR2_X1 U369 ( .A(KEYINPUT89), .B(G141GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U371 ( .A(KEYINPUT3), .B(n318), .Z(n435) );
  INV_X1 U372 ( .A(n435), .ZN(n324) );
  XOR2_X1 U373 ( .A(G197GAT), .B(KEYINPUT21), .Z(n320) );
  XNOR2_X1 U374 ( .A(G218GAT), .B(KEYINPUT88), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n340) );
  XOR2_X1 U376 ( .A(G204GAT), .B(n340), .Z(n322) );
  NAND2_X1 U377 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U379 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n328) );
  XOR2_X1 U381 ( .A(n328), .B(n327), .Z(n331) );
  XOR2_X1 U382 ( .A(G162GAT), .B(G50GAT), .Z(n348) );
  XNOR2_X1 U383 ( .A(G155GAT), .B(G22GAT), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n329), .B(G78GAT), .ZN(n395) );
  XNOR2_X1 U385 ( .A(n348), .B(n395), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n475) );
  XNOR2_X1 U387 ( .A(G183GAT), .B(G211GAT), .ZN(n332) );
  XOR2_X1 U388 ( .A(n332), .B(G8GAT), .Z(n388) );
  XNOR2_X1 U389 ( .A(G36GAT), .B(KEYINPUT76), .ZN(n333) );
  XNOR2_X1 U390 ( .A(n333), .B(G190GAT), .ZN(n363) );
  XOR2_X1 U391 ( .A(KEYINPUT97), .B(n363), .Z(n335) );
  NAND2_X1 U392 ( .A1(G226GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U394 ( .A(n337), .B(n336), .Z(n342) );
  XOR2_X1 U395 ( .A(G169GAT), .B(KEYINPUT19), .Z(n339) );
  XNOR2_X1 U396 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n453) );
  XNOR2_X1 U398 ( .A(n340), .B(n453), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n388), .B(n343), .ZN(n530) );
  XOR2_X1 U401 ( .A(KEYINPUT47), .B(KEYINPUT117), .Z(n402) );
  XOR2_X1 U402 ( .A(G106GAT), .B(KEYINPUT9), .Z(n345) );
  XNOR2_X1 U403 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n367) );
  XOR2_X1 U405 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n347) );
  XNOR2_X1 U406 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n349) );
  XOR2_X1 U408 ( .A(n349), .B(n348), .Z(n361) );
  INV_X1 U409 ( .A(KEYINPUT7), .ZN(n350) );
  NAND2_X1 U410 ( .A1(G43GAT), .A2(n350), .ZN(n353) );
  INV_X1 U411 ( .A(G43GAT), .ZN(n351) );
  NAND2_X1 U412 ( .A1(n351), .A2(KEYINPUT7), .ZN(n352) );
  NAND2_X1 U413 ( .A1(n353), .A2(n352), .ZN(n355) );
  XNOR2_X1 U414 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n374) );
  XOR2_X1 U416 ( .A(n356), .B(n374), .Z(n359) );
  XOR2_X1 U417 ( .A(KEYINPUT75), .B(G134GAT), .Z(n421) );
  NAND2_X1 U418 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XOR2_X1 U419 ( .A(n361), .B(n360), .Z(n365) );
  XNOR2_X1 U420 ( .A(KEYINPUT64), .B(G92GAT), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n565) );
  XOR2_X1 U422 ( .A(G113GAT), .B(G1GAT), .Z(n427) );
  XOR2_X1 U423 ( .A(G169GAT), .B(G15GAT), .Z(n369) );
  XNOR2_X1 U424 ( .A(G36GAT), .B(G50GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U426 ( .A(n427), .B(n370), .Z(n372) );
  NAND2_X1 U427 ( .A1(G229GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(n373), .B(KEYINPUT29), .Z(n376) );
  XNOR2_X1 U430 ( .A(n374), .B(KEYINPUT65), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n384) );
  XOR2_X1 U432 ( .A(G197GAT), .B(G22GAT), .Z(n378) );
  XNOR2_X1 U433 ( .A(G141GAT), .B(G8GAT), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U435 ( .A(KEYINPUT66), .B(KEYINPUT68), .Z(n380) );
  XNOR2_X1 U436 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U438 ( .A(n382), .B(n381), .Z(n383) );
  XOR2_X1 U439 ( .A(n384), .B(n383), .Z(n575) );
  INV_X1 U440 ( .A(n575), .ZN(n568) );
  NOR2_X1 U441 ( .A1(n544), .A2(n568), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n385), .B(KEYINPUT46), .ZN(n386) );
  NOR2_X1 U443 ( .A1(n565), .A2(n386), .ZN(n400) );
  XOR2_X1 U444 ( .A(n388), .B(n387), .Z(n399) );
  XOR2_X1 U445 ( .A(G127GAT), .B(G15GAT), .Z(n449) );
  XOR2_X1 U446 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n390) );
  XNOR2_X1 U447 ( .A(G1GAT), .B(G64GAT), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U449 ( .A(n449), .B(n391), .Z(n393) );
  NAND2_X1 U450 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U452 ( .A(n394), .B(KEYINPUT78), .Z(n397) );
  XNOR2_X1 U453 ( .A(n395), .B(KEYINPUT14), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n583) );
  XOR2_X1 U456 ( .A(KEYINPUT116), .B(n583), .Z(n571) );
  NAND2_X1 U457 ( .A1(n400), .A2(n571), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n408) );
  XNOR2_X1 U459 ( .A(n565), .B(KEYINPUT36), .ZN(n494) );
  NAND2_X1 U460 ( .A1(n494), .A2(n583), .ZN(n404) );
  XOR2_X1 U461 ( .A(KEYINPUT45), .B(KEYINPUT118), .Z(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n406) );
  NOR2_X1 U463 ( .A1(n579), .A2(n575), .ZN(n405) );
  AND2_X1 U464 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U465 ( .A(KEYINPUT48), .B(n409), .ZN(n554) );
  NOR2_X1 U466 ( .A1(n530), .A2(n554), .ZN(n412) );
  XOR2_X1 U467 ( .A(KEYINPUT123), .B(KEYINPUT54), .Z(n410) );
  XNOR2_X1 U468 ( .A(KEYINPUT122), .B(n410), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n436) );
  XOR2_X1 U470 ( .A(KEYINPUT94), .B(KEYINPUT6), .Z(n414) );
  XNOR2_X1 U471 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U473 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n416) );
  XNOR2_X1 U474 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U476 ( .A(n418), .B(n417), .Z(n433) );
  XOR2_X1 U477 ( .A(G120GAT), .B(KEYINPUT0), .Z(n420) );
  XNOR2_X1 U478 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n419) );
  XOR2_X1 U479 ( .A(n421), .B(n448), .Z(n423) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n431) );
  XOR2_X1 U482 ( .A(G155GAT), .B(G148GAT), .Z(n425) );
  XNOR2_X1 U483 ( .A(G85GAT), .B(G162GAT), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U485 ( .A(n426), .B(G127GAT), .Z(n429) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U490 ( .A(n435), .B(n434), .Z(n501) );
  INV_X1 U491 ( .A(n501), .ZN(n528) );
  NAND2_X1 U492 ( .A1(n436), .A2(n528), .ZN(n574) );
  NOR2_X1 U493 ( .A1(n475), .A2(n574), .ZN(n439) );
  INV_X1 U494 ( .A(KEYINPUT55), .ZN(n437) );
  XOR2_X1 U495 ( .A(KEYINPUT83), .B(KEYINPUT86), .Z(n441) );
  XNOR2_X1 U496 ( .A(G176GAT), .B(KEYINPUT82), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n458) );
  XOR2_X1 U498 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n443) );
  XNOR2_X1 U499 ( .A(G113GAT), .B(G183GAT), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U501 ( .A(G43GAT), .B(G99GAT), .Z(n445) );
  XNOR2_X1 U502 ( .A(G134GAT), .B(G190GAT), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n456) );
  XOR2_X1 U505 ( .A(n449), .B(n448), .Z(n451) );
  NAND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U508 ( .A(G71GAT), .B(n453), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n293), .B(n454), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X2 U511 ( .A(n458), .B(n457), .Z(n534) );
  INV_X1 U512 ( .A(n534), .ZN(n541) );
  NAND2_X1 U513 ( .A1(n459), .A2(n541), .ZN(n570) );
  NOR2_X1 U514 ( .A1(n544), .A2(n570), .ZN(n462) );
  XNOR2_X1 U515 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n460) );
  INV_X1 U516 ( .A(KEYINPUT58), .ZN(n465) );
  INV_X1 U517 ( .A(n565), .ZN(n551) );
  NOR2_X1 U518 ( .A1(n570), .A2(n551), .ZN(n463) );
  XNOR2_X1 U519 ( .A(G190GAT), .B(n463), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  NOR2_X1 U521 ( .A1(n579), .A2(n568), .ZN(n498) );
  NAND2_X1 U522 ( .A1(n534), .A2(n475), .ZN(n467) );
  XNOR2_X1 U523 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n467), .B(n466), .ZN(n573) );
  INV_X1 U525 ( .A(n530), .ZN(n504) );
  XOR2_X1 U526 ( .A(n504), .B(KEYINPUT27), .Z(n476) );
  NOR2_X1 U527 ( .A1(n573), .A2(n476), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT101), .ZN(n472) );
  NOR2_X1 U529 ( .A1(n534), .A2(n530), .ZN(n469) );
  NOR2_X1 U530 ( .A1(n475), .A2(n469), .ZN(n470) );
  XNOR2_X1 U531 ( .A(KEYINPUT25), .B(n470), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n473), .B(KEYINPUT102), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n474), .A2(n528), .ZN(n480) );
  XNOR2_X1 U535 ( .A(n475), .B(KEYINPUT28), .ZN(n513) );
  INV_X1 U536 ( .A(n513), .ZN(n537) );
  NOR2_X1 U537 ( .A1(n528), .A2(n476), .ZN(n477) );
  XNOR2_X1 U538 ( .A(KEYINPUT98), .B(n477), .ZN(n556) );
  NAND2_X1 U539 ( .A1(n537), .A2(n556), .ZN(n540) );
  NOR2_X1 U540 ( .A1(n541), .A2(n540), .ZN(n478) );
  XNOR2_X1 U541 ( .A(KEYINPUT99), .B(n478), .ZN(n479) );
  NAND2_X1 U542 ( .A1(n480), .A2(n479), .ZN(n481) );
  XOR2_X1 U543 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n483) );
  NAND2_X1 U544 ( .A1(n551), .A2(n583), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n484) );
  NOR2_X1 U546 ( .A1(n495), .A2(n484), .ZN(n515) );
  NAND2_X1 U547 ( .A1(n498), .A2(n515), .ZN(n492) );
  NOR2_X1 U548 ( .A1(n528), .A2(n492), .ZN(n485) );
  XOR2_X1 U549 ( .A(KEYINPUT34), .B(n485), .Z(n486) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  NOR2_X1 U551 ( .A1(n530), .A2(n492), .ZN(n487) );
  XOR2_X1 U552 ( .A(KEYINPUT104), .B(n487), .Z(n488) );
  XNOR2_X1 U553 ( .A(G8GAT), .B(n488), .ZN(G1325GAT) );
  NOR2_X1 U554 ( .A1(n534), .A2(n492), .ZN(n490) );
  XNOR2_X1 U555 ( .A(KEYINPUT105), .B(KEYINPUT35), .ZN(n489) );
  XNOR2_X1 U556 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U557 ( .A(G15GAT), .B(n491), .Z(G1326GAT) );
  NOR2_X1 U558 ( .A1(n537), .A2(n492), .ZN(n493) );
  XOR2_X1 U559 ( .A(G22GAT), .B(n493), .Z(G1327GAT) );
  XOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .Z(n503) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(KEYINPUT38), .Z(n500) );
  NOR2_X1 U562 ( .A1(n583), .A2(n495), .ZN(n496) );
  NAND2_X1 U563 ( .A1(n494), .A2(n496), .ZN(n497) );
  NAND2_X1 U564 ( .A1(n498), .A2(n527), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n512) );
  NAND2_X1 U566 ( .A1(n512), .A2(n501), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  XOR2_X1 U568 ( .A(G36GAT), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U569 ( .A1(n512), .A2(n504), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(G1329GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT40), .B(KEYINPUT110), .Z(n508) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(KEYINPUT109), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n511) );
  NAND2_X1 U574 ( .A1(n512), .A2(n541), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1330GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U579 ( .A1(n575), .A2(n544), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n526), .A2(n515), .ZN(n523) );
  NOR2_X1 U581 ( .A1(n528), .A2(n523), .ZN(n520) );
  XOR2_X1 U582 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n517) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(KEYINPUT111), .B(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1332GAT) );
  NOR2_X1 U587 ( .A1(n530), .A2(n523), .ZN(n521) );
  XOR2_X1 U588 ( .A(G64GAT), .B(n521), .Z(G1333GAT) );
  NOR2_X1 U589 ( .A1(n534), .A2(n523), .ZN(n522) );
  XOR2_X1 U590 ( .A(G71GAT), .B(n522), .Z(G1334GAT) );
  NOR2_X1 U591 ( .A1(n537), .A2(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n536) );
  NOR2_X1 U595 ( .A1(n528), .A2(n536), .ZN(n529) );
  XOR2_X1 U596 ( .A(G85GAT), .B(n529), .Z(G1336GAT) );
  NOR2_X1 U597 ( .A1(n530), .A2(n536), .ZN(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G92GAT), .B(n533), .ZN(G1337GAT) );
  NOR2_X1 U601 ( .A1(n534), .A2(n536), .ZN(n535) );
  XOR2_X1 U602 ( .A(G99GAT), .B(n535), .Z(G1338GAT) );
  NOR2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U604 ( .A(KEYINPUT44), .B(n538), .Z(n539) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  NOR2_X1 U606 ( .A1(n540), .A2(n554), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n568), .A2(n550), .ZN(n543) );
  XOR2_X1 U609 ( .A(G113GAT), .B(n543), .Z(G1340GAT) );
  NOR2_X1 U610 ( .A1(n544), .A2(n550), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NOR2_X1 U613 ( .A1(n571), .A2(n550), .ZN(n548) );
  XNOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NOR2_X1 U620 ( .A1(n573), .A2(n554), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(n557), .Z(n566) );
  NAND2_X1 U623 ( .A1(n566), .A2(n575), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT53), .Z(n561) );
  NAND2_X1 U626 ( .A1(n566), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n583), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n570), .ZN(n569) );
  XOR2_X1 U635 ( .A(G169GAT), .B(n569), .Z(G1348GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U637 ( .A(G183GAT), .B(n572), .Z(G1350GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n577) );
  NOR2_X1 U639 ( .A1(n573), .A2(n574), .ZN(n587) );
  NAND2_X1 U640 ( .A1(n587), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U644 ( .A1(n587), .A2(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n585) );
  NAND2_X1 U648 ( .A1(n587), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  NAND2_X1 U651 ( .A1(n587), .A2(n494), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

