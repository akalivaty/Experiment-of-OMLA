

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U554 ( .A(KEYINPUT29), .B(n729), .Z(n521) );
  XNOR2_X2 U555 ( .A(n690), .B(KEYINPUT94), .ZN(n731) );
  INV_X1 U556 ( .A(G2105), .ZN(n528) );
  NOR2_X1 U557 ( .A1(n684), .A2(n683), .ZN(n686) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n680) );
  XOR2_X1 U559 ( .A(KEYINPUT65), .B(n533), .Z(n642) );
  NAND2_X1 U560 ( .A1(n522), .A2(n826), .ZN(n816) );
  AND2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n892) );
  AND2_X1 U562 ( .A1(n820), .A2(n803), .ZN(n522) );
  INV_X1 U563 ( .A(KEYINPUT96), .ZN(n708) );
  XNOR2_X1 U564 ( .A(n709), .B(n708), .ZN(n715) );
  INV_X1 U565 ( .A(KEYINPUT97), .ZN(n692) );
  XNOR2_X1 U566 ( .A(n695), .B(KEYINPUT30), .ZN(n696) );
  INV_X1 U567 ( .A(KEYINPUT31), .ZN(n699) );
  INV_X1 U568 ( .A(G40), .ZN(n681) );
  OR2_X1 U569 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U570 ( .A(KEYINPUT12), .B(KEYINPUT70), .ZN(n563) );
  INV_X1 U571 ( .A(KEYINPUT88), .ZN(n685) );
  XNOR2_X1 U572 ( .A(n564), .B(n563), .ZN(n566) );
  XNOR2_X1 U573 ( .A(n686), .B(n685), .ZN(n798) );
  INV_X1 U574 ( .A(KEYINPUT17), .ZN(n523) );
  XNOR2_X1 U575 ( .A(KEYINPUT71), .B(n588), .ZN(n1027) );
  NOR2_X1 U576 ( .A1(G651), .A2(n629), .ZN(n641) );
  AND2_X2 U577 ( .A1(n528), .A2(G2104), .ZN(n895) );
  INV_X1 U578 ( .A(n1013), .ZN(n703) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n629) );
  NAND2_X1 U580 ( .A1(n896), .A2(G138), .ZN(n525) );
  NOR2_X2 U581 ( .A1(n572), .A2(n571), .ZN(n1013) );
  AND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(G164) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XNOR2_X2 U584 ( .A(n524), .B(n523), .ZN(n896) );
  XNOR2_X1 U585 ( .A(n525), .B(KEYINPUT86), .ZN(n532) );
  NAND2_X1 U586 ( .A1(G102), .A2(n895), .ZN(n527) );
  NAND2_X1 U587 ( .A1(G114), .A2(n892), .ZN(n526) );
  NAND2_X1 U588 ( .A1(n527), .A2(n526), .ZN(n530) );
  NOR2_X2 U589 ( .A1(G2104), .A2(n528), .ZN(n891) );
  AND2_X1 U590 ( .A1(G126), .A2(n891), .ZN(n529) );
  NOR2_X1 U591 ( .A1(n530), .A2(n529), .ZN(n531) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G108), .ZN(G238) );
  INV_X1 U594 ( .A(G120), .ZN(G236) );
  INV_X1 U595 ( .A(G57), .ZN(G237) );
  INV_X1 U596 ( .A(G82), .ZN(G220) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n533) );
  NAND2_X1 U598 ( .A1(G88), .A2(n642), .ZN(n536) );
  INV_X1 U599 ( .A(G651), .ZN(n537) );
  OR2_X1 U600 ( .A1(n537), .A2(n629), .ZN(n534) );
  XOR2_X1 U601 ( .A(KEYINPUT66), .B(n534), .Z(n643) );
  NAND2_X1 U602 ( .A1(G75), .A2(n643), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n542) );
  NOR2_X1 U604 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n538), .Z(n646) );
  NAND2_X1 U606 ( .A1(G62), .A2(n646), .ZN(n540) );
  NAND2_X1 U607 ( .A1(G50), .A2(n641), .ZN(n539) );
  NAND2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(G166) );
  NAND2_X1 U610 ( .A1(G76), .A2(n643), .ZN(n543) );
  XNOR2_X1 U611 ( .A(KEYINPUT74), .B(n543), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT73), .B(KEYINPUT4), .Z(n545) );
  NAND2_X1 U613 ( .A1(G89), .A2(n642), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(KEYINPUT5), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n646), .A2(G63), .ZN(n549) );
  XOR2_X1 U618 ( .A(KEYINPUT75), .B(n549), .Z(n551) );
  NAND2_X1 U619 ( .A1(n641), .A2(G51), .ZN(n550) );
  NAND2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U621 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(n896), .A2(G137), .ZN(n558) );
  NAND2_X1 U626 ( .A1(G101), .A2(n895), .ZN(n556) );
  XOR2_X1 U627 ( .A(KEYINPUT23), .B(n556), .Z(n557) );
  NAND2_X1 U628 ( .A1(n558), .A2(n557), .ZN(n684) );
  NAND2_X1 U629 ( .A1(G125), .A2(n891), .ZN(n560) );
  NAND2_X1 U630 ( .A1(G113), .A2(n892), .ZN(n559) );
  NAND2_X1 U631 ( .A1(n560), .A2(n559), .ZN(n682) );
  NOR2_X1 U632 ( .A1(n684), .A2(n682), .ZN(G160) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U634 ( .A(n561), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U635 ( .A(G567), .ZN(n675) );
  NOR2_X1 U636 ( .A1(n675), .A2(G223), .ZN(n562) );
  XNOR2_X1 U637 ( .A(n562), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U638 ( .A1(G81), .A2(n642), .ZN(n564) );
  NAND2_X1 U639 ( .A1(G68), .A2(n643), .ZN(n565) );
  NAND2_X1 U640 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U641 ( .A(n567), .B(KEYINPUT13), .ZN(n569) );
  NAND2_X1 U642 ( .A1(G43), .A2(n641), .ZN(n568) );
  NAND2_X1 U643 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n646), .A2(G56), .ZN(n570) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n570), .Z(n571) );
  NAND2_X1 U646 ( .A1(n1013), .A2(G860), .ZN(G153) );
  NAND2_X1 U647 ( .A1(G64), .A2(n646), .ZN(n574) );
  NAND2_X1 U648 ( .A1(G52), .A2(n641), .ZN(n573) );
  AND2_X1 U649 ( .A1(n574), .A2(n573), .ZN(n580) );
  XNOR2_X1 U650 ( .A(KEYINPUT9), .B(KEYINPUT68), .ZN(n578) );
  NAND2_X1 U651 ( .A1(G90), .A2(n642), .ZN(n576) );
  NAND2_X1 U652 ( .A1(G77), .A2(n643), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U654 ( .A(n578), .B(n577), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n580), .A2(n579), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G66), .A2(n646), .ZN(n582) );
  NAND2_X1 U657 ( .A1(G92), .A2(n642), .ZN(n581) );
  NAND2_X1 U658 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n643), .A2(G79), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n641), .A2(G54), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U662 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n587), .Z(n588) );
  INV_X1 U664 ( .A(G868), .ZN(n660) );
  NAND2_X1 U665 ( .A1(n1027), .A2(n660), .ZN(n589) );
  XNOR2_X1 U666 ( .A(n589), .B(KEYINPUT72), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U669 ( .A1(G65), .A2(n646), .ZN(n593) );
  NAND2_X1 U670 ( .A1(G53), .A2(n641), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U672 ( .A1(G91), .A2(n642), .ZN(n595) );
  NAND2_X1 U673 ( .A1(G78), .A2(n643), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n1026) );
  INV_X1 U676 ( .A(n1026), .ZN(G299) );
  NOR2_X1 U677 ( .A1(G286), .A2(n660), .ZN(n598) );
  XNOR2_X1 U678 ( .A(n598), .B(KEYINPUT76), .ZN(n600) );
  NOR2_X1 U679 ( .A1(G299), .A2(G868), .ZN(n599) );
  NOR2_X1 U680 ( .A1(n600), .A2(n599), .ZN(G297) );
  INV_X1 U681 ( .A(G559), .ZN(n601) );
  NOR2_X1 U682 ( .A1(G860), .A2(n601), .ZN(n602) );
  XNOR2_X1 U683 ( .A(KEYINPUT77), .B(n602), .ZN(n603) );
  INV_X1 U684 ( .A(n1027), .ZN(n639) );
  NAND2_X1 U685 ( .A1(n603), .A2(n639), .ZN(n604) );
  XNOR2_X1 U686 ( .A(n604), .B(KEYINPUT16), .ZN(n605) );
  XNOR2_X1 U687 ( .A(KEYINPUT78), .B(n605), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G868), .A2(n703), .ZN(n608) );
  NAND2_X1 U689 ( .A1(G868), .A2(n639), .ZN(n606) );
  NOR2_X1 U690 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G99), .A2(n895), .ZN(n610) );
  NAND2_X1 U693 ( .A1(G111), .A2(n892), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U695 ( .A(n611), .B(KEYINPUT79), .ZN(n613) );
  NAND2_X1 U696 ( .A1(G135), .A2(n896), .ZN(n612) );
  NAND2_X1 U697 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n891), .A2(G123), .ZN(n614) );
  XOR2_X1 U699 ( .A(KEYINPUT18), .B(n614), .Z(n615) );
  NOR2_X1 U700 ( .A1(n616), .A2(n615), .ZN(n935) );
  XNOR2_X1 U701 ( .A(G2096), .B(n935), .ZN(n618) );
  INV_X1 U702 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U703 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G85), .A2(n642), .ZN(n620) );
  NAND2_X1 U705 ( .A1(G47), .A2(n641), .ZN(n619) );
  NAND2_X1 U706 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U707 ( .A1(G72), .A2(n643), .ZN(n622) );
  NAND2_X1 U708 ( .A1(n646), .A2(G60), .ZN(n621) );
  NAND2_X1 U709 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U711 ( .A(n625), .B(KEYINPUT67), .ZN(G290) );
  NAND2_X1 U712 ( .A1(G49), .A2(n641), .ZN(n627) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U714 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U715 ( .A1(n646), .A2(n628), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n629), .A2(G87), .ZN(n630) );
  NAND2_X1 U717 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G86), .A2(n642), .ZN(n633) );
  NAND2_X1 U719 ( .A1(G48), .A2(n641), .ZN(n632) );
  NAND2_X1 U720 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n643), .A2(G73), .ZN(n634) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n634), .Z(n635) );
  NOR2_X1 U723 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U724 ( .A1(n646), .A2(G61), .ZN(n637) );
  NAND2_X1 U725 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G559), .A2(n639), .ZN(n640) );
  XNOR2_X1 U727 ( .A(n640), .B(n703), .ZN(n845) );
  NAND2_X1 U728 ( .A1(G55), .A2(n641), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G93), .A2(n642), .ZN(n645) );
  NAND2_X1 U730 ( .A1(G80), .A2(n643), .ZN(n644) );
  NAND2_X1 U731 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n646), .A2(G67), .ZN(n647) );
  XOR2_X1 U733 ( .A(KEYINPUT80), .B(n647), .Z(n648) );
  NOR2_X1 U734 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U736 ( .A(n652), .B(KEYINPUT81), .Z(n846) );
  XOR2_X1 U737 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n653) );
  XNOR2_X1 U738 ( .A(G288), .B(n653), .ZN(n654) );
  XNOR2_X1 U739 ( .A(G166), .B(n654), .ZN(n656) );
  XNOR2_X1 U740 ( .A(G305), .B(n1026), .ZN(n655) );
  XNOR2_X1 U741 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U742 ( .A(n846), .B(n657), .ZN(n658) );
  XNOR2_X1 U743 ( .A(G290), .B(n658), .ZN(n919) );
  XNOR2_X1 U744 ( .A(n845), .B(n919), .ZN(n659) );
  NAND2_X1 U745 ( .A1(n659), .A2(G868), .ZN(n662) );
  NAND2_X1 U746 ( .A1(n660), .A2(n846), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n664), .ZN(n666) );
  XOR2_X1 U751 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n665) );
  XNOR2_X1 U752 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U753 ( .A1(n667), .A2(G2072), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n668), .B(KEYINPUT84), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U756 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U759 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U760 ( .A1(G96), .A2(n671), .ZN(n842) );
  NAND2_X1 U761 ( .A1(G2106), .A2(n842), .ZN(n672) );
  XNOR2_X1 U762 ( .A(n672), .B(KEYINPUT85), .ZN(n677) );
  NOR2_X1 U763 ( .A1(G236), .A2(G238), .ZN(n673) );
  NAND2_X1 U764 ( .A1(G69), .A2(n673), .ZN(n674) );
  NOR2_X1 U765 ( .A1(G237), .A2(n674), .ZN(n844) );
  NOR2_X1 U766 ( .A1(n675), .A2(n844), .ZN(n676) );
  NOR2_X1 U767 ( .A1(n677), .A2(n676), .ZN(G319) );
  INV_X1 U768 ( .A(G319), .ZN(n679) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U770 ( .A1(n679), .A2(n678), .ZN(n841) );
  NAND2_X1 U771 ( .A1(n841), .A2(G36), .ZN(G176) );
  INV_X1 U772 ( .A(G166), .ZN(G303) );
  INV_X1 U773 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U774 ( .A(n680), .B(KEYINPUT64), .ZN(n799) );
  XNOR2_X1 U775 ( .A(KEYINPUT93), .B(n798), .ZN(n687) );
  NAND2_X1 U776 ( .A1(n799), .A2(n687), .ZN(n691) );
  INV_X1 U777 ( .A(G1961), .ZN(n974) );
  NAND2_X1 U778 ( .A1(n691), .A2(n974), .ZN(n689) );
  INV_X1 U779 ( .A(n691), .ZN(n720) );
  XNOR2_X1 U780 ( .A(KEYINPUT25), .B(G2078), .ZN(n995) );
  NAND2_X1 U781 ( .A1(n720), .A2(n995), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n702) );
  NOR2_X1 U783 ( .A1(G171), .A2(n702), .ZN(n698) );
  NAND2_X1 U784 ( .A1(n691), .A2(G8), .ZN(n690) );
  NOR2_X1 U785 ( .A1(n731), .A2(G1966), .ZN(n748) );
  BUF_X1 U786 ( .A(n691), .Z(n732) );
  NOR2_X1 U787 ( .A1(G2084), .A2(n732), .ZN(n745) );
  NOR2_X1 U788 ( .A1(n748), .A2(n745), .ZN(n693) );
  XNOR2_X1 U789 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n694), .A2(G8), .ZN(n695) );
  NOR2_X1 U791 ( .A1(G168), .A2(n696), .ZN(n697) );
  NOR2_X1 U792 ( .A1(n698), .A2(n697), .ZN(n700) );
  XNOR2_X1 U793 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U794 ( .A(n701), .B(KEYINPUT98), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n702), .A2(G171), .ZN(n730) );
  NOR2_X1 U796 ( .A1(n1027), .A2(n703), .ZN(n710) );
  AND2_X1 U797 ( .A1(n720), .A2(G1996), .ZN(n705) );
  XNOR2_X1 U798 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n704) );
  XNOR2_X1 U799 ( .A(n705), .B(n704), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n732), .A2(G1341), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n710), .A2(n715), .ZN(n714) );
  NOR2_X1 U803 ( .A1(n720), .A2(G1348), .ZN(n712) );
  NOR2_X1 U804 ( .A1(G2067), .A2(n732), .ZN(n711) );
  NOR2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n715), .A2(n1013), .ZN(n716) );
  NAND2_X1 U808 ( .A1(n716), .A2(n1027), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n724) );
  NAND2_X1 U810 ( .A1(n720), .A2(G2072), .ZN(n719) );
  XNOR2_X1 U811 ( .A(n719), .B(KEYINPUT27), .ZN(n722) );
  INV_X1 U812 ( .A(G1956), .ZN(n962) );
  NOR2_X1 U813 ( .A1(n962), .A2(n720), .ZN(n721) );
  NOR2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n1026), .A2(n725), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U817 ( .A1(n1026), .A2(n725), .ZN(n726) );
  XOR2_X1 U818 ( .A(n726), .B(KEYINPUT28), .Z(n727) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n730), .A2(n521), .ZN(n747) );
  INV_X1 U821 ( .A(G8), .ZN(n737) );
  NOR2_X1 U822 ( .A1(n731), .A2(G1971), .ZN(n734) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U825 ( .A1(n735), .A2(G303), .ZN(n736) );
  OR2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n739) );
  AND2_X1 U827 ( .A1(n747), .A2(n739), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n746), .A2(n738), .ZN(n743) );
  INV_X1 U829 ( .A(n739), .ZN(n741) );
  AND2_X1 U830 ( .A1(G286), .A2(G8), .ZN(n740) );
  OR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U833 ( .A(n744), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U834 ( .A1(G8), .A2(n745), .ZN(n751) );
  AND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n749) );
  NOR2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n753), .A2(n752), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n764), .B(KEYINPUT99), .ZN(n757) );
  NAND2_X1 U840 ( .A1(G8), .A2(G166), .ZN(n754) );
  NOR2_X1 U841 ( .A1(G2090), .A2(n754), .ZN(n755) );
  XOR2_X1 U842 ( .A(KEYINPUT101), .B(n755), .Z(n756) );
  NOR2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n758) );
  INV_X1 U844 ( .A(n731), .ZN(n767) );
  NOR2_X1 U845 ( .A1(n758), .A2(n767), .ZN(n759) );
  INV_X1 U846 ( .A(n759), .ZN(n763) );
  NOR2_X1 U847 ( .A1(G1981), .A2(G305), .ZN(n760) );
  XNOR2_X1 U848 ( .A(n760), .B(KEYINPUT24), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n761), .A2(n767), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n782) );
  XOR2_X1 U851 ( .A(KEYINPUT99), .B(n764), .Z(n773) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n765) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n1032) );
  XNOR2_X1 U855 ( .A(KEYINPUT100), .B(n1032), .ZN(n771) );
  AND2_X1 U856 ( .A1(n766), .A2(KEYINPUT33), .ZN(n768) );
  AND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U858 ( .A(G1981), .B(G305), .ZN(n1017) );
  NOR2_X1 U859 ( .A1(n769), .A2(n1017), .ZN(n775) );
  AND2_X1 U860 ( .A1(n775), .A2(KEYINPUT33), .ZN(n778) );
  INV_X1 U861 ( .A(n778), .ZN(n770) );
  AND2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n780) );
  NAND2_X1 U864 ( .A1(G1976), .A2(G288), .ZN(n1025) );
  INV_X1 U865 ( .A(n1025), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n731), .A2(n774), .ZN(n776) );
  AND2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  OR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  AND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n817) );
  NAND2_X1 U871 ( .A1(G141), .A2(n896), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G117), .A2(n892), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n895), .A2(G105), .ZN(n785) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(n785), .Z(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n891), .A2(G129), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n904) );
  NAND2_X1 U879 ( .A1(G1996), .A2(n904), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G95), .A2(n895), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G107), .A2(n892), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G131), .A2(n896), .ZN(n793) );
  NAND2_X1 U884 ( .A1(G119), .A2(n891), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n794) );
  OR2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n905) );
  NAND2_X1 U887 ( .A1(G1991), .A2(n905), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n942) );
  NOR2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n831) );
  NAND2_X1 U890 ( .A1(n942), .A2(n831), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n800), .B(KEYINPUT92), .ZN(n820) );
  XNOR2_X1 U892 ( .A(G1986), .B(KEYINPUT87), .ZN(n801) );
  XNOR2_X1 U893 ( .A(n801), .B(G290), .ZN(n1023) );
  INV_X1 U894 ( .A(n831), .ZN(n814) );
  NOR2_X1 U895 ( .A1(n1023), .A2(n814), .ZN(n802) );
  XNOR2_X1 U896 ( .A(n802), .B(KEYINPUT89), .ZN(n803) );
  NAND2_X1 U897 ( .A1(G128), .A2(n891), .ZN(n805) );
  NAND2_X1 U898 ( .A1(G116), .A2(n892), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U900 ( .A(KEYINPUT35), .B(n806), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n895), .A2(G104), .ZN(n807) );
  XNOR2_X1 U902 ( .A(n807), .B(KEYINPUT90), .ZN(n809) );
  NAND2_X1 U903 ( .A1(G140), .A2(n896), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U905 ( .A(KEYINPUT34), .B(n810), .Z(n811) );
  NAND2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U907 ( .A(KEYINPUT36), .B(n813), .Z(n916) );
  XNOR2_X1 U908 ( .A(G2067), .B(KEYINPUT37), .ZN(n828) );
  OR2_X1 U909 ( .A1(n916), .A2(n828), .ZN(n936) );
  NOR2_X1 U910 ( .A1(n936), .A2(n814), .ZN(n815) );
  XNOR2_X1 U911 ( .A(n815), .B(KEYINPUT91), .ZN(n826) );
  OR2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U913 ( .A(n818), .B(KEYINPUT102), .ZN(n834) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n904), .ZN(n946) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n905), .ZN(n938) );
  NOR2_X1 U917 ( .A1(n819), .A2(n938), .ZN(n822) );
  INV_X1 U918 ( .A(n820), .ZN(n821) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U920 ( .A(KEYINPUT103), .B(n823), .Z(n824) );
  NOR2_X1 U921 ( .A1(n946), .A2(n824), .ZN(n825) );
  XNOR2_X1 U922 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n916), .A2(n828), .ZN(n943) );
  NAND2_X1 U925 ( .A1(n829), .A2(n943), .ZN(n830) );
  XNOR2_X1 U926 ( .A(KEYINPUT104), .B(n830), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n835), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U930 ( .A(G223), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n836), .A2(G2106), .ZN(n837) );
  XNOR2_X1 U932 ( .A(n837), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U934 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n839) );
  XOR2_X1 U936 ( .A(KEYINPUT107), .B(n839), .Z(n840) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(n842), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(G261) );
  INV_X1 U942 ( .A(G261), .ZN(G325) );
  NOR2_X1 U943 ( .A1(n845), .A2(G860), .ZN(n847) );
  XOR2_X1 U944 ( .A(n847), .B(n846), .Z(G145) );
  XNOR2_X1 U945 ( .A(G1341), .B(G2454), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n848), .B(G2430), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n849), .B(G1348), .ZN(n855) );
  XOR2_X1 U948 ( .A(G2443), .B(G2427), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2438), .B(G2446), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U951 ( .A(G2451), .B(G2435), .Z(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  NAND2_X1 U954 ( .A1(n856), .A2(G14), .ZN(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT105), .B(n857), .ZN(G401) );
  XOR2_X1 U956 ( .A(G1956), .B(G1966), .Z(n859) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1981), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U959 ( .A(G1976), .B(G1971), .Z(n861) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1961), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U962 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U963 ( .A(G2474), .B(KEYINPUT109), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n867) );
  XOR2_X1 U965 ( .A(G1991), .B(KEYINPUT41), .Z(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(G229) );
  XOR2_X1 U967 ( .A(G2096), .B(KEYINPUT43), .Z(n869) );
  XNOR2_X1 U968 ( .A(G2090), .B(G2678), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U970 ( .A(n870), .B(KEYINPUT108), .Z(n872) );
  XNOR2_X1 U971 ( .A(G2067), .B(G2072), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U973 ( .A(KEYINPUT42), .B(G2100), .Z(n874) );
  XNOR2_X1 U974 ( .A(G2084), .B(G2078), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(G227) );
  NAND2_X1 U977 ( .A1(G124), .A2(n891), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n877), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n895), .A2(G100), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G136), .A2(n896), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G112), .A2(n892), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(G162) );
  XNOR2_X1 U985 ( .A(G164), .B(n935), .ZN(n915) );
  NAND2_X1 U986 ( .A1(G103), .A2(n895), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G139), .A2(n896), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G127), .A2(n891), .ZN(n887) );
  NAND2_X1 U990 ( .A1(G115), .A2(n892), .ZN(n886) );
  NAND2_X1 U991 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n930) );
  XNOR2_X1 U994 ( .A(n930), .B(G162), .ZN(n903) );
  NAND2_X1 U995 ( .A1(G130), .A2(n891), .ZN(n894) );
  NAND2_X1 U996 ( .A1(G118), .A2(n892), .ZN(n893) );
  NAND2_X1 U997 ( .A1(n894), .A2(n893), .ZN(n901) );
  NAND2_X1 U998 ( .A1(G106), .A2(n895), .ZN(n898) );
  NAND2_X1 U999 ( .A1(G142), .A2(n896), .ZN(n897) );
  NAND2_X1 U1000 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U1001 ( .A(KEYINPUT45), .B(n899), .Z(n900) );
  NOR2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(G160), .B(n904), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1006 ( .A(n908), .B(n907), .Z(n913) );
  XOR2_X1 U1007 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n910) );
  XNOR2_X1 U1008 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT110), .B(n911), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1013 ( .A(n917), .B(n916), .Z(n918) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n918), .ZN(G395) );
  XNOR2_X1 U1015 ( .A(G286), .B(n919), .ZN(n921) );
  XNOR2_X1 U1016 ( .A(n1027), .B(n1013), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n922), .B(G301), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n923), .ZN(G397) );
  NOR2_X1 U1020 ( .A1(G229), .A2(G227), .ZN(n924) );
  XOR2_X1 U1021 ( .A(KEYINPUT49), .B(n924), .Z(n925) );
  NAND2_X1 U1022 ( .A1(G319), .A2(n925), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(G401), .A2(n926), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n927) );
  XOR2_X1 U1025 ( .A(KEYINPUT113), .B(n927), .Z(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1029 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n933), .Z(n952) );
  XOR2_X1 U1033 ( .A(G2084), .B(G160), .Z(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT114), .B(n940), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n949) );
  XOR2_X1 U1040 ( .A(G2090), .B(G162), .Z(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n947), .B(KEYINPUT51), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT115), .B(n950), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1046 ( .A(n953), .B(KEYINPUT116), .Z(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n954), .ZN(n955) );
  NOR2_X1 U1048 ( .A1(KEYINPUT55), .A2(n955), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT117), .B(n956), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(G29), .ZN(n1012) );
  XOR2_X1 U1051 ( .A(G1966), .B(G21), .Z(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT125), .B(n958), .ZN(n972) );
  XOR2_X1 U1053 ( .A(G4), .B(KEYINPUT124), .Z(n960) );
  XNOR2_X1 U1054 ( .A(G1348), .B(KEYINPUT59), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(n960), .B(n959), .ZN(n969) );
  XNOR2_X1 U1056 ( .A(G1341), .B(G19), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n961), .B(KEYINPUT122), .ZN(n966) );
  XOR2_X1 U1058 ( .A(G1981), .B(G6), .Z(n964) );
  XNOR2_X1 U1059 ( .A(n962), .B(G20), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n967), .B(KEYINPUT123), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1064 ( .A(KEYINPUT60), .B(n970), .Z(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT126), .B(n973), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n974), .B(G5), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n984) );
  XNOR2_X1 U1069 ( .A(G1971), .B(G22), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G23), .B(G1976), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G1986), .B(KEYINPUT127), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(n979), .B(G24), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(KEYINPUT58), .B(n982), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1077 ( .A(KEYINPUT61), .B(n985), .Z(n986) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n986), .ZN(n1010) );
  XOR2_X1 U1079 ( .A(G29), .B(KEYINPUT120), .Z(n1007) );
  XNOR2_X1 U1080 ( .A(G1996), .B(G32), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(G33), .B(G2072), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n994) );
  XOR2_X1 U1083 ( .A(G2067), .B(G26), .Z(n989) );
  NAND2_X1 U1084 ( .A1(n989), .A2(G28), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G25), .B(G1991), .ZN(n990) );
  XNOR2_X1 U1086 ( .A(KEYINPUT118), .B(n990), .ZN(n991) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1089 ( .A(G27), .B(n995), .Z(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(n998), .B(KEYINPUT119), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(n999), .B(KEYINPUT53), .ZN(n1002) );
  XOR2_X1 U1093 ( .A(G2084), .B(G34), .Z(n1000) );
  XNOR2_X1 U1094 ( .A(KEYINPUT54), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1096 ( .A(G35), .B(G2090), .ZN(n1003) );
  NOR2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1098 ( .A(n1005), .B(KEYINPUT55), .ZN(n1006) );
  NAND2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1100 ( .A1(G11), .A2(n1008), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1039) );
  XOR2_X1 U1103 ( .A(KEYINPUT56), .B(G16), .Z(n1037) );
  XNOR2_X1 U1104 ( .A(n1013), .B(G1341), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(G171), .B(G1961), .ZN(n1014) );
  NAND2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(G168), .B(G1966), .Z(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1109 ( .A(KEYINPUT121), .B(n1018), .Z(n1019) );
  XNOR2_X1 U1110 ( .A(n1019), .B(KEYINPUT57), .ZN(n1020) );
  NOR2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1035) );
  NAND2_X1 U1113 ( .A1(G1971), .A2(G303), .ZN(n1024) );
  NAND2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(n1026), .B(G1956), .ZN(n1029) );
  XOR2_X1 U1116 ( .A(G1348), .B(n1027), .Z(n1028) );
  NAND2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  NAND2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1122 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1123 ( .A(n1040), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

