//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n189), .A2(new_n190), .B1(G134), .B2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(G134), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(G131), .B1(new_n192), .B2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n194), .B1(new_n199), .B2(new_n193), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  XNOR2_X1  g015(.A(G134), .B(G137), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n200), .B(new_n201), .C1(new_n193), .C2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  OR2_X1    g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n205), .B(new_n206), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT65), .B1(new_n207), .B2(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n209), .A3(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(new_n205), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n211), .A2(new_n217), .A3(KEYINPUT70), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n204), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G116), .B(G119), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT69), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT2), .B(G113), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G119), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G116), .ZN(new_n231));
  OAI211_X1 g045(.A(KEYINPUT68), .B(new_n227), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n225), .A2(new_n226), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n226), .B1(new_n225), .B2(new_n232), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n208), .A2(new_n210), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n209), .A2(G143), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n236), .B1(new_n240), .B2(KEYINPUT1), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n238), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n202), .A2(new_n201), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n203), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n222), .A2(new_n235), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(G237), .A2(G953), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT27), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n218), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n211), .A2(new_n217), .A3(KEYINPUT66), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n204), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n244), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n244), .A2(KEYINPUT30), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n235), .B1(new_n260), .B2(new_n222), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n251), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n188), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n235), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n204), .A2(new_n220), .A3(new_n221), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n244), .A2(KEYINPUT30), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n257), .B1(new_n255), .B2(new_n244), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n245), .B(new_n250), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n245), .A2(KEYINPUT28), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n222), .A2(new_n235), .A3(new_n277), .A4(new_n244), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n276), .A2(new_n278), .B1(new_n256), .B2(new_n265), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n275), .B1(new_n279), .B2(new_n250), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n256), .A2(new_n265), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n250), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n272), .A2(new_n274), .A3(new_n280), .A4(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(G472), .A2(G902), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT32), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n287), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT32), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n261), .A2(new_n259), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n245), .A2(new_n250), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n188), .B(new_n263), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT71), .B1(new_n270), .B2(KEYINPUT31), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n274), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n285), .A2(new_n280), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n291), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n281), .A2(new_n299), .A3(new_n282), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n235), .B1(new_n244), .B2(new_n222), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n276), .B2(new_n278), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n300), .B(new_n250), .C1(new_n299), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n245), .A2(new_n284), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n259), .B2(new_n261), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n305), .B2(new_n299), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G472), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n298), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n187), .B1(new_n288), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G472), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n303), .B2(new_n306), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n286), .B2(new_n291), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n287), .B1(new_n296), .B2(new_n297), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n290), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT74), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  INV_X1    g131(.A(G902), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(G234), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT22), .B(G137), .Z(new_n320));
  INV_X1    g134(.A(G953), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n321), .A2(G221), .A3(G234), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n320), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G140), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n326), .A2(new_n328), .A3(G146), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n325), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  XNOR2_X1  g144(.A(G125), .B(G140), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n332), .B2(G146), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n230), .A2(G128), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n230), .B2(G128), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n336), .B2(KEYINPUT23), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n236), .A2(G119), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n335), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n337), .A2(G110), .A3(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n339), .A2(new_n334), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT24), .B(G110), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT24), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G110), .ZN(new_n347));
  INV_X1    g161(.A(G110), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT24), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT75), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n342), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n333), .B1(new_n341), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n353));
  OAI21_X1  g167(.A(G110), .B1(new_n337), .B2(new_n340), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n345), .A2(new_n350), .A3(new_n342), .ZN(new_n355));
  INV_X1    g169(.A(new_n330), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n327), .A2(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n325), .A2(G140), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT16), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n356), .A2(new_n359), .A3(G146), .ZN(new_n360));
  AOI21_X1  g174(.A(G146), .B1(new_n356), .B2(new_n359), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n354), .B(new_n355), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n352), .A2(new_n353), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n353), .B1(new_n352), .B2(new_n362), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n324), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n352), .A2(new_n362), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n323), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT25), .B1(new_n368), .B2(new_n318), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n370));
  AOI211_X1 g184(.A(new_n370), .B(G902), .C1(new_n365), .C2(new_n367), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n319), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n365), .A2(new_n367), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n319), .A2(G902), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n310), .A2(new_n316), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(G214), .B1(G237), .B2(G902), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT86), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n218), .A2(G125), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(G125), .B2(new_n242), .ZN(new_n384));
  INV_X1    g198(.A(G224), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G953), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT90), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n384), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G104), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n389), .A2(KEYINPUT3), .A3(G104), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT3), .B1(new_n389), .B2(G104), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G101), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(KEYINPUT79), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n399));
  INV_X1    g213(.A(G104), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n389), .A2(KEYINPUT3), .A3(G104), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n390), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n396), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n394), .A2(G101), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n391), .B(new_n395), .C1(new_n392), .C2(new_n393), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT4), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n406), .B(new_n409), .C1(new_n233), .C2(new_n234), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT5), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n229), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT87), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n223), .A2(KEYINPUT5), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n229), .A2(new_n415), .A3(new_n411), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n413), .A2(new_n414), .A3(G113), .A4(new_n416), .ZN(new_n417));
  OR3_X1    g231(.A1(new_n226), .A2(new_n229), .A3(new_n231), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT80), .B1(new_n389), .B2(G104), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n400), .A3(G107), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n389), .A2(G104), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G101), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n417), .A2(new_n418), .A3(new_n408), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n410), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G122), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n410), .A2(new_n425), .A3(new_n427), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(KEYINPUT6), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n427), .B1(new_n410), .B2(new_n425), .ZN(new_n432));
  XOR2_X1   g246(.A(KEYINPUT88), .B(KEYINPUT6), .Z(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n432), .A2(KEYINPUT89), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT89), .B1(new_n432), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n388), .B(new_n431), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n386), .A2(new_n438), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n384), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n384), .A2(new_n439), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n417), .A2(new_n418), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n424), .A2(new_n408), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n425), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n427), .B(KEYINPUT8), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n440), .A2(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(G902), .B1(new_n447), .B2(new_n430), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n437), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n437), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n382), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT94), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n326), .B2(new_n328), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT91), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT19), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT19), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT92), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n458), .A2(KEYINPUT92), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n331), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n209), .A3(new_n461), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n246), .A2(G143), .A3(G214), .ZN(new_n463));
  AOI21_X1  g277(.A(G143), .B1(new_n246), .B2(G214), .ZN(new_n464));
  OAI21_X1  g278(.A(G131), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G237), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n321), .A3(G214), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n207), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n246), .A2(G143), .A3(G214), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n201), .A3(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n465), .A2(new_n470), .B1(new_n332), .B2(G146), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT18), .A2(G131), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n468), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n472), .B1(new_n468), .B2(new_n469), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n455), .A2(G146), .A3(new_n456), .ZN(new_n476));
  INV_X1    g290(.A(new_n329), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n462), .A2(new_n471), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  XOR2_X1   g293(.A(G113), .B(G122), .Z(new_n480));
  XOR2_X1   g294(.A(KEYINPUT93), .B(G104), .Z(new_n481));
  XOR2_X1   g295(.A(new_n480), .B(new_n481), .Z(new_n482));
  OAI21_X1  g296(.A(new_n453), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n471), .A2(new_n462), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n475), .A2(new_n478), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n482), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(KEYINPUT94), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n356), .A2(new_n359), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n209), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n332), .A2(G146), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT95), .B1(new_n360), .B2(new_n361), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n465), .A2(new_n496), .A3(new_n470), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n496), .B2(new_n465), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n482), .B(new_n485), .C1(new_n495), .C2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n483), .A2(new_n488), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT96), .ZN(new_n501));
  NOR2_X1   g315(.A1(G475), .A2(G902), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n502), .B(KEYINPUT97), .Z(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n483), .A2(new_n488), .A3(new_n499), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT20), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n503), .A2(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n485), .B1(new_n495), .B2(new_n498), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n487), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n499), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n318), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G475), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT9), .B(G234), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n518), .A2(new_n317), .A3(G953), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT14), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n228), .A3(G122), .ZN(new_n521));
  INV_X1    g335(.A(G122), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT14), .B1(new_n522), .B2(G116), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(G116), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT101), .B(new_n521), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT101), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n228), .A2(G122), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n228), .A2(G122), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(KEYINPUT14), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(G107), .A3(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n530), .A2(KEYINPUT102), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(KEYINPUT102), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n236), .A2(G143), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n207), .A2(G128), .ZN(new_n535));
  OAI21_X1  g349(.A(G134), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n207), .A2(G128), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n236), .A2(G143), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n195), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT100), .ZN(new_n541));
  OR3_X1    g355(.A1(new_n528), .A2(new_n524), .A3(G107), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT100), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n536), .A2(new_n543), .A3(new_n539), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n533), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n207), .A2(KEYINPUT13), .A3(G128), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n535), .B2(KEYINPUT99), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(KEYINPUT99), .B2(new_n548), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT13), .B1(new_n207), .B2(G128), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(KEYINPUT98), .ZN(new_n552));
  OAI21_X1  g366(.A(G134), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n539), .ZN(new_n554));
  OAI21_X1  g368(.A(G107), .B1(new_n528), .B2(new_n524), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n542), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n519), .B1(new_n547), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n545), .B1(new_n531), .B2(new_n532), .ZN(new_n559));
  INV_X1    g373(.A(new_n557), .ZN(new_n560));
  INV_X1    g374(.A(new_n519), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n318), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G952), .ZN(new_n567));
  AOI211_X1 g381(.A(G953), .B(new_n567), .C1(G234), .C2(G237), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n318), .B(new_n321), .C1(G234), .C2(G237), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n547), .A2(new_n557), .A3(new_n519), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n561), .B1(new_n559), .B2(new_n560), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n565), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n566), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n452), .A2(new_n517), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G128), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n238), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n408), .A3(new_n424), .ZN(new_n585));
  AND4_X1   g399(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n237), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n581), .A2(G128), .B1(new_n240), .B2(new_n215), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n443), .ZN(new_n589));
  AOI221_X4 g403(.A(KEYINPUT12), .B1(new_n203), .B2(new_n198), .C1(new_n585), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n585), .A2(new_n589), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n204), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT10), .B1(new_n586), .B2(new_n587), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n443), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT4), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n394), .B2(G101), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n408), .A2(new_n598), .B1(new_n397), .B2(new_n405), .ZN(new_n599));
  INV_X1    g413(.A(new_n221), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT70), .B1(new_n211), .B2(new_n217), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n596), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n204), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT82), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n606));
  AND3_X1   g420(.A1(new_n585), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n585), .B2(new_n606), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n603), .B(new_n604), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(G110), .B(G140), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n321), .A2(G227), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n594), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT85), .ZN(new_n615));
  INV_X1    g429(.A(new_n609), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n586), .B1(new_n580), .B2(new_n582), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n606), .B1(new_n617), .B2(new_n443), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT82), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n585), .A2(new_n605), .A3(new_n606), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n604), .B1(new_n621), .B2(new_n603), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n612), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT85), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n594), .A2(new_n609), .A3(new_n624), .A4(new_n613), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n615), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G469), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n318), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n594), .A2(new_n609), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n612), .B(KEYINPUT78), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n607), .A2(new_n608), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n599), .A2(new_n602), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n595), .A2(new_n443), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n204), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n613), .A3(new_n609), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT83), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n632), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n639), .B1(new_n632), .B2(new_n638), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n640), .A2(new_n641), .A3(G902), .ZN(new_n642));
  OAI211_X1 g456(.A(KEYINPUT84), .B(new_n628), .C1(new_n642), .C2(new_n627), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n632), .A2(new_n638), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT83), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n632), .A2(new_n638), .A3(new_n639), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n318), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT84), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n648), .A3(G469), .ZN(new_n649));
  INV_X1    g463(.A(G221), .ZN(new_n650));
  INV_X1    g464(.A(new_n518), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n651), .B2(new_n318), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n579), .A2(new_n643), .A3(new_n649), .A4(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n379), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT103), .B(G101), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G3));
  AND3_X1   g471(.A1(new_n643), .A2(new_n649), .A3(new_n653), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n285), .A2(new_n280), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n292), .A2(new_n293), .A3(new_n273), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n264), .B2(new_n271), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n378), .B(new_n314), .C1(new_n662), .C2(new_n311), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n452), .A2(KEYINPUT104), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n667), .B(new_n382), .C1(new_n450), .C2(new_n451), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n564), .A2(new_n318), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n563), .B2(G478), .ZN(new_n672));
  OAI21_X1  g486(.A(KEYINPUT33), .B1(new_n558), .B2(new_n562), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT33), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n573), .A2(new_n574), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n672), .B1(G478), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n510), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n507), .B2(KEYINPUT20), .ZN(new_n679));
  INV_X1    g493(.A(new_n516), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n669), .A2(new_n572), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n665), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT105), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT34), .B(G104), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G6));
  NAND2_X1  g501(.A1(new_n566), .A2(new_n577), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n501), .A2(new_n506), .ZN(new_n689));
  INV_X1    g503(.A(new_n509), .ZN(new_n690));
  OAI22_X1  g504(.A1(new_n508), .A2(KEYINPUT106), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n507), .B2(KEYINPUT20), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n516), .B(new_n688), .C1(new_n691), .C2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n669), .A3(new_n572), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n665), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT35), .B(G107), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G9));
  AND2_X1   g513(.A1(new_n649), .A2(new_n653), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n363), .A2(new_n364), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n324), .A2(KEYINPUT36), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n703), .A2(new_n375), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n372), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n314), .B(new_n705), .C1(new_n662), .C2(new_n311), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n700), .A2(new_n707), .A3(new_n643), .A4(new_n579), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT37), .B(G110), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G12));
  INV_X1    g524(.A(new_n705), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n666), .B2(new_n668), .ZN(new_n712));
  INV_X1    g526(.A(G900), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n569), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n568), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n694), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT74), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT74), .B1(new_n313), .B2(new_n315), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n722), .A3(new_n658), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G128), .ZN(G30));
  XNOR2_X1  g538(.A(new_n716), .B(KEYINPUT39), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n658), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n726), .A2(KEYINPUT40), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(KEYINPUT40), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n517), .A2(new_n688), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n284), .B1(new_n292), .B2(new_n245), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n318), .B1(new_n304), .B2(new_n301), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n298), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n729), .B1(new_n733), .B2(new_n315), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n450), .A2(new_n451), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT38), .Z(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n737), .A2(new_n381), .A3(new_n705), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n727), .A2(new_n728), .A3(new_n734), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G143), .ZN(G45));
  NAND2_X1  g554(.A1(new_n682), .A2(new_n716), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n722), .A2(new_n658), .A3(new_n712), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G146), .ZN(G48));
  AOI211_X1 g558(.A(new_n571), .B(new_n681), .C1(new_n666), .C2(new_n668), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n626), .A2(new_n318), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(G469), .ZN(new_n747));
  AND4_X1   g561(.A1(new_n378), .A2(new_n747), .A3(new_n628), .A4(new_n653), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n722), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT41), .B(G113), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NAND3_X1  g565(.A1(new_n310), .A2(new_n748), .A3(new_n316), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n696), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n228), .ZN(G18));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n679), .A2(new_n578), .A3(new_n680), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n628), .A2(new_n756), .A3(new_n653), .A4(new_n747), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n722), .A2(new_n755), .A3(new_n712), .A4(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n712), .A2(new_n757), .A3(new_n310), .A4(new_n316), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT107), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G119), .ZN(G21));
  AOI21_X1  g576(.A(new_n729), .B1(new_n666), .B2(new_n668), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n660), .B1(KEYINPUT31), .B2(new_n270), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n302), .A2(new_n250), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n289), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n372), .B1(new_n373), .B2(new_n375), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n286), .A2(new_n318), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(G472), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n628), .A2(new_n747), .A3(new_n653), .A4(new_n572), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n763), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT108), .B(G122), .Z(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G24));
  AOI21_X1  g587(.A(new_n766), .B1(new_n768), .B2(G472), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n682), .A3(new_n705), .A4(new_n716), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n747), .A2(new_n628), .A3(new_n653), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n669), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n325), .ZN(G27));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n437), .A2(new_n448), .ZN(new_n781));
  INV_X1    g595(.A(new_n449), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n437), .A2(new_n448), .A3(new_n449), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n652), .A2(new_n381), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n627), .A2(new_n318), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n638), .A2(KEYINPUT109), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n637), .A2(new_n789), .A3(new_n613), .A4(new_n609), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n788), .A2(new_n790), .B1(new_n629), .B2(new_n631), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n787), .B1(new_n791), .B2(G469), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n786), .B1(new_n792), .B2(new_n628), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n310), .A2(new_n316), .A3(new_n378), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n780), .B1(new_n794), .B2(new_n741), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n378), .B1(new_n288), .B2(new_n309), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n742), .A3(KEYINPUT42), .A4(new_n793), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G131), .ZN(G33));
  NAND4_X1  g614(.A1(new_n722), .A2(new_n378), .A3(new_n718), .A4(new_n793), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NOR2_X1   g616(.A1(new_n679), .A2(new_n680), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n677), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT43), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(KEYINPUT43), .ZN(new_n808));
  MUX2_X1   g622(.A(new_n807), .B(new_n804), .S(new_n808), .Z(new_n809));
  NAND2_X1  g623(.A1(new_n768), .A2(G472), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n711), .B1(new_n810), .B2(new_n314), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT44), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n809), .A2(KEYINPUT44), .A3(new_n811), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n735), .A2(new_n382), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n627), .B1(new_n791), .B2(KEYINPUT45), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n645), .A2(new_n820), .A3(new_n646), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n787), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT46), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n822), .A2(KEYINPUT46), .A3(new_n823), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n628), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n653), .A3(new_n725), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n818), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n814), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  AOI21_X1  g646(.A(KEYINPUT47), .B1(new_n828), .B2(new_n653), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(KEYINPUT47), .A3(new_n653), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n722), .A2(new_n378), .A3(new_n741), .A4(new_n816), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G140), .ZN(G42));
  AND2_X1   g653(.A1(new_n747), .A2(new_n628), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT49), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n733), .A2(new_n315), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n804), .A2(new_n767), .A3(new_n652), .A4(new_n381), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n737), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n372), .A2(new_n704), .A3(new_n653), .A4(new_n716), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n792), .B2(new_n628), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI211_X1 g662(.A(KEYINPUT116), .B(new_n845), .C1(new_n792), .C2(new_n628), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n669), .B(new_n734), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n775), .A2(new_n777), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n723), .A2(new_n743), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n310), .A2(new_n700), .A3(new_n316), .A4(new_n643), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n778), .B1(new_n855), .B2(new_n719), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT52), .A3(new_n743), .A4(new_n850), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT112), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n759), .B(new_n755), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n310), .A2(new_n748), .A3(new_n316), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n695), .A2(new_n669), .A3(new_n572), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n749), .A3(new_n771), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n859), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n793), .A2(new_n682), .A3(new_n716), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(new_n796), .A3(new_n780), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n722), .A2(new_n378), .A3(new_n742), .A4(new_n793), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n867), .B1(new_n868), .B2(new_n780), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n516), .B1(new_n691), .B2(new_n693), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n566), .A2(new_n577), .A3(new_n716), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n870), .A2(new_n816), .A3(new_n711), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n722), .A2(new_n658), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n774), .A2(new_n705), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n742), .A3(new_n793), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n801), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n382), .B(new_n572), .C1(new_n450), .C2(new_n451), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n511), .A2(new_n516), .A3(new_n688), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n803), .A2(KEYINPUT113), .A3(new_n688), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n700), .A3(new_n664), .A4(new_n643), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n708), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n885), .B1(new_n884), .B2(new_n708), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n681), .A2(new_n878), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n700), .A2(new_n664), .A3(new_n643), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n379), .B2(new_n654), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n771), .B1(new_n752), .B2(new_n683), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n753), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(KEYINPUT112), .A3(new_n761), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n865), .A2(new_n877), .A3(new_n892), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n858), .B1(new_n896), .B2(KEYINPUT115), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n799), .A2(new_n801), .A3(new_n873), .A4(new_n875), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n884), .A2(new_n708), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT114), .ZN(new_n900));
  INV_X1    g714(.A(new_n891), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n886), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT115), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n865), .A4(new_n895), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT53), .B1(new_n897), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n854), .A2(new_n857), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT53), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT117), .B1(new_n908), .B2(new_n896), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n865), .A2(new_n895), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n854), .B2(new_n857), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(new_n911), .A3(new_n913), .A4(new_n903), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT54), .B1(new_n906), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n809), .A2(new_n568), .ZN(new_n917));
  INV_X1    g731(.A(new_n776), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n816), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g734(.A(KEYINPUT120), .B(KEYINPUT48), .Z(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n797), .A3(new_n921), .ZN(new_n922));
  AND4_X1   g736(.A1(new_n378), .A2(new_n919), .A3(new_n568), .A4(new_n842), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n567), .B(G953), .C1(new_n923), .C2(new_n682), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n917), .A2(new_n797), .A3(new_n919), .ZN(new_n925));
  NOR2_X1   g739(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n917), .A2(new_n669), .A3(new_n776), .A4(new_n769), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n922), .A2(new_n924), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n736), .A2(new_n918), .A3(new_n382), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n917), .A2(new_n769), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT50), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n517), .A2(new_n677), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n920), .A2(new_n874), .B1(new_n923), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(KEYINPUT51), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n917), .A2(new_n769), .A3(new_n817), .ZN(new_n937));
  INV_X1    g751(.A(new_n835), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n833), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n840), .A2(new_n652), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n929), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n939), .A2(KEYINPUT119), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT119), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n836), .A2(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n943), .A2(new_n945), .A3(new_n940), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n933), .B(new_n935), .C1(new_n946), .C2(new_n937), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT51), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n912), .B1(new_n896), .B2(new_n858), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT54), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n894), .A2(KEYINPUT118), .A3(new_n761), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT118), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n860), .B2(new_n864), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n913), .A2(new_n903), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n950), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n916), .A2(new_n949), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(G952), .A2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n844), .B1(new_n957), .B2(new_n958), .ZN(G75));
  NAND2_X1  g773(.A1(new_n950), .A2(new_n955), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT121), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n961), .A3(G210), .A4(G902), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(new_n388), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT55), .ZN(new_n965));
  XOR2_X1   g779(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n318), .B1(new_n950), .B2(new_n955), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n961), .B1(new_n968), .B2(G210), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n321), .A2(G952), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT56), .B1(new_n968), .B2(G210), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(new_n965), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n970), .A2(new_n974), .ZN(G51));
  XNOR2_X1  g789(.A(new_n787), .B(KEYINPUT57), .ZN(new_n976));
  INV_X1    g790(.A(new_n956), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n951), .B1(new_n950), .B2(new_n955), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n626), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n968), .A2(new_n821), .A3(new_n819), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n971), .B1(new_n980), .B2(new_n981), .ZN(G54));
  INV_X1    g796(.A(KEYINPUT124), .ZN(new_n983));
  INV_X1    g797(.A(new_n689), .ZN(new_n984));
  NAND2_X1  g798(.A1(KEYINPUT58), .A2(G475), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT123), .Z(new_n986));
  NAND3_X1  g800(.A1(new_n968), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n972), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n984), .B1(new_n968), .B2(new_n986), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n983), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n968), .A2(new_n986), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n689), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n992), .A2(KEYINPUT124), .A3(new_n972), .A4(new_n987), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n990), .A2(new_n993), .ZN(G60));
  XNOR2_X1  g808(.A(new_n670), .B(KEYINPUT59), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n676), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n977), .B2(new_n978), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n972), .ZN(new_n998));
  INV_X1    g812(.A(new_n995), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n909), .A2(new_n914), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n896), .A2(KEYINPUT115), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1001), .A2(new_n905), .A3(new_n907), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n912), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n951), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n999), .B1(new_n1004), .B2(new_n977), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n998), .B1(new_n1005), .B2(new_n676), .ZN(G63));
  XNOR2_X1  g820(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n317), .A2(new_n318), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n960), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n971), .B1(new_n1010), .B2(new_n373), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1011), .B(KEYINPUT61), .C1(new_n703), .C2(new_n1010), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT61), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1010), .A2(new_n703), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1009), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n950), .B2(new_n955), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n972), .B1(new_n1016), .B2(new_n368), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1013), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1012), .A2(new_n1018), .ZN(G66));
  AOI21_X1  g833(.A(G953), .B1(new_n910), .B2(new_n892), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT126), .ZN(new_n1021));
  OAI21_X1  g835(.A(G953), .B1(new_n570), .B2(new_n385), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n963), .B1(G898), .B2(new_n321), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(G69));
  AOI22_X1  g839(.A1(new_n814), .A2(new_n830), .B1(new_n836), .B2(new_n837), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n856), .A2(new_n743), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n739), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n881), .A2(new_n681), .A3(new_n882), .ZN(new_n1030));
  OR4_X1    g844(.A1(new_n379), .A2(new_n726), .A3(new_n816), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT62), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1027), .A2(new_n739), .A3(new_n1032), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n1026), .A2(new_n1029), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n321), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n269), .B1(new_n222), .B2(new_n260), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n457), .A2(new_n461), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT127), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1038), .B1(G900), .B2(G953), .ZN(new_n1041));
  INV_X1    g855(.A(new_n763), .ZN(new_n1042));
  OR3_X1    g856(.A1(new_n829), .A2(new_n1042), .A3(new_n796), .ZN(new_n1043));
  AND2_X1   g857(.A1(new_n1027), .A2(new_n801), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1026), .A2(new_n799), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1041), .B1(new_n1045), .B2(G953), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1039), .A2(new_n1040), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n321), .B1(G227), .B2(G900), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1047), .B(new_n1048), .ZN(G72));
  NAND2_X1  g863(.A1(G472), .A2(G902), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1050), .B(KEYINPUT63), .Z(new_n1051));
  NAND2_X1  g865(.A1(new_n910), .A2(new_n892), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1051), .B1(new_n1034), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1053), .A2(new_n730), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1051), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1055), .A2(new_n305), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1054), .A2(new_n972), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1058));
  INV_X1    g872(.A(new_n305), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1059), .A2(new_n1051), .ZN(new_n1060));
  NOR2_X1   g874(.A1(new_n1060), .A2(new_n730), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1057), .B1(new_n1058), .B2(new_n1061), .ZN(G57));
endmodule


