//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272, new_n1273;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n207), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT64), .Z(new_n218));
  OAI22_X1  g0018(.A1(new_n212), .A2(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n223), .B(new_n229), .C1(G58), .C2(G232), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n208), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT1), .Z(new_n232));
  AOI211_X1 g0032(.A(new_n219), .B(new_n232), .C1(new_n213), .C2(new_n212), .ZN(G361));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n222), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G58), .ZN(new_n244));
  INV_X1    g0044(.A(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G97), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G87), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n221), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  OAI211_X1 g0053(.A(G226), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  OAI211_X1 g0054(.A(G232), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n227), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n254), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G238), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT71), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n263), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n259), .A2(new_n262), .B1(new_n266), .B2(G238), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT13), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n273), .A3(new_n269), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(G179), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT73), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n271), .A2(new_n277), .A3(G179), .A4(new_n274), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n273), .B1(new_n272), .B2(new_n269), .ZN(new_n281));
  OAI21_X1  g0081(.A(G169), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT14), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n271), .A2(new_n274), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT74), .B1(new_n279), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n256), .A2(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n289), .A2(G77), .B1(new_n290), .B2(G50), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n207), .B2(G68), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n214), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT11), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n225), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n300), .B(KEYINPUT12), .Z(new_n301));
  AOI21_X1  g0101(.A(KEYINPUT11), .B1(new_n292), .B2(new_n294), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n294), .B1(new_n206), .B2(G20), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n303), .A2(G68), .ZN(new_n304));
  NOR4_X1   g0104(.A1(new_n297), .A2(new_n301), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  XOR2_X1   g0105(.A(new_n305), .B(KEYINPUT75), .Z(new_n306));
  AOI21_X1  g0106(.A(new_n285), .B1(new_n284), .B2(G169), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI211_X1 g0108(.A(KEYINPUT14), .B(new_n308), .C1(new_n271), .C2(new_n274), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT74), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n276), .A2(new_n278), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n288), .A2(new_n306), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n284), .A2(G200), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n271), .A2(G190), .A3(new_n274), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(new_n305), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n317), .A2(KEYINPUT72), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(KEYINPUT72), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n303), .A2(G77), .ZN(new_n321));
  XOR2_X1   g0121(.A(KEYINPUT15), .B(G87), .Z(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n323));
  OR2_X1    g0123(.A1(KEYINPUT8), .A2(G58), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT8), .A2(G58), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n290), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT69), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT69), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n290), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n294), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n321), .B1(G77), .B2(new_n298), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n268), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT3), .B(G33), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G232), .A3(new_n251), .ZN(new_n337));
  OR2_X1    g0137(.A1(KEYINPUT68), .A2(G107), .ZN(new_n338));
  NAND2_X1  g0138(.A1(KEYINPUT68), .A2(G107), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n251), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n337), .B1(new_n336), .B2(new_n340), .C1(new_n344), .C2(new_n226), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n335), .B1(new_n345), .B2(new_n262), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n266), .A2(G244), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n334), .B1(new_n348), .B2(G200), .ZN(new_n349));
  INV_X1    g0149(.A(G190), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n348), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n314), .A2(new_n320), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n203), .A2(KEYINPUT67), .A3(G20), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT67), .ZN(new_n354));
  NOR3_X1   g0154(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(new_n207), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n290), .A2(G150), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n289), .A2(new_n324), .A3(new_n325), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n353), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n294), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n299), .A2(new_n202), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n303), .A2(G50), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n252), .A2(new_n253), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G77), .ZN(new_n365));
  OAI211_X1 g0165(.A(G223), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n366));
  OAI211_X1 g0166(.A(G222), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT66), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n365), .A2(KEYINPUT66), .A3(new_n366), .A4(new_n367), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n262), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n335), .B1(new_n266), .B2(G226), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n363), .B1(new_n374), .B2(G179), .ZN(new_n375));
  AOI21_X1  g0175(.A(G169), .B1(new_n372), .B2(new_n373), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G179), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n346), .A2(new_n378), .A3(new_n347), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n334), .ZN(new_n380));
  AOI21_X1  g0180(.A(G169), .B1(new_n346), .B2(new_n347), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n374), .A2(G200), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT9), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n363), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n372), .A2(G190), .A3(new_n373), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n363), .A2(new_n384), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n383), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT10), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT70), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G200), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n372), .B2(new_n373), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT10), .B1(new_n394), .B2(KEYINPUT70), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n374), .A2(G200), .B1(new_n363), .B2(new_n384), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n385), .A3(new_n386), .A4(new_n396), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n377), .B(new_n382), .C1(new_n392), .C2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(G223), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n336), .A2(KEYINPUT76), .A3(G223), .A4(new_n251), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n336), .A2(G226), .A3(G1698), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n401), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n262), .ZN(new_n406));
  INV_X1    g0206(.A(G232), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n268), .B1(new_n265), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(G200), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  AOI211_X1 g0210(.A(G190), .B(new_n408), .C1(new_n405), .C2(new_n262), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n341), .A2(new_n207), .A3(new_n342), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n341), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n342), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n225), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G58), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n225), .ZN(new_n420));
  OAI21_X1  g0220(.A(G20), .B1(new_n420), .B2(new_n201), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n290), .A2(G159), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n413), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT7), .B1(new_n364), .B2(new_n207), .ZN(new_n425));
  NOR4_X1   g0225(.A1(new_n252), .A2(new_n253), .A3(new_n415), .A4(G20), .ZN(new_n426));
  OAI21_X1  g0226(.A(G68), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n423), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(KEYINPUT16), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n424), .A2(new_n429), .A3(new_n294), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n326), .A2(new_n298), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n303), .B2(new_n326), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT17), .B1(new_n412), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n406), .A2(new_n350), .A3(new_n409), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n408), .B1(new_n405), .B2(new_n262), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(G200), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(new_n430), .A4(new_n432), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n434), .A2(KEYINPUT77), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT77), .B1(new_n434), .B2(new_n439), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n436), .A2(G169), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n436), .A2(new_n378), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n433), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n433), .A2(KEYINPUT18), .A3(new_n443), .A4(new_n444), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n398), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n352), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n343), .B2(G250), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT4), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(G244), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n456), .A2(new_n457), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n336), .A2(G244), .A3(new_n251), .A4(new_n460), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n455), .A2(new_n458), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n262), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n206), .A2(G45), .ZN(new_n469));
  OAI211_X1 g0269(.A(G257), .B(new_n261), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G274), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n308), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n464), .B2(new_n262), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n378), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT78), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n206), .A2(G33), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n333), .A2(new_n481), .A3(new_n298), .A4(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n298), .A2(new_n482), .A3(new_n214), .A4(new_n293), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT78), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n227), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n298), .A2(G97), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n340), .B1(new_n416), .B2(new_n417), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n247), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n207), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n327), .A2(new_n245), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n490), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n487), .B(new_n489), .C1(new_n497), .C2(new_n333), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n478), .A2(new_n480), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n393), .B1(new_n465), .B2(new_n476), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n350), .B(new_n475), .C1(new_n464), .C2(new_n262), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n336), .A2(new_n207), .A3(G68), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n289), .A2(G97), .ZN(new_n504));
  NOR2_X1   g0304(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n505));
  AND2_X1   g0305(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n505), .ZN(new_n508));
  AOI21_X1  g0308(.A(G20), .B1(new_n508), .B2(new_n257), .ZN(new_n509));
  INV_X1    g0309(.A(G87), .ZN(new_n510));
  AND2_X1   g0310(.A1(KEYINPUT68), .A2(G107), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT68), .A2(G107), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n510), .B(new_n227), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n503), .B(new_n507), .C1(new_n509), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n294), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n483), .A2(new_n485), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n322), .ZN(new_n518));
  INV_X1    g0318(.A(new_n322), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n299), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G238), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n522));
  OAI211_X1 g0322(.A(G244), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n262), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n261), .A2(G250), .A3(new_n469), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n308), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n526), .A2(new_n378), .A3(new_n527), .A4(new_n528), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n521), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(G200), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n515), .A2(new_n294), .B1(new_n299), .B2(new_n519), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n517), .A2(G87), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n526), .A2(G190), .A3(new_n527), .A4(new_n528), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n499), .A2(new_n502), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n207), .B1(new_n338), .B2(new_n339), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT23), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n511), .A2(new_n512), .ZN(new_n544));
  OAI211_X1 g0344(.A(KEYINPUT84), .B(KEYINPUT23), .C1(new_n544), .C2(new_n207), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(G20), .B1(KEYINPUT23), .B2(G107), .ZN(new_n547));
  INV_X1    g0347(.A(new_n524), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(G20), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n510), .A2(KEYINPUT83), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n550), .B(new_n207), .C1(new_n252), .C2(new_n253), .ZN(new_n551));
  NAND2_X1  g0351(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT22), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n510), .B1(KEYINPUT83), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n336), .A2(new_n556), .A3(new_n207), .A4(new_n552), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n546), .A2(new_n549), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT85), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT85), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n546), .A2(new_n558), .A3(new_n561), .A4(new_n549), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(KEYINPUT24), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n559), .A2(KEYINPUT85), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n294), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n299), .A2(new_n493), .ZN(new_n567));
  XNOR2_X1  g0367(.A(new_n567), .B(KEYINPUT25), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n517), .B2(G107), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n336), .A2(G250), .A3(new_n251), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G294), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n344), .C2(new_n228), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n262), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n473), .A2(new_n262), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G264), .ZN(new_n576));
  AND4_X1   g0376(.A1(G179), .A2(new_n574), .A3(new_n474), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT86), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT86), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(new_n474), .A3(new_n576), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n579), .B1(new_n580), .B2(G169), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n578), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n570), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n393), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(G190), .B2(new_n580), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n566), .A2(new_n585), .A3(new_n569), .ZN(new_n586));
  OAI211_X1 g0386(.A(G257), .B(new_n251), .C1(new_n252), .C2(new_n253), .ZN(new_n587));
  OAI211_X1 g0387(.A(G264), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n341), .A2(G303), .A3(new_n342), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n262), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n575), .A2(G270), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n474), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n484), .A2(new_n221), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n299), .A2(new_n221), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n293), .A2(new_n214), .B1(G20), .B2(new_n221), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n453), .B(new_n207), .C1(G33), .C2(new_n227), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n596), .A2(KEYINPUT20), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT20), .B1(new_n596), .B2(new_n597), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n594), .B(new_n595), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(G169), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT81), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n593), .A2(new_n600), .A3(KEYINPUT81), .A4(G169), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n593), .A2(KEYINPUT21), .A3(G169), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n593), .A2(new_n378), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n600), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n593), .A2(G200), .ZN(new_n610));
  INV_X1    g0410(.A(new_n600), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n610), .B(new_n611), .C1(new_n350), .C2(new_n593), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n606), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n539), .A2(new_n583), .A3(new_n586), .A4(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n452), .A2(new_n614), .ZN(G372));
  OAI21_X1  g0415(.A(new_n382), .B1(new_n318), .B2(new_n319), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n314), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT88), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n314), .A2(KEYINPUT88), .A3(new_n616), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n442), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n449), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n392), .A2(new_n397), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n377), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n532), .A2(new_n537), .ZN(new_n625));
  XNOR2_X1  g0425(.A(KEYINPUT87), .B(KEYINPUT26), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n499), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n478), .A2(new_n480), .A3(new_n498), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT26), .B1(new_n538), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n630), .A3(new_n532), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n566), .A2(new_n569), .A3(new_n585), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n544), .B1(new_n425), .B2(new_n426), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n492), .A2(new_n494), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G20), .ZN(new_n635));
  INV_X1    g0435(.A(new_n496), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n486), .B(new_n488), .C1(new_n637), .C2(new_n294), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n477), .A2(G200), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n479), .A2(G190), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(new_n629), .A3(new_n532), .A4(new_n537), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n632), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n606), .A2(new_n609), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n583), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n631), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n624), .B1(new_n452), .B2(new_n647), .ZN(G369));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n209), .A2(G20), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n206), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n570), .A2(new_n649), .A3(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n657), .A2(new_n583), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n570), .A2(new_n656), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n632), .B1(new_n659), .B2(KEYINPUT89), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n656), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n583), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n613), .B1(new_n611), .B2(new_n662), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n644), .A2(new_n600), .A3(new_n656), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n645), .A2(new_n656), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n658), .A2(new_n660), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n570), .A2(new_n582), .A3(new_n662), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n669), .A2(new_n674), .ZN(G399));
  NAND2_X1  g0475(.A1(new_n514), .A2(new_n221), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n210), .A2(G41), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n676), .A2(new_n206), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n677), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n217), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT90), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(KEYINPUT90), .B2(new_n678), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT31), .B1(new_n614), .B2(new_n656), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n591), .A2(new_n592), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n529), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n577), .A2(new_n479), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n477), .A2(new_n593), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n378), .A3(new_n580), .A4(new_n529), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n656), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n684), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n690), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT91), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n692), .A2(new_n690), .A3(KEYINPUT91), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n689), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT92), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n538), .A2(new_n629), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(new_n626), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT26), .ZN(new_n707));
  OAI211_X1 g0507(.A(KEYINPUT92), .B(new_n627), .C1(new_n538), .C2(new_n629), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n499), .A2(new_n502), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n625), .A3(new_n586), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n644), .B1(new_n570), .B2(new_n582), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n532), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n662), .C1(new_n709), .C2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n647), .B2(new_n656), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n703), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n683), .B1(new_n719), .B2(G1), .ZN(G364));
  INV_X1    g0520(.A(new_n668), .ZN(new_n721));
  INV_X1    g0521(.A(G45), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n209), .A2(new_n722), .A3(G20), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n677), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n666), .A2(new_n667), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n721), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G13), .A2(G33), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n666), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n214), .B1(G20), .B2(new_n308), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n207), .A2(new_n378), .A3(new_n393), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G190), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n336), .B1(new_n738), .B2(G326), .ZN(new_n739));
  INV_X1    g0539(.A(G303), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n207), .A2(new_n350), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n393), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n739), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n736), .A2(new_n350), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT33), .B(G317), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n207), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n378), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G311), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n741), .A2(new_n750), .ZN(new_n754));
  INV_X1    g0554(.A(G322), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n749), .A2(new_n742), .ZN(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n749), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n753), .B(new_n758), .C1(G329), .C2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n207), .B1(new_n759), .B2(G190), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n748), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT97), .Z(new_n766));
  XNOR2_X1  g0566(.A(new_n754), .B(KEYINPUT94), .ZN(new_n767));
  INV_X1    g0567(.A(new_n751), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n767), .A2(G58), .B1(G77), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT95), .ZN(new_n770));
  INV_X1    g0570(.A(new_n764), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n746), .A2(G68), .B1(G97), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G159), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n760), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT32), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n336), .B1(new_n743), .B2(new_n510), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT96), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n776), .A2(new_n777), .B1(new_n202), .B2(new_n737), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n777), .B2(new_n776), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n770), .A2(new_n772), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n756), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(G107), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n735), .B1(new_n766), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n210), .A2(new_n336), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n218), .A2(G45), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(new_n246), .C2(new_n722), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n210), .A2(new_n364), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G355), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n786), .B(new_n788), .C1(G116), .C2(new_n211), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n733), .A2(new_n735), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n734), .A2(new_n783), .A3(new_n791), .A4(new_n727), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n730), .A2(new_n792), .ZN(G396));
  NAND2_X1  g0593(.A1(new_n382), .A2(KEYINPUT99), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT99), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n380), .B2(new_n381), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n334), .A2(new_n656), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT100), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n797), .A2(new_n351), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n711), .A2(new_n712), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n801), .B(new_n662), .C1(new_n802), .C2(new_n631), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n647), .A2(new_n656), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n382), .A2(new_n656), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n703), .B(new_n807), .Z(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n728), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n746), .A2(G150), .B1(new_n738), .B2(G137), .ZN(new_n810));
  INV_X1    g0610(.A(new_n767), .ZN(new_n811));
  INV_X1    g0611(.A(G143), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n773), .B2(new_n751), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n781), .A2(G68), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n336), .B1(new_n760), .B2(new_n816), .C1(new_n202), .C2(new_n743), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G58), .B2(new_n771), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n737), .A2(new_n740), .B1(new_n227), .B2(new_n764), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n364), .B1(new_n751), .B2(new_n221), .C1(new_n493), .C2(new_n743), .ZN(new_n821));
  INV_X1    g0621(.A(new_n754), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n821), .C1(G294), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n756), .A2(new_n510), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G311), .B2(new_n761), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT98), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n823), .B(new_n826), .C1(new_n757), .C2(new_n745), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n819), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n728), .B1(new_n828), .B2(new_n735), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n735), .A2(new_n731), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(G77), .B2(new_n831), .C1(new_n806), .C2(new_n732), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n809), .A2(new_n832), .ZN(G384));
  NAND3_X1  g0633(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n695), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n434), .A2(new_n439), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT77), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n434), .A2(KEYINPUT77), .A3(new_n439), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(new_n449), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n654), .B1(new_n430), .B2(new_n432), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n841), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n430), .B(new_n432), .C1(new_n410), .C2(new_n411), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n445), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT102), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n433), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n841), .B1(new_n849), .B2(new_n437), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n850), .B(new_n445), .C1(KEYINPUT102), .C2(KEYINPUT37), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n848), .A2(new_n851), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n843), .B1(new_n449), .B2(new_n836), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  AND4_X1   g0658(.A1(new_n311), .A2(new_n312), .A3(new_n283), .A4(new_n286), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n311), .B1(new_n310), .B2(new_n312), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n318), .A2(new_n319), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n306), .B(new_n656), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n306), .A2(new_n656), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n314), .A2(new_n320), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n835), .A2(new_n858), .A3(new_n806), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT40), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n843), .B1(new_n442), .B2(new_n449), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n854), .B1(new_n869), .B2(new_n855), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT40), .B1(new_n870), .B2(new_n853), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n695), .A2(new_n834), .B1(new_n805), .B2(new_n800), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n835), .A2(new_n451), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(G330), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n451), .A2(new_n714), .A3(new_n716), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT103), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT103), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n451), .A2(new_n714), .A3(new_n716), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n624), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n877), .B(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n852), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n842), .B2(new_n852), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT39), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n853), .A2(new_n888), .A3(new_n857), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n314), .A2(new_n656), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n654), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n449), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n797), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n662), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n803), .A2(new_n897), .B1(new_n863), .B2(new_n865), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n885), .B2(new_n886), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n892), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n884), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n206), .B2(new_n650), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n221), .B1(new_n634), .B2(KEYINPUT35), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n215), .C1(KEYINPUT35), .C2(new_n634), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n420), .A2(new_n217), .A3(new_n245), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT101), .Z(new_n908));
  NOR2_X1   g0708(.A1(new_n225), .A2(G50), .ZN(new_n909));
  OAI211_X1 g0709(.A(G1), .B(new_n209), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n903), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT104), .Z(G367));
  OAI21_X1  g0712(.A(new_n710), .B1(new_n638), .B2(new_n662), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n499), .A2(new_n656), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n915), .A2(new_n658), .A3(new_n660), .A4(new_n670), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT42), .Z(new_n917));
  OAI21_X1  g0717(.A(new_n629), .B1(new_n913), .B2(new_n583), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n662), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n662), .B1(new_n534), .B2(new_n535), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n532), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n625), .B2(new_n921), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT105), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT43), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n920), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n920), .B2(new_n927), .ZN(new_n929));
  INV_X1    g0729(.A(new_n669), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n915), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n928), .A2(new_n929), .B1(KEYINPUT106), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(KEYINPUT106), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(KEYINPUT106), .B(new_n931), .C1(new_n928), .C2(new_n929), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n677), .B(KEYINPUT41), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n671), .A2(new_n672), .A3(new_n915), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT107), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n671), .A2(KEYINPUT107), .A3(new_n672), .A4(new_n915), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT44), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n674), .B2(new_n915), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n673), .A2(KEYINPUT44), .A3(new_n914), .A4(new_n913), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n945), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n930), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n671), .B1(new_n663), .B2(new_n670), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(new_n721), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n718), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n945), .A2(new_n949), .A3(new_n669), .A4(new_n950), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n952), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n937), .B1(new_n957), .B2(new_n719), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n934), .B(new_n935), .C1(new_n958), .C2(new_n726), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n924), .A2(new_n733), .ZN(new_n960));
  AOI22_X1  g0760(.A1(G150), .A2(new_n822), .B1(new_n768), .B2(G50), .ZN(new_n961));
  INV_X1    g0761(.A(G137), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n961), .B1(new_n419), .B2(new_n743), .C1(new_n962), .C2(new_n760), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n764), .A2(new_n225), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n738), .A2(G143), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n746), .A2(G159), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n781), .A2(G77), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n336), .A4(new_n967), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n963), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n364), .B1(new_n751), .B2(new_n757), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n743), .A2(new_n221), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n971), .A2(KEYINPUT46), .B1(new_n745), .B2(new_n763), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n970), .B(new_n972), .C1(G317), .C2(new_n761), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n737), .A2(new_n752), .B1(new_n340), .B2(new_n764), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(KEYINPUT46), .B2(new_n971), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n973), .B(new_n975), .C1(new_n740), .C2(new_n811), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n756), .A2(new_n227), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n969), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n728), .B1(new_n979), .B2(new_n735), .ZN(new_n980));
  INV_X1    g0780(.A(new_n784), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n790), .B1(new_n211), .B2(new_n519), .C1(new_n241), .C2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n960), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n959), .A2(new_n983), .ZN(G387));
  INV_X1    g0784(.A(new_n955), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n954), .A2(new_n718), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n677), .A3(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n746), .A2(G311), .B1(new_n738), .B2(G322), .ZN(new_n988));
  INV_X1    g0788(.A(G317), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n988), .B1(new_n740), .B2(new_n751), .C1(new_n811), .C2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT48), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n757), .B2(new_n764), .C1(new_n763), .C2(new_n743), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT49), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n761), .A2(G326), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n993), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n336), .B1(new_n781), .B2(G116), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n336), .B1(new_n227), .B2(new_n756), .C1(new_n737), .C2(new_n773), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n746), .A2(new_n326), .B1(new_n768), .B2(G68), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT110), .Z(new_n1001));
  NOR2_X1   g0801(.A1(new_n519), .A2(new_n764), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n743), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(G77), .ZN(new_n1004));
  INV_X1    g0804(.A(G150), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1004), .B1(new_n202), .B2(new_n754), .C1(new_n1005), .C2(new_n760), .ZN(new_n1006));
  OR4_X1    g0806(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n998), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n735), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n981), .B1(new_n238), .B2(G45), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n676), .B2(new_n787), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n326), .A2(new_n202), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT50), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n225), .B2(new_n245), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n1014), .A2(G45), .A3(new_n676), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1011), .A2(new_n1015), .B1(G107), .B2(new_n211), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n728), .B1(new_n1016), .B2(new_n790), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT109), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n733), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1009), .B(new_n1018), .C1(new_n663), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n726), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n987), .B(new_n1020), .C1(new_n1021), .C2(new_n954), .ZN(G393));
  NAND3_X1  g0822(.A1(new_n952), .A2(new_n726), .A3(new_n956), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n913), .A2(new_n733), .A3(new_n914), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n790), .B1(new_n227), .B2(new_n211), .C1(new_n249), .C2(new_n981), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n737), .A2(new_n1005), .B1(new_n773), .B2(new_n754), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT51), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n764), .A2(new_n245), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n743), .A2(new_n225), .B1(new_n760), .B2(new_n812), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n326), .C2(new_n768), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n364), .B(new_n824), .C1(G50), .C2(new_n746), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n737), .A2(new_n989), .B1(new_n752), .B2(new_n754), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT52), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G283), .A2(new_n1003), .B1(new_n761), .B2(G322), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n336), .B1(new_n771), .B2(G116), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n746), .A2(G303), .B1(G107), .B2(new_n781), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n751), .A2(new_n763), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1032), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n728), .B1(new_n1040), .B2(new_n735), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1024), .A2(new_n1025), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n952), .A2(new_n956), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n985), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT111), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n957), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n955), .B1(new_n952), .B2(new_n956), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n677), .B1(new_n1047), .B2(KEYINPUT111), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1023), .B(new_n1042), .C1(new_n1046), .C2(new_n1048), .ZN(G390));
  AOI21_X1  g0849(.A(new_n891), .B1(new_n853), .B2(new_n857), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n532), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n643), .B2(new_n646), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n656), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1054), .A2(new_n801), .B1(new_n662), .B2(new_n896), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n863), .A2(new_n865), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1050), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n702), .A2(G330), .A3(new_n806), .A4(new_n866), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n803), .A2(new_n897), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n891), .B1(new_n1059), .B2(new_n866), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1057), .B(new_n1058), .C1(new_n890), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT112), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1057), .B1(new_n890), .B2(new_n1060), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n835), .A2(G330), .A3(new_n866), .A4(new_n806), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n887), .B(new_n889), .C1(new_n898), .C2(new_n891), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT112), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1062), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(new_n1021), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n336), .B1(new_n745), .B2(new_n962), .ZN(new_n1072));
  INV_X1    g0872(.A(G128), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n737), .A2(new_n1073), .B1(new_n773), .B2(new_n764), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(G50), .C2(new_n781), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT54), .B(G143), .Z(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(G125), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1077), .A2(new_n751), .B1(new_n1078), .B2(new_n760), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n743), .B2(new_n1005), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1003), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1075), .B(new_n1083), .C1(new_n816), .C2(new_n754), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n815), .B1(new_n221), .B2(new_n754), .C1(new_n763), .C2(new_n760), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G97), .B2(new_n768), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n757), .A2(new_n737), .B1(new_n745), .B2(new_n340), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G87), .B2(new_n1003), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(new_n245), .C2(new_n764), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1084), .B1(new_n1089), .B2(new_n336), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n728), .B1(new_n1090), .B2(new_n735), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n326), .B2(new_n831), .C1(new_n890), .C2(new_n732), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n643), .A2(new_n583), .A3(new_n613), .A4(new_n662), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1093), .A2(KEYINPUT31), .B1(new_n656), .B2(new_n693), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n1095));
  OAI211_X1 g0895(.A(G330), .B(new_n806), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n1056), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1064), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1059), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n835), .A2(G330), .A3(new_n806), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n1056), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n835), .A2(G330), .A3(new_n451), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n882), .A2(new_n624), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1070), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n677), .B1(new_n1070), .B2(new_n1106), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1071), .B(new_n1092), .C1(new_n1108), .C2(new_n1109), .ZN(G378));
  INV_X1    g0910(.A(KEYINPUT115), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n377), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n623), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1111), .B1(new_n623), .B2(new_n1112), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n363), .B(new_n893), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1115), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n363), .A2(new_n893), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1116), .A2(new_n1121), .A3(new_n1119), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n874), .B2(G330), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n667), .B(new_n1125), .C1(new_n868), .C2(new_n873), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n901), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n835), .A2(new_n806), .A3(new_n866), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1130), .A2(new_n871), .B1(new_n867), .B2(KEYINPUT40), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1131), .B2(new_n667), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n874), .A2(G330), .A3(new_n1126), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n900), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1105), .B1(new_n1070), .B2(new_n1106), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1136), .A3(KEYINPUT57), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n677), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT117), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1134), .A2(KEYINPUT116), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1129), .A2(KEYINPUT116), .A3(new_n1134), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n1136), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT57), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT117), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1137), .A2(new_n1145), .A3(new_n677), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1139), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1140), .A2(new_n1141), .A3(new_n726), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n746), .A2(G132), .B1(new_n738), .B2(G125), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G128), .A2(new_n822), .B1(new_n768), .B2(G137), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n771), .A2(G150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1003), .A2(new_n1076), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G33), .B1(new_n761), .B2(G124), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G41), .B1(new_n781), .B2(G159), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n519), .A2(new_n751), .B1(new_n745), .B2(new_n227), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT114), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1004), .B(new_n364), .C1(new_n221), .C2(new_n737), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(G41), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n754), .A2(new_n493), .B1(new_n760), .B2(new_n757), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n756), .A2(new_n419), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1163), .A2(new_n964), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1160), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT58), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n202), .B1(new_n252), .B2(G41), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1166), .A2(new_n1167), .B1(KEYINPUT113), .B2(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1169), .A2(KEYINPUT113), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1158), .A2(new_n1168), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n728), .B1(new_n1172), .B2(new_n735), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(G50), .B2(new_n831), .C1(new_n1125), .C2(new_n732), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1148), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1147), .A2(new_n1175), .ZN(G375));
  OR2_X1    g0976(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n936), .A3(new_n1106), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G283), .A2(new_n822), .B1(new_n1003), .B2(G97), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n740), .B2(new_n760), .C1(new_n340), .C2(new_n751), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n967), .B1(new_n745), .B2(new_n221), .C1(new_n763), .C2(new_n737), .ZN(new_n1181));
  OR3_X1    g0981(.A1(new_n1180), .A2(new_n1002), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n336), .B1(new_n1077), .B2(new_n745), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1164), .B(new_n1183), .C1(G50), .C2(new_n771), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n737), .A2(new_n816), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT118), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n767), .A2(G137), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G159), .A2(new_n1003), .B1(new_n761), .B2(G128), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n751), .A2(new_n1005), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1182), .A2(new_n336), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n728), .B1(new_n1191), .B2(new_n735), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n866), .B2(new_n732), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n225), .B2(new_n830), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1103), .B2(new_n726), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1178), .A2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT119), .Z(G381));
  XOR2_X1   g0997(.A(G375), .B(KEYINPUT120), .Z(new_n1198));
  INV_X1    g0998(.A(G378), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(G381), .A2(G384), .A3(G387), .A4(G390), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(G393), .A2(G396), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(G407));
  NAND3_X1  g1002(.A1(new_n1198), .A2(new_n655), .A3(new_n1199), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(G407), .A2(G213), .A3(new_n1203), .ZN(G409));
  NAND3_X1  g1004(.A1(new_n1147), .A2(G378), .A3(new_n1175), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1135), .A2(new_n726), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1174), .B(new_n1206), .C1(new_n1142), .C2(new_n937), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1199), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G213), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(G343), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1177), .A2(KEYINPUT121), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT60), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT60), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1177), .A2(KEYINPUT121), .A3(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1214), .A2(new_n677), .A3(new_n1106), .A4(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(G384), .A3(new_n1195), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G384), .B1(new_n1217), .B2(new_n1195), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1209), .A2(KEYINPUT122), .A3(new_n1212), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT127), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT62), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT61), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1211), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G2897), .B(new_n1211), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1220), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1211), .A2(G2897), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1218), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1226), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1227), .B2(new_n1221), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1209), .A2(new_n1212), .A3(new_n1221), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT122), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1225), .A2(new_n1236), .A3(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(G393), .A2(G396), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(new_n1201), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1042), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n957), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(KEYINPUT111), .B2(new_n1047), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n679), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1243), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(G387), .A2(new_n1023), .A3(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G390), .A2(new_n983), .A3(new_n959), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(G390), .A2(KEYINPUT125), .A3(new_n983), .A4(new_n959), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1241), .B2(new_n1201), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1242), .B1(new_n1255), .B2(KEYINPUT124), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1255), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G387), .A2(KEYINPUT126), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(G390), .Z(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1240), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT63), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1239), .A2(new_n1262), .A3(new_n1222), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT123), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1237), .A2(new_n1262), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1266), .A2(new_n1260), .A3(new_n1233), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1239), .A2(KEYINPUT123), .A3(new_n1262), .A4(new_n1222), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1261), .A2(new_n1269), .ZN(G405));
  NAND2_X1  g1070(.A1(G375), .A2(new_n1199), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1205), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(new_n1221), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(new_n1260), .ZN(G402));
endmodule


