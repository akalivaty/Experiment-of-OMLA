//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1191, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT64), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT65), .B2(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(G58), .A2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n206), .B(new_n226), .C1(new_n229), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n220), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n211), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(KEYINPUT66), .B(G87), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G222), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G223), .A2(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  OAI211_X1 g0062(.A(G1), .B(G13), .C1(new_n252), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n261), .B(new_n264), .C1(G77), .C2(new_n257), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n267), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n265), .B(new_n269), .C1(new_n215), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G200), .ZN(new_n272));
  INV_X1    g0072(.A(G190), .ZN(new_n273));
  OAI21_X1  g0073(.A(G20), .B1(new_n231), .B2(G50), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT8), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n219), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT68), .B(G58), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(new_n278), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n228), .A2(G33), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n274), .B1(new_n275), .B2(new_n277), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n227), .ZN(new_n285));
  INV_X1    g0085(.A(G13), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n286), .A2(new_n228), .A3(G1), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n283), .A2(new_n285), .B1(new_n214), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n285), .B1(new_n266), .B2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT9), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n272), .B1(new_n273), .B2(new_n271), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n292), .B2(new_n291), .ZN(new_n294));
  XOR2_X1   g0094(.A(new_n294), .B(KEYINPUT10), .Z(new_n295));
  AND2_X1   g0095(.A1(new_n270), .A2(KEYINPUT71), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n270), .A2(KEYINPUT71), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n296), .A2(new_n297), .A3(new_n209), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n220), .A2(G1698), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(G226), .B2(G1698), .ZN(new_n300));
  INV_X1    g0100(.A(G97), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n300), .A2(new_n256), .B1(new_n252), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n264), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n269), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT13), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(new_n298), .B2(new_n304), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(G169), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT14), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n306), .A2(new_n311), .A3(G169), .A4(new_n308), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n307), .A2(KEYINPUT72), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n305), .B(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n310), .B(new_n312), .C1(new_n313), .C2(new_n315), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n277), .A2(new_n214), .B1(new_n282), .B2(new_n216), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n228), .A2(G68), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n285), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n320));
  XNOR2_X1  g0120(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n286), .A2(G1), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n318), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n289), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n321), .B(new_n325), .C1(new_n208), .C2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n323), .A2(new_n328), .A3(new_n324), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n316), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n306), .A2(G200), .A3(new_n308), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n330), .B(new_n333), .C1(new_n315), .C2(new_n273), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n295), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n290), .A2(new_n288), .B1(new_n271), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT69), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(G179), .B2(new_n271), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT70), .ZN(new_n340));
  XOR2_X1   g0140(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n254), .A2(KEYINPUT75), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n345), .A3(new_n252), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n255), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n348));
  OR2_X1    g0148(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n349));
  NAND2_X1  g0149(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n256), .A2(new_n228), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n208), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n231), .B1(new_n280), .B2(new_n208), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(G20), .B1(G159), .B2(new_n276), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n342), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT79), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT76), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(KEYINPUT3), .B2(new_n252), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n252), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n254), .A2(KEYINPUT75), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n359), .B(G33), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n228), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT7), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n349), .A2(new_n350), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n362), .A2(new_n228), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(G68), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT16), .A3(new_n355), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT79), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n342), .C1(new_n353), .C2(new_n356), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n358), .A2(new_n285), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n362), .A2(new_n365), .ZN(new_n375));
  NOR2_X1   g0175(.A1(G223), .A2(G1698), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n215), .B2(G1698), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G87), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n252), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n264), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n269), .B1(new_n270), .B2(new_n220), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT80), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT80), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n269), .B(new_n386), .C1(new_n270), .C2(new_n220), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(new_n273), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G200), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n263), .B1(new_n378), .B2(new_n381), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n384), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n322), .A2(G20), .ZN(new_n394));
  MUX2_X1   g0194(.A(new_n326), .B(new_n394), .S(new_n281), .Z(new_n395));
  NAND3_X1  g0195(.A1(new_n374), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n374), .A2(new_n393), .A3(KEYINPUT17), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n374), .A2(new_n395), .ZN(new_n401));
  AOI21_X1  g0201(.A(G179), .B1(new_n385), .B2(new_n387), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n383), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n336), .B1(new_n391), .B2(new_n384), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT18), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  AOI211_X1 g0208(.A(new_n408), .B(new_n405), .C1(new_n374), .C2(new_n395), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  XOR2_X1   g0210(.A(KEYINPUT8), .B(G58), .Z(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT15), .B(G87), .Z(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n412), .B1(new_n414), .B2(new_n282), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n285), .B1(G77), .B2(new_n289), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n287), .A2(new_n216), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G238), .A2(G1698), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n257), .B(new_n420), .C1(new_n220), .C2(G1698), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(new_n264), .C1(G107), .C2(new_n257), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n263), .A2(G244), .A3(new_n267), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n269), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n336), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n424), .A2(G179), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n419), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR4_X1   g0228(.A1(new_n340), .A2(new_n400), .A3(new_n410), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n424), .A2(G200), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n418), .B(new_n430), .C1(new_n273), .C2(new_n424), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n335), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(G257), .A2(G1698), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n211), .B2(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n362), .B2(new_n365), .ZN(new_n436));
  INV_X1    g0236(.A(G303), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n257), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n264), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n266), .A2(G45), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT82), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT5), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G41), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT82), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n266), .A4(G45), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n442), .A2(new_n446), .A3(G274), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n264), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n442), .A2(new_n447), .A3(new_n446), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(G270), .A3(new_n263), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n439), .A2(G179), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n253), .A2(KEYINPUT76), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n343), .A2(new_n345), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(G33), .ZN(new_n456));
  AOI211_X1 g0256(.A(KEYINPUT76), .B(new_n252), .C1(new_n343), .C2(new_n345), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n434), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n438), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n263), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n452), .B1(new_n264), .B2(new_n448), .ZN(new_n461));
  OAI21_X1  g0261(.A(G169), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT21), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n453), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(G20), .B1(G33), .B2(G283), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n301), .A2(KEYINPUT81), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT81), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n465), .B1(new_n469), .B2(G33), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G20), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n285), .A2(KEYINPUT85), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT85), .B1(new_n285), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT20), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n470), .B(KEYINPUT20), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n285), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(new_n394), .C1(G1), .C2(new_n252), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n471), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n287), .A2(new_n471), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT84), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n464), .A2(new_n488), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n483), .B(new_n486), .C1(new_n478), .C2(new_n479), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n463), .B1(new_n490), .B2(new_n462), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT86), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT86), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n493), .B(new_n463), .C1(new_n490), .C2(new_n462), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n460), .A2(new_n461), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G190), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n496), .B(new_n490), .C1(new_n390), .C2(new_n495), .ZN(new_n497));
  AND4_X1   g0297(.A1(new_n489), .A2(new_n492), .A3(new_n494), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n263), .A2(G250), .A3(new_n441), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n441), .A2(new_n268), .ZN(new_n500));
  XOR2_X1   g0300(.A(new_n500), .B(KEYINPUT83), .Z(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n252), .A2(new_n471), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n362), .A2(new_n365), .B1(new_n217), .B2(G1698), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n209), .A2(new_n258), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n499), .B(new_n502), .C1(new_n506), .C2(new_n263), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n336), .ZN(new_n508));
  INV_X1    g0308(.A(new_n499), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n217), .A2(G1698), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n505), .B(new_n510), .C1(new_n456), .C2(new_n457), .ZN(new_n511));
  INV_X1    g0311(.A(new_n503), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n509), .B1(new_n513), .B2(new_n264), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(new_n313), .A3(new_n502), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n375), .A2(new_n228), .A3(G68), .ZN(new_n516));
  INV_X1    g0316(.A(new_n469), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n379), .A2(new_n210), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT19), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n519), .A2(new_n252), .A3(new_n301), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n517), .A2(new_n518), .B1(G20), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n469), .B2(new_n282), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n285), .ZN(new_n524));
  INV_X1    g0324(.A(new_n482), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n413), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n413), .A2(new_n394), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n508), .A2(new_n515), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n482), .A2(new_n301), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n394), .A2(G97), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n301), .A2(new_n210), .ZN(new_n534));
  NOR2_X1   g0334(.A1(G97), .A2(G107), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT6), .A4(new_n210), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n539));
  AOI21_X1  g0339(.A(G20), .B1(new_n346), .B2(new_n255), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n351), .B1(new_n540), .B2(KEYINPUT7), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(new_n210), .ZN(new_n542));
  AOI211_X1 g0342(.A(new_n531), .B(new_n532), .C1(new_n542), .C2(new_n285), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n253), .A2(new_n255), .A3(G250), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT4), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n217), .B1(new_n362), .B2(new_n365), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n544), .B(new_n547), .C1(new_n548), .C2(KEYINPUT4), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n264), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n451), .A2(new_n263), .ZN(new_n551));
  INV_X1    g0351(.A(G257), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n550), .A2(G190), .A3(new_n450), .A4(new_n554), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n449), .B(new_n553), .C1(new_n549), .C2(new_n264), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n543), .B(new_n555), .C1(new_n556), .C2(new_n390), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n550), .A2(new_n313), .A3(new_n450), .A4(new_n554), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n210), .B1(new_n348), .B2(new_n352), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n536), .A2(new_n537), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n560), .A2(new_n228), .B1(new_n216), .B2(new_n277), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n285), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n531), .ZN(new_n563));
  INV_X1    g0363(.A(new_n532), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n558), .B(new_n565), .C1(new_n556), .C2(G169), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n507), .A2(G200), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n482), .A2(new_n379), .ZN(new_n568));
  AOI211_X1 g0368(.A(new_n527), .B(new_n568), .C1(new_n523), .C2(new_n285), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n514), .A2(G190), .A3(new_n502), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AND4_X1   g0371(.A1(new_n530), .A2(new_n557), .A3(new_n566), .A4(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT88), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n552), .A2(G1698), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(G250), .B2(G1698), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n362), .B2(new_n365), .ZN(new_n576));
  INV_X1    g0376(.A(G294), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n252), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n264), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n451), .A2(G264), .A3(new_n263), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n579), .A2(new_n450), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n573), .B1(new_n581), .B2(new_n336), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(G179), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n450), .A3(new_n580), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(KEYINPUT88), .A3(G169), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n228), .A2(G87), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT22), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n362), .B2(new_n365), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n256), .B2(new_n587), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n210), .A2(G20), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n503), .A2(new_n228), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n591), .A2(KEYINPUT24), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT24), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n590), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n285), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n322), .A2(G20), .A3(new_n210), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(KEYINPUT87), .B2(KEYINPUT25), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(KEYINPUT87), .B2(KEYINPUT25), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(KEYINPUT87), .A3(KEYINPUT25), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n525), .A2(G107), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n603), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n581), .A2(new_n390), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n581), .A2(G190), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n586), .A2(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n498), .A2(new_n572), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n432), .A2(new_n614), .ZN(G372));
  NAND2_X1  g0415(.A1(new_n401), .A2(new_n406), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n408), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n401), .A2(KEYINPUT18), .A3(new_n406), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n334), .A2(new_n428), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n332), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n619), .B1(new_n622), .B2(new_n400), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n340), .B1(new_n623), .B2(new_n295), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n557), .A2(new_n566), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n586), .A2(new_n609), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n492), .A2(new_n489), .A3(new_n494), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n515), .A2(new_n529), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n508), .A2(KEYINPUT89), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n508), .A2(KEYINPUT89), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n611), .A2(new_n612), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(new_n571), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n571), .A2(new_n530), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(new_n566), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n628), .A2(new_n634), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n566), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n632), .A2(new_n635), .A3(new_n571), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n632), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n624), .B1(new_n432), .B2(new_n643), .ZN(G369));
  INV_X1    g0444(.A(new_n322), .ZN(new_n645));
  OR3_X1    g0445(.A1(new_n645), .A2(KEYINPUT27), .A3(G20), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT27), .B1(new_n645), .B2(G20), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n627), .A2(new_n488), .A3(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT90), .ZN(new_n652));
  INV_X1    g0452(.A(new_n650), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n498), .B1(new_n490), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(KEYINPUT90), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  INV_X1    g0457(.A(new_n613), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n609), .A2(new_n650), .ZN(new_n659));
  INV_X1    g0459(.A(new_n626), .ZN(new_n660));
  OAI22_X1  g0460(.A1(new_n658), .A2(new_n659), .B1(new_n660), .B2(new_n653), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n627), .A2(new_n653), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n663), .A2(new_n613), .B1(new_n626), .B2(new_n653), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(G399));
  NOR3_X1   g0465(.A1(new_n517), .A2(G116), .A3(new_n518), .ZN(new_n666));
  INV_X1    g0466(.A(new_n204), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n669), .A3(G1), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n232), .B2(new_n669), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT28), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n637), .A2(new_n635), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n673), .B(new_n632), .C1(new_n628), .C2(new_n634), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n632), .A2(new_n571), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n635), .B1(new_n675), .B2(new_n639), .ZN(new_n676));
  OAI211_X1 g0476(.A(KEYINPUT29), .B(new_n653), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(KEYINPUT93), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT93), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n642), .A2(new_n653), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n678), .B1(new_n682), .B2(new_n677), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n550), .A2(new_n450), .A3(new_n554), .ZN(new_n684));
  INV_X1    g0484(.A(new_n551), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n449), .B1(new_n685), .B2(G270), .ZN(new_n686));
  AOI21_X1  g0486(.A(G179), .B1(new_n686), .B2(new_n439), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n684), .A2(new_n507), .A3(new_n687), .A4(new_n584), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT92), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n553), .B1(new_n549), .B2(new_n264), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n579), .A2(new_n580), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n450), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT92), .A3(new_n507), .A4(new_n687), .ZN(new_n694));
  NOR2_X1   g0494(.A1(KEYINPUT91), .A2(KEYINPUT30), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n514), .A2(new_n495), .A3(G179), .A4(new_n502), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n581), .A2(new_n691), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n507), .A2(new_n453), .ZN(new_n699));
  INV_X1    g0499(.A(new_n695), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n691), .A3(new_n581), .A4(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n690), .A2(new_n694), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n650), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n498), .A2(new_n572), .A3(new_n613), .A4(new_n653), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n698), .A2(new_n701), .A3(new_n688), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n650), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n683), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n672), .B1(new_n712), .B2(G1), .ZN(G364));
  NOR2_X1   g0513(.A1(new_n286), .A2(G20), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G45), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n669), .A2(G1), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n657), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(G330), .B2(new_n656), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT95), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n656), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n228), .B1(KEYINPUT96), .B2(new_n336), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n336), .A2(KEYINPUT96), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n227), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n228), .A2(new_n273), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n313), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n280), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G179), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G190), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n301), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n228), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n729), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n256), .B(new_n736), .C1(G77), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n390), .A2(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G107), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n728), .A2(new_n741), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n379), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n313), .A2(new_n390), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n728), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n746), .B1(G50), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n737), .A2(new_n732), .ZN(new_n751));
  INV_X1    g0551(.A(G159), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n740), .A2(new_n744), .A3(new_n750), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n747), .A2(new_n737), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n731), .B(new_n755), .C1(G68), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G317), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n751), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G329), .ZN(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n762), .B(new_n764), .C1(new_n765), .C2(new_n742), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G326), .B2(new_n749), .ZN(new_n767));
  INV_X1    g0567(.A(new_n745), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G303), .ZN(new_n769));
  INV_X1    g0569(.A(new_n730), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n257), .B1(new_n770), .B2(G322), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n734), .A2(G294), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n767), .A2(new_n769), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(G311), .B2(new_n739), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n727), .B1(new_n758), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n257), .A2(new_n204), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT94), .Z(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G355), .ZN(new_n778));
  INV_X1    g0578(.A(G45), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n250), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n375), .A2(new_n667), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G45), .B2(new_n232), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n778), .B1(G116), .B2(new_n204), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n722), .A2(new_n727), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n724), .A2(new_n775), .A3(new_n785), .A4(new_n717), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n719), .A2(new_n786), .ZN(G396));
  OAI21_X1  g0587(.A(new_n431), .B1(new_n418), .B2(new_n653), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n427), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n428), .A2(new_n653), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n680), .B(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(new_n710), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n716), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n256), .B1(new_n742), .B2(new_n379), .C1(new_n471), .C2(new_n738), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n736), .B1(G311), .B2(new_n763), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n765), .B2(new_n756), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(G303), .C2(new_n749), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n799), .B1(new_n210), .B2(new_n745), .C1(new_n577), .C2(new_n730), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G143), .A2(new_n770), .B1(new_n739), .B2(G159), .ZN(new_n801));
  INV_X1    g0601(.A(G137), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n802), .B2(new_n748), .C1(new_n275), .C2(new_n756), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT34), .Z(new_n804));
  AOI22_X1  g0604(.A1(new_n768), .A2(G50), .B1(new_n763), .B2(G132), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n743), .A2(G68), .ZN(new_n806));
  INV_X1    g0606(.A(new_n280), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n734), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n805), .A2(new_n375), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n800), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n727), .ZN(new_n811));
  INV_X1    g0611(.A(new_n721), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n727), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n216), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n791), .A2(new_n812), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n811), .A2(new_n717), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n795), .A2(new_n816), .ZN(G384));
  INV_X1    g0617(.A(KEYINPUT99), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n653), .B(new_n792), .C1(new_n638), .C2(new_n641), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n790), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT97), .B1(new_n332), .B2(new_n653), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n331), .A2(new_n650), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n332), .A2(new_n334), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n332), .A2(KEYINPUT97), .A3(new_n334), .A4(new_n822), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT98), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n371), .A2(new_n285), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n341), .B1(new_n370), .B2(new_n355), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n395), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n648), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n831), .A2(new_n828), .A3(new_n832), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n410), .B2(new_n400), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n831), .A2(new_n828), .A3(new_n832), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n833), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n831), .A2(new_n406), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n396), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n838), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n401), .A2(new_n832), .ZN(new_n845));
  AND4_X1   g0645(.A1(new_n838), .A2(new_n616), .A3(new_n845), .A4(new_n396), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n837), .B(KEYINPUT38), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n374), .A2(new_n393), .A3(new_n395), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n648), .B1(new_n374), .B2(new_n395), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n838), .A3(new_n616), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n842), .A2(new_n839), .A3(new_n833), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(new_n838), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT38), .B1(new_n854), .B2(new_n837), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n827), .A2(new_n856), .B1(new_n619), .B2(new_n832), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n838), .B1(new_n851), .B2(new_n616), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n846), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n398), .A2(new_n399), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n845), .B1(new_n619), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n858), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n847), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT101), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT39), .B1(new_n848), .B2(new_n855), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT101), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n863), .A2(new_n847), .A3(new_n868), .A4(new_n864), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n332), .A2(new_n650), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n818), .A2(new_n857), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n857), .A2(new_n818), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n624), .B1(new_n683), .B2(new_n432), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n791), .B1(new_n824), .B2(new_n825), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n650), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n705), .A2(new_n706), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n863), .A2(new_n847), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n878), .A2(new_n877), .A3(new_n880), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n856), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n880), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n432), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n886), .B(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(G330), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n876), .B(new_n890), .Z(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n266), .B2(new_n714), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n471), .B1(new_n538), .B2(KEYINPUT35), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n893), .B(new_n229), .C1(KEYINPUT35), .C2(new_n538), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT36), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n233), .B1(new_n280), .B2(new_n208), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n896), .A2(new_n216), .B1(G50), .B2(new_n208), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(G1), .A3(new_n286), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n892), .A2(new_n895), .A3(new_n898), .ZN(G367));
  OR2_X1    g0699(.A1(new_n569), .A2(new_n653), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n675), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT102), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n632), .A2(new_n900), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n675), .A2(KEYINPUT102), .A3(new_n900), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n722), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n256), .B1(new_n749), .B2(G143), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n734), .A2(G68), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n743), .A2(G77), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n770), .A2(G150), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n745), .A2(new_n280), .B1(new_n751), .B2(new_n802), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT106), .Z(new_n915));
  AOI211_X1 g0715(.A(new_n913), .B(new_n915), .C1(G50), .C2(new_n739), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n757), .A2(G159), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n734), .A2(G107), .ZN(new_n918));
  INV_X1    g0718(.A(new_n375), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n919), .B1(new_n759), .B2(new_n751), .C1(new_n469), .C2(new_n742), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n749), .A2(G311), .B1(new_n739), .B2(G283), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n921), .B1(new_n577), .B2(new_n756), .C1(new_n437), .C2(new_n730), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n745), .A2(new_n471), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT46), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT47), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n727), .ZN(new_n928));
  INV_X1    g0728(.A(new_n781), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n784), .B1(new_n204), .B2(new_n414), .C1(new_n241), .C2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n928), .A2(new_n717), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n908), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n625), .B1(new_n543), .B2(new_n653), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n566), .B1(new_n934), .B2(new_n660), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT103), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(KEYINPUT103), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n653), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n663), .A2(new_n625), .A3(new_n613), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT42), .Z(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT104), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n933), .B1(new_n940), .B2(new_n938), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT43), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n907), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n639), .A2(new_n650), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n662), .B1(new_n934), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n946), .B(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n715), .A2(G1), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n934), .A2(new_n947), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n664), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT45), .Z(new_n954));
  NOR2_X1   g0754(.A1(new_n664), .A2(new_n952), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n657), .A2(new_n661), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n663), .A2(new_n613), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n661), .B2(new_n663), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT105), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n657), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n961), .B(KEYINPUT105), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n964), .B1(new_n965), .B2(new_n657), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n712), .B1(new_n959), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n668), .B(KEYINPUT41), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n951), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n932), .B1(new_n950), .B2(new_n969), .ZN(G387));
  OR2_X1    g0770(.A1(new_n711), .A2(new_n966), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n669), .B1(new_n711), .B2(new_n966), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n951), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n966), .A2(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G322), .A2(new_n749), .B1(new_n757), .B2(G311), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n437), .B2(new_n738), .C1(new_n759), .C2(new_n730), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT48), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n765), .B2(new_n735), .C1(new_n577), .C2(new_n745), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT49), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n763), .A2(G326), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n375), .B1(G116), .B2(new_n743), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G159), .A2(new_n749), .B1(new_n743), .B2(G97), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n214), .B2(new_n730), .C1(new_n414), .C2(new_n735), .ZN(new_n985));
  XOR2_X1   g0785(.A(KEYINPUT108), .B(G150), .Z(new_n986));
  OAI22_X1  g0786(.A1(new_n986), .A2(new_n751), .B1(new_n745), .B2(new_n216), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n985), .A2(new_n919), .A3(new_n987), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n208), .B2(new_n738), .C1(new_n281), .C2(new_n756), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n727), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n661), .A2(new_n723), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n238), .A2(G45), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT107), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n411), .A2(new_n214), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT50), .Z(new_n996));
  AOI21_X1  g0796(.A(G45), .B1(G68), .B2(G77), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n666), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n994), .A2(new_n781), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n777), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n999), .B1(G107), .B2(new_n204), .C1(new_n666), .C2(new_n1000), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n716), .B(new_n992), .C1(new_n784), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n975), .B1(new_n991), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n973), .A2(new_n1003), .ZN(G393));
  NOR2_X1   g0804(.A1(new_n742), .A2(new_n379), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n756), .A2(new_n214), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1006), .B(new_n919), .C1(new_n411), .C2(new_n739), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n748), .A2(new_n275), .B1(new_n730), .B2(new_n752), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT51), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n734), .A2(G77), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n768), .A2(G68), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1005), .B(new_n1012), .C1(G143), .C2(new_n763), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT109), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n757), .A2(G303), .B1(new_n763), .B2(G322), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n765), .B2(new_n745), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G317), .A2(new_n749), .B1(new_n770), .B2(G311), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT52), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(G294), .C2(new_n739), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n734), .A2(G116), .ZN(new_n1020));
  AND4_X1   g0820(.A1(new_n256), .A2(new_n1019), .A3(new_n744), .A4(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n727), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n784), .B1(new_n204), .B2(new_n469), .C1(new_n246), .C2(new_n929), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n934), .A2(new_n722), .A3(new_n947), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1022), .A2(new_n717), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n959), .B2(new_n974), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n971), .A2(new_n959), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n669), .B1(new_n971), .B2(new_n959), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(G390));
  OR2_X1    g0830(.A1(new_n870), .A2(new_n721), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n813), .A2(new_n281), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G283), .A2(new_n749), .B1(new_n739), .B2(new_n517), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n210), .B2(new_n756), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1034), .A2(KEYINPUT115), .B1(G77), .B2(new_n734), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n256), .C1(KEYINPUT115), .C2(new_n1034), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n806), .B1(new_n471), .B2(new_n730), .C1(new_n577), .C2(new_n751), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1036), .A2(new_n746), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n986), .A2(new_n745), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT53), .ZN(new_n1040));
  INV_X1    g0840(.A(G128), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1040), .B1(new_n1041), .B2(new_n748), .C1(new_n752), .C2(new_n735), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n756), .A2(new_n802), .ZN(new_n1043));
  INV_X1    g0843(.A(G132), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n730), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(KEYINPUT54), .B(G143), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(G125), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1047), .A2(new_n738), .B1(new_n1048), .B2(new_n751), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n257), .C1(new_n214), .C2(new_n742), .ZN(new_n1051));
  NOR4_X1   g0851(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n727), .B1(new_n1038), .B2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1031), .A2(new_n717), .A3(new_n1032), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n871), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n653), .B(new_n789), .C1(new_n674), .C2(new_n676), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1056), .A2(new_n790), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n826), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n882), .B(new_n1055), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n871), .B1(new_n820), .B2(new_n826), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n870), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n881), .A2(G330), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT110), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n826), .A2(G330), .A3(new_n709), .A4(new_n792), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1059), .B(new_n1066), .C1(new_n870), .C2(new_n1060), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT110), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1061), .A2(new_n1068), .A3(new_n1063), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1054), .B1(new_n1070), .B2(new_n974), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1061), .A2(new_n1068), .A3(new_n1063), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1068), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1067), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT114), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1058), .B1(new_n710), .B2(new_n791), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1062), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n820), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n880), .A2(KEYINPUT111), .A3(G330), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n792), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT111), .B1(new_n880), .B2(G330), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1058), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT112), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT112), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1087), .B(new_n1058), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1086), .A2(new_n1088), .A3(new_n1066), .A4(new_n1057), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT113), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1088), .A2(new_n1066), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT113), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1056), .A2(new_n790), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1085), .B2(KEYINPUT112), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1081), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n888), .A2(G330), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n624), .C1(new_n683), .C2(new_n432), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1077), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1092), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1080), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1098), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(KEYINPUT114), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1076), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n668), .B1(new_n1106), .B2(new_n1070), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1072), .B1(new_n1105), .B2(new_n1107), .ZN(G378));
  NAND2_X1  g0908(.A1(new_n295), .A2(new_n339), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n291), .A2(new_n832), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1109), .B(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(G330), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n886), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1113), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n1116), .C1(new_n883), .C2(new_n885), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n874), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1115), .A2(new_n872), .A3(new_n873), .A4(new_n1117), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n951), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n716), .B1(new_n1116), .B2(new_n812), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n813), .A2(new_n214), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n919), .A2(new_n262), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(G33), .A2(G41), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT116), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n214), .A3(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT117), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n730), .A2(new_n1041), .B1(new_n738), .B2(new_n802), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n735), .A2(new_n275), .B1(new_n1047), .B2(new_n745), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(G125), .C2(new_n749), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1044), .B2(new_n756), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT59), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1126), .B1(G159), .B2(new_n743), .ZN(new_n1134));
  INV_X1    g0934(.A(G124), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n751), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1128), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n910), .B1(new_n301), .B2(new_n756), .C1(new_n280), .C2(new_n742), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n414), .A2(new_n738), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n216), .A2(new_n745), .B1(new_n730), .B2(new_n210), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1124), .A2(new_n1138), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1141), .B1(new_n471), .B2(new_n748), .C1(new_n765), .C2(new_n751), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n727), .B1(new_n1137), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT119), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1122), .A2(new_n1123), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1121), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1103), .B1(new_n1070), .B2(new_n1096), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1152), .A3(KEYINPUT57), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n668), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT57), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1149), .B1(new_n1154), .B2(new_n1155), .ZN(G375));
  OAI211_X1 g0956(.A(new_n1080), .B(new_n1098), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n968), .B(KEYINPUT120), .Z(new_n1158));
  NOR3_X1   g0958(.A1(new_n1096), .A2(new_n1077), .A3(new_n1098), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT114), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1157), .B(new_n1158), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G137), .A2(new_n770), .B1(new_n743), .B2(new_n807), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n1041), .B2(new_n751), .C1(new_n275), .C2(new_n738), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G50), .B2(new_n734), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n919), .B1(new_n757), .B2(new_n1046), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n1044), .C2(new_n748), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G159), .B2(new_n768), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n735), .A2(new_n414), .B1(new_n748), .B2(new_n577), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n911), .B1(new_n210), .B2(new_n738), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(G303), .C2(new_n763), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n257), .B1(new_n768), .B2(G97), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n765), .C2(new_n730), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G116), .B2(new_n757), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n727), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n717), .B(new_n1174), .C1(new_n826), .C2(new_n721), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n208), .B2(new_n813), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1102), .B2(new_n951), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1161), .A2(new_n1177), .ZN(G381));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1098), .B1(new_n1076), .B2(new_n1102), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1180), .B2(new_n1151), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n668), .A3(new_n1153), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1070), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n669), .B1(new_n1184), .B2(new_n1076), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1071), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1182), .A2(new_n1186), .A3(new_n1149), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n973), .A2(new_n786), .A3(new_n719), .A4(new_n1003), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(G387), .A2(G390), .A3(G384), .A4(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n1177), .A3(new_n1161), .A4(new_n1189), .ZN(G407));
  NAND3_X1  g0990(.A1(new_n1182), .A2(new_n1186), .A3(new_n1149), .ZN(new_n1191));
  OAI211_X1 g0991(.A(G407), .B(G213), .C1(G343), .C2(new_n1191), .ZN(G409));
  INV_X1    g0992(.A(KEYINPUT121), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1194), .A2(new_n1102), .A3(new_n1103), .A4(new_n1067), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1151), .B1(new_n1195), .B2(new_n1103), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1148), .B1(new_n1196), .B2(new_n1158), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1193), .B1(new_n1197), .B2(G378), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G378), .B(new_n1149), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1150), .A2(new_n1152), .A3(new_n1158), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1149), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1186), .A2(KEYINPUT121), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1198), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT60), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1157), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1096), .A2(KEYINPUT60), .A3(new_n1098), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1106), .A4(new_n668), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1177), .ZN(new_n1208));
  INV_X1    g1008(.A(G384), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1207), .A2(G384), .A3(new_n1177), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n649), .A2(G213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1203), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT62), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1203), .A2(new_n1214), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n649), .A2(KEYINPUT122), .A3(G213), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1210), .A2(new_n1211), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n649), .A2(G213), .A3(G2897), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1220), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1210), .A2(new_n1211), .A3(new_n1222), .A4(new_n1218), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1217), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT61), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT62), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1203), .A2(new_n1227), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1216), .A2(new_n1225), .A3(new_n1226), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G387), .A2(new_n1029), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1188), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1230), .A2(new_n1232), .A3(KEYINPUT123), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(G387), .A2(new_n1029), .B1(new_n1232), .B2(KEYINPUT123), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n969), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1235), .A2(new_n949), .B1(new_n908), .B2(new_n931), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1236), .A2(G390), .A3(new_n1188), .A4(new_n1231), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1233), .B1(new_n1238), .B2(new_n1230), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1229), .A2(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1203), .A2(new_n1214), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT63), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1215), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1203), .A2(new_n1214), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1244), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1213), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT125), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1215), .B2(new_n1242), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT124), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1239), .B2(KEYINPUT61), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1234), .A2(new_n1237), .B1(G387), .B2(new_n1029), .ZN(new_n1250));
  OAI211_X1 g1050(.A(KEYINPUT124), .B(new_n1226), .C1(new_n1250), .C2(new_n1233), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1243), .A2(new_n1245), .A3(new_n1247), .A4(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1240), .A2(new_n1253), .ZN(G405));
  AOI21_X1  g1054(.A(new_n1186), .B1(new_n1182), .B2(new_n1149), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1212), .B1(new_n1187), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT127), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1212), .B(KEYINPUT127), .C1(new_n1187), .C2(new_n1255), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G375), .A2(G378), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n1191), .A3(new_n1213), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1261), .A2(new_n1213), .A3(KEYINPUT126), .A4(new_n1191), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1260), .A2(new_n1239), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1239), .B1(new_n1260), .B2(new_n1266), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(G402));
endmodule


