//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n203), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(G20), .A3(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n202), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n212), .B1(new_n206), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT64), .ZN(new_n247));
  INV_X1    g0047(.A(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G33), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT65), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n247), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n247), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(G50), .A3(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n259), .B(new_n267), .C1(G50), .C2(new_n262), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n213), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G226), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n279), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G223), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n284), .B1(new_n221), .B2(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  AOI211_X1 g0087(.A(new_n278), .B(new_n281), .C1(new_n287), .C2(new_n279), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n268), .A2(new_n269), .B1(new_n288), .B2(G190), .ZN(new_n289));
  INV_X1    g0089(.A(G200), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n289), .B(new_n291), .C1(new_n269), .C2(new_n268), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n268), .C1(G169), .C2(new_n288), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G107), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n282), .A2(new_n283), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n302), .B1(new_n303), .B2(new_n230), .C1(new_n216), .C2(new_n285), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n279), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n279), .A2(new_n276), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n278), .B1(G244), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G179), .B2(new_n308), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT15), .B(G87), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT66), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT67), .A3(new_n250), .ZN(new_n315));
  INV_X1    g0115(.A(new_n252), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT67), .B1(new_n314), .B2(new_n250), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n247), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n221), .B1(new_n265), .B2(G20), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n264), .A2(new_n321), .B1(new_n221), .B2(new_n263), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n312), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n323), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n308), .A2(G200), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n325), .B(new_n326), .C1(new_n327), .C2(new_n308), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n297), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT68), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n332), .B1(new_n303), .B2(new_n280), .C1(new_n230), .C2(new_n285), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n279), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n278), .B1(G238), .B2(new_n306), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n335), .B1(new_n334), .B2(new_n336), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n309), .A2(KEYINPUT70), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT14), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n339), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n337), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(new_n341), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n343), .B(new_n347), .C1(new_n294), .C2(new_n345), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n264), .A2(G68), .A3(new_n266), .ZN(new_n349));
  XOR2_X1   g0149(.A(new_n349), .B(KEYINPUT69), .Z(new_n350));
  INV_X1    g0150(.A(KEYINPUT64), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n246), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n250), .A2(G77), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n355), .A2(KEYINPUT11), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n263), .A2(new_n202), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT12), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(KEYINPUT11), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n350), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n348), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n340), .A2(G190), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n345), .A2(G200), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n330), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n352), .A2(new_n262), .A3(new_n316), .A4(new_n266), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n263), .A2(new_n252), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT75), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n372), .A3(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT73), .B1(new_n201), .B2(new_n202), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(G58), .A3(G68), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n377), .A3(new_n203), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(G20), .B1(G159), .B2(new_n256), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n245), .A2(KEYINPUT71), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT71), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G33), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT3), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT72), .B1(new_n245), .B2(KEYINPUT3), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT72), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n381), .A2(new_n383), .A3(new_n389), .A4(KEYINPUT3), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n387), .A2(new_n388), .A3(new_n248), .A4(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n391), .A2(G68), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n387), .A2(new_n248), .A3(new_n390), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT7), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n380), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n352), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT74), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n388), .A2(G20), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT3), .B1(new_n381), .B2(new_n383), .ZN(new_n399));
  INV_X1    g0199(.A(new_n300), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n388), .B1(new_n282), .B2(G20), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n202), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n380), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n397), .B1(new_n404), .B2(KEYINPUT16), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT74), .B(new_n406), .C1(new_n403), .C2(new_n380), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n374), .B1(new_n396), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n306), .A2(G232), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n277), .B2(new_n273), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n387), .A2(new_n390), .ZN(new_n412));
  NOR2_X1   g0212(.A1(G223), .A2(G1698), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n280), .B2(G1698), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n411), .B1(new_n417), .B2(new_n279), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G179), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n412), .A2(new_n414), .B1(G33), .B2(G87), .ZN(new_n420));
  INV_X1    g0220(.A(new_n279), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(G169), .B1(new_n422), .B2(new_n411), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT18), .B1(new_n409), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n394), .A2(G68), .A3(new_n391), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(KEYINPUT16), .A3(new_n379), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT71), .B(G33), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n300), .B1(new_n429), .B2(KEYINPUT3), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n301), .A2(new_n248), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n430), .A2(new_n398), .B1(new_n431), .B2(new_n388), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n379), .B1(new_n432), .B2(new_n202), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT74), .B1(new_n433), .B2(new_n406), .ZN(new_n434));
  INV_X1    g0234(.A(new_n407), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n247), .B(new_n428), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n371), .A2(new_n373), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(new_n424), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n426), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n411), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(new_n327), .C1(new_n421), .C2(new_n420), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n418), .B2(G200), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n434), .A2(new_n435), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n428), .A2(new_n247), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n437), .B(new_n444), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT17), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n437), .A4(new_n444), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n441), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n367), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n275), .A2(G1), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(new_n218), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n421), .A2(new_n456), .B1(new_n272), .B2(new_n455), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n216), .A2(G1698), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n385), .B1(new_n429), .B2(KEYINPUT3), .ZN(new_n460));
  AND4_X1   g0260(.A1(new_n389), .A2(new_n381), .A3(new_n383), .A4(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT81), .B(G116), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n429), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G244), .B(G1698), .C1(new_n460), .C2(new_n461), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n222), .B1(new_n387), .B2(new_n390), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT80), .B1(new_n472), .B2(G1698), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n468), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n458), .B1(new_n474), .B2(new_n279), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT19), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n250), .A2(G97), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n248), .B1(new_n332), .B2(new_n476), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n217), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n476), .A2(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n412), .A2(new_n248), .A3(G68), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g0283(.A(new_n313), .B(KEYINPUT66), .Z(new_n484));
  AOI22_X1  g0284(.A1(new_n483), .A2(new_n247), .B1(new_n263), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n265), .A2(G33), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n264), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n314), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n475), .A2(new_n294), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n469), .A2(new_n470), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n472), .A2(KEYINPUT80), .A3(G1698), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n467), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n457), .B1(new_n493), .B2(new_n421), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n309), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n475), .A2(G190), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(G200), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n488), .A2(G87), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n497), .A2(new_n485), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT79), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT4), .B1(new_n472), .B2(new_n283), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n282), .A2(G250), .A3(G1698), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT4), .A2(G244), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n504), .B(new_n505), .C1(new_n303), .C2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n279), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G41), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n455), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n274), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT77), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n509), .B2(G41), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n511), .A2(new_n272), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n514), .A2(new_n512), .A3(new_n455), .A4(new_n510), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n421), .A3(G257), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT78), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n517), .A2(new_n421), .A3(KEYINPUT78), .A4(G257), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n502), .B1(new_n508), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G244), .B(new_n283), .C1(new_n460), .C2(new_n461), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n507), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n502), .B(new_n522), .C1(new_n526), .C2(new_n421), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G190), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT76), .B1(new_n432), .B2(new_n223), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n223), .A2(KEYINPUT6), .A3(G97), .ZN(new_n532));
  INV_X1    g0332(.A(G97), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n223), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n479), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n532), .B1(new_n535), .B2(KEYINPUT6), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n432), .A2(KEYINPUT76), .A3(new_n223), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n247), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n262), .A2(G97), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n488), .B2(G97), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n522), .B1(new_n526), .B2(new_n421), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(G200), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n508), .A2(new_n294), .A3(new_n522), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(KEYINPUT79), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n527), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n309), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n530), .A2(new_n545), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n465), .A2(new_n464), .A3(new_n248), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n248), .A2(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT23), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n217), .A2(G20), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT22), .B1(new_n282), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n412), .A2(KEYINPUT22), .A3(new_n248), .A4(G87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT24), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT24), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n562), .A3(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n247), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n223), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT82), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT25), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n262), .B2(G107), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n569), .B(KEYINPUT83), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n223), .B2(new_n487), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n517), .A2(new_n421), .A3(G264), .ZN(new_n574));
  MUX2_X1   g0374(.A(G250), .B(G257), .S(G1698), .Z(new_n575));
  AOI22_X1  g0375(.A1(new_n412), .A2(new_n575), .B1(G294), .B2(new_n465), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(new_n576), .B2(new_n421), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n516), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n575), .B1(new_n460), .B2(new_n461), .ZN(new_n580));
  INV_X1    g0380(.A(G294), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n429), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n279), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n515), .A3(new_n574), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n565), .A2(new_n573), .A3(new_n579), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(new_n294), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n309), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n352), .B1(new_n561), .B2(new_n563), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(new_n572), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n505), .B(new_n248), .C1(G33), .C2(new_n533), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n246), .B(new_n592), .C1(new_n464), .C2(new_n248), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT20), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n264), .A2(G116), .A3(new_n486), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n463), .A2(G20), .A3(new_n261), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n517), .A2(new_n421), .A3(G270), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n515), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(G257), .A2(G1698), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n224), .B2(G1698), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n412), .A2(new_n603), .B1(G303), .B2(new_n301), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n601), .B1(new_n604), .B2(new_n421), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n598), .A2(G169), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n598), .A2(KEYINPUT21), .A3(G169), .A4(new_n605), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n603), .B1(new_n460), .B2(new_n461), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n301), .A2(G303), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n600), .B1(new_n612), .B2(new_n279), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n598), .A2(G179), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n598), .B1(G200), .B2(new_n605), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(G190), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n551), .A2(new_n591), .A3(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n454), .A2(new_n501), .A3(new_n620), .ZN(G372));
  XNOR2_X1  g0421(.A(new_n441), .B(KEYINPUT85), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n366), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n312), .A2(new_n625), .A3(new_n323), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT86), .B1(new_n311), .B2(new_n325), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI211_X1 g0428(.A(new_n451), .B(new_n624), .C1(new_n363), .C2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n293), .B1(new_n623), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n296), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n474), .A2(KEYINPUT84), .A3(new_n279), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT84), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n493), .B2(new_n421), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n458), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n490), .B1(new_n636), .B2(G169), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n496), .A2(new_n500), .A3(new_n547), .A4(new_n550), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n547), .A2(new_n550), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n485), .A2(new_n499), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(G190), .B2(new_n475), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n636), .B2(new_n290), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n642), .A2(new_n645), .A3(new_n646), .A4(new_n637), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n551), .A2(new_n586), .A3(new_n637), .A4(new_n645), .ZN(new_n648));
  INV_X1    g0448(.A(new_n590), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n615), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n640), .B(new_n647), .C1(new_n648), .C2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n632), .B1(new_n454), .B2(new_n652), .ZN(G369));
  NAND2_X1  g0453(.A1(new_n261), .A2(new_n248), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT87), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT87), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n598), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n619), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n665), .B2(new_n663), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n662), .B1(new_n589), .B2(new_n572), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n591), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n662), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n590), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n615), .A2(new_n671), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n591), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n590), .B2(new_n662), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n673), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n207), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n480), .A2(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n210), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n651), .A2(new_n687), .A3(new_n671), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT89), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n649), .B2(new_n615), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n665), .A2(KEYINPUT89), .A3(new_n590), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n645), .A2(new_n637), .ZN(new_n693));
  INV_X1    g0493(.A(new_n543), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n544), .A2(G200), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n694), .B(new_n695), .C1(new_n327), .C2(new_n549), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n641), .A2(new_n696), .A3(new_n586), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n638), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n642), .A2(new_n645), .A3(KEYINPUT26), .A4(new_n637), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n639), .A2(new_n646), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n662), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n688), .B1(new_n703), .B2(new_n687), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT31), .B1(new_n620), .B2(new_n501), .ZN(new_n706));
  AND4_X1   g0506(.A1(new_n294), .A2(new_n584), .A3(new_n544), .A4(new_n605), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n633), .A2(new_n635), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n458), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n613), .A2(new_n583), .A3(G179), .A4(new_n574), .ZN(new_n710));
  NOR4_X1   g0510(.A1(new_n549), .A2(KEYINPUT30), .A3(new_n494), .A4(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n494), .A2(new_n710), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n529), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n709), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT88), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT88), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n709), .C1(new_n711), .C2(new_n714), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT31), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n706), .B1(new_n719), .B2(new_n671), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n662), .A2(KEYINPUT31), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n715), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n705), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n686), .B1(new_n726), .B2(G1), .ZN(G364));
  NOR2_X1   g0527(.A1(new_n260), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n265), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n681), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n668), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G330), .B2(new_n666), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n212), .B1(G20), .B2(new_n309), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n327), .A2(G200), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n248), .B1(new_n736), .B2(new_n294), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n533), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n248), .A2(new_n294), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT92), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n736), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n201), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n248), .A2(G179), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G190), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G159), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n738), .B(new_n743), .C1(KEYINPUT32), .C2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n744), .A2(G190), .A3(G200), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n282), .B1(new_n750), .B2(new_n217), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT94), .Z(new_n752));
  NAND2_X1  g0552(.A1(new_n741), .A2(new_n745), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G77), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n744), .A2(new_n327), .A3(G200), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(new_n223), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n739), .A2(new_n327), .A3(G200), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n757), .B1(new_n202), .B2(new_n758), .C1(new_n748), .C2(KEYINPUT32), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n739), .A2(G190), .A3(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT93), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n760), .A2(KEYINPUT93), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n759), .B1(G50), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n749), .A2(new_n752), .A3(new_n755), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n282), .B1(new_n747), .B2(G329), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n769), .B2(new_n756), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n754), .B2(G311), .ZN(new_n771));
  INV_X1    g0571(.A(new_n742), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G322), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n765), .A2(G326), .ZN(new_n774));
  INV_X1    g0574(.A(G303), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n737), .A2(new_n581), .B1(new_n750), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n758), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n771), .A2(new_n773), .A3(new_n774), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n735), .B1(new_n767), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n734), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n240), .A2(new_n275), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT91), .Z(new_n788));
  NOR2_X1   g0588(.A1(new_n412), .A2(new_n680), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n789), .C1(G45), .C2(new_n210), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n680), .A2(new_n301), .ZN(new_n791));
  INV_X1    g0591(.A(G116), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n791), .A2(G355), .B1(new_n792), .B2(new_n680), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n786), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n731), .B(KEYINPUT90), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n781), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n784), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n666), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n733), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n662), .A2(new_n323), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n626), .A2(new_n627), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT98), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n324), .A2(new_n328), .A3(new_n802), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n807), .A2(new_n805), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n806), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n652), .B2(new_n662), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n651), .A2(new_n671), .A3(new_n809), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n731), .B1(new_n814), .B2(new_n724), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n814), .A2(new_n724), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n764), .A2(new_n818), .B1(new_n255), .B2(new_n758), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT96), .ZN(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  INV_X1    g0621(.A(G159), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n742), .C1(new_n822), .C2(new_n753), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT97), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n412), .ZN(new_n827));
  INV_X1    g0627(.A(new_n737), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(G58), .B1(new_n747), .B2(G132), .ZN(new_n829));
  INV_X1    g0629(.A(G50), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n750), .C1(new_n202), .C2(new_n756), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n826), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n825), .B2(new_n824), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n738), .B1(new_n772), .B2(G294), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT95), .Z(new_n835));
  OAI22_X1  g0635(.A1(new_n758), .A2(new_n769), .B1(new_n750), .B2(new_n223), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n282), .B1(new_n747), .B2(G311), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n217), .B2(new_n756), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n836), .B(new_n838), .C1(new_n754), .C2(new_n464), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n835), .B(new_n839), .C1(new_n775), .C2(new_n764), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n735), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n734), .A2(new_n782), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n795), .B1(G77), .B2(new_n843), .C1(new_n809), .C2(new_n783), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n816), .A2(new_n817), .B1(new_n841), .B2(new_n844), .ZN(G384));
  NOR2_X1   g0645(.A1(new_n728), .A2(new_n265), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n419), .A2(new_n423), .A3(new_n660), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT102), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n427), .B2(new_n379), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n848), .B1(new_n849), .B2(new_n352), .ZN(new_n850));
  OAI211_X1 g0650(.A(KEYINPUT102), .B(new_n247), .C1(new_n395), .C2(KEYINPUT16), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n851), .A3(new_n428), .ZN(new_n852));
  INV_X1    g0652(.A(new_n370), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n447), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n438), .A2(new_n424), .ZN(new_n857));
  INV_X1    g0657(.A(new_n660), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n438), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n857), .A2(new_n859), .A3(new_n860), .A4(new_n447), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n660), .B1(new_n852), .B2(new_n853), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n441), .B2(new_n451), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n862), .A2(new_n864), .A3(KEYINPUT38), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT38), .B1(new_n862), .B2(new_n864), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT103), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n862), .A2(new_n864), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT103), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n862), .A2(new_n864), .A3(KEYINPUT38), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n362), .A2(new_n662), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n363), .A2(new_n366), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n362), .B(new_n662), .C1(new_n624), .C2(new_n348), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n809), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n716), .A2(new_n721), .A3(new_n718), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n720), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT105), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(KEYINPUT105), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n451), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n859), .B1(new_n622), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n857), .A2(new_n447), .ZN(new_n892));
  INV_X1    g0692(.A(new_n859), .ZN(new_n893));
  OR4_X1    g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(KEYINPUT37), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n892), .B2(new_n893), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n891), .A3(new_n861), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n869), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n883), .B1(new_n898), .B2(new_n872), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n881), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n888), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n720), .A2(new_n880), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n453), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n901), .B2(new_n903), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT39), .B1(new_n898), .B2(new_n872), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n870), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n363), .A2(new_n662), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n324), .A2(new_n662), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n812), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n878), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n918), .A2(new_n874), .B1(new_n623), .B2(new_n660), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n631), .B1(new_n704), .B2(new_n453), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n920), .B(new_n921), .Z(new_n922));
  AOI21_X1  g0722(.A(new_n846), .B1(new_n907), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n922), .B2(new_n907), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n212), .A2(new_n248), .A3(new_n792), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT99), .Z(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT36), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(KEYINPUT36), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n211), .A2(G77), .A3(new_n377), .A4(new_n375), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(KEYINPUT100), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(KEYINPUT100), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(G50), .C2(new_n202), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(G1), .A3(new_n260), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT101), .Z(new_n938));
  NAND4_X1  g0738(.A1(new_n924), .A2(new_n931), .A3(new_n932), .A4(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT106), .ZN(G367));
  INV_X1    g0740(.A(new_n789), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n236), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n785), .B1(new_n484), .B2(new_n207), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n795), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(KEYINPUT46), .A2(G116), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n533), .A2(new_n756), .B1(new_n750), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(G107), .B2(new_n828), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n777), .A2(G294), .B1(new_n747), .B2(G317), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n827), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT46), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n750), .B2(new_n463), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n951), .B1(new_n753), .B2(new_n769), .C1(new_n775), .C2(new_n742), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n949), .B(new_n952), .C1(G311), .C2(new_n765), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n772), .A2(G150), .B1(G68), .B2(new_n828), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n821), .B2(new_n764), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT109), .Z(new_n956));
  OAI221_X1 g0756(.A(new_n282), .B1(new_n746), .B2(new_n818), .C1(new_n201), .C2(new_n750), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n758), .A2(new_n822), .B1(new_n756), .B2(new_n221), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n957), .B(new_n958), .C1(new_n754), .C2(G50), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n953), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT47), .Z(new_n961));
  AOI21_X1  g0761(.A(new_n944), .B1(new_n961), .B2(new_n734), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n643), .A2(new_n662), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n645), .A2(new_n637), .A3(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n637), .A2(new_n963), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n962), .B1(new_n798), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n551), .B1(new_n694), .B2(new_n671), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n642), .A2(new_n662), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n677), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT108), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT44), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n970), .A2(new_n677), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT45), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(new_n673), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n676), .B1(new_n672), .B2(new_n675), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n667), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n725), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n726), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n681), .B(KEYINPUT41), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n730), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n968), .A2(new_n969), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n987), .A2(new_n591), .A3(new_n675), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT107), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n696), .A2(new_n649), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n662), .B1(new_n991), .B2(new_n641), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n988), .B2(KEYINPUT42), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n990), .A2(new_n993), .B1(KEYINPUT43), .B2(new_n966), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n673), .A2(new_n970), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n967), .B1(new_n986), .B2(new_n998), .ZN(G387));
  INV_X1    g0799(.A(new_n791), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n1000), .A2(new_n683), .B1(G107), .B2(new_n207), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n233), .A2(new_n275), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT110), .Z(new_n1003));
  OAI211_X1 g0803(.A(new_n683), .B(new_n275), .C1(new_n202), .C2(new_n221), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT111), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(KEYINPUT111), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n252), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT50), .B1(new_n252), .B2(G50), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1009), .A2(new_n789), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1001), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n795), .B1(new_n1011), .B2(new_n786), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n756), .A2(new_n533), .B1(new_n746), .B2(new_n255), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n758), .A2(new_n252), .B1(new_n750), .B2(new_n221), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n765), .C2(G159), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n827), .B1(new_n772), .B2(G50), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n484), .A2(new_n737), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n754), .B2(G68), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n737), .A2(new_n769), .B1(new_n750), .B2(new_n581), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n754), .A2(G303), .B1(G311), .B2(new_n777), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n772), .A2(G317), .ZN(new_n1022));
  INV_X1    g0822(.A(G322), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1021), .B(new_n1022), .C1(new_n1023), .C2(new_n764), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n756), .A2(new_n463), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1030), .B(new_n412), .C1(G326), .C2(new_n747), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1019), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1012), .B1(new_n1033), .B2(new_n734), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n672), .B2(new_n798), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n725), .A2(KEYINPUT112), .A3(new_n981), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n681), .C1(new_n725), .C2(new_n981), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT112), .B1(new_n725), .B2(new_n981), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1035), .B1(new_n729), .B2(new_n981), .C1(new_n1037), .C2(new_n1038), .ZN(G393));
  OR2_X1    g0839(.A1(new_n979), .A2(new_n982), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n682), .B1(new_n979), .B2(new_n982), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n979), .A2(new_n730), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n785), .B1(new_n533), .B2(new_n207), .C1(new_n941), .C2(new_n243), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n795), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT113), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n772), .A2(G311), .B1(new_n765), .B2(G317), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT52), .Z(new_n1048));
  AOI22_X1  g0848(.A1(new_n464), .A2(new_n828), .B1(new_n777), .B2(G303), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1049), .A2(new_n301), .A3(new_n757), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n754), .B2(G294), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n750), .A2(new_n769), .B1(new_n746), .B2(new_n1023), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT114), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1048), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n742), .A2(new_n822), .B1(new_n764), .B2(new_n255), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT51), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n758), .A2(new_n830), .B1(new_n750), .B2(new_n202), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n737), .A2(new_n221), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n756), .A2(new_n217), .B1(new_n746), .B2(new_n821), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n827), .B(new_n1060), .C1(new_n754), .C2(new_n316), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1056), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1054), .A2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1046), .B1(new_n735), .B2(new_n1063), .C1(new_n987), .C2(new_n798), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1042), .A2(new_n1043), .A3(new_n1064), .ZN(G390));
  NAND2_X1  g0865(.A1(new_n690), .A2(new_n691), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n637), .B1(new_n648), .B2(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n700), .A2(new_n701), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n671), .B(new_n809), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n915), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(KEYINPUT115), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT115), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(new_n1072), .A3(new_n915), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n878), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n912), .B1(new_n898), .B2(new_n872), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n912), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n917), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n908), .B2(new_n910), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n723), .A2(G330), .A3(new_n809), .A4(new_n878), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n908), .A2(new_n910), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1082), .A2(new_n1078), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1083));
  INV_X1    g0883(.A(G330), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n720), .B2(new_n880), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n879), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1081), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n453), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT116), .B1(new_n921), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n702), .B(new_n637), .C1(new_n648), .C2(new_n1066), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n687), .B1(new_n1091), .B2(new_n671), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n651), .A2(new_n687), .A3(new_n671), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n453), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AND4_X1   g0894(.A1(KEYINPUT116), .A2(new_n1094), .A3(new_n632), .A4(new_n1089), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1085), .A2(new_n809), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n878), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1097), .A2(new_n1100), .A3(new_n1080), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n916), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n723), .A2(G330), .A3(new_n809), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1103), .A2(new_n1099), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1101), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1096), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n682), .B1(new_n1088), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1087), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1110), .A2(new_n1096), .A3(new_n1105), .A4(new_n1081), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n730), .A3(new_n1081), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n795), .B1(new_n316), .B2(new_n843), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n772), .A2(G132), .B1(new_n765), .B2(G128), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT119), .Z(new_n1116));
  NAND2_X1  g0916(.A1(new_n747), .A2(G125), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n282), .B1(new_n756), .B2(new_n830), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT117), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1119), .B2(new_n1118), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT118), .Z(new_n1122));
  INV_X1    g0922(.A(new_n750), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(G150), .ZN(new_n1124));
  XOR2_X1   g0924(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n818), .B2(new_n758), .C1(new_n822), .C2(new_n737), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n753), .A2(new_n1128), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1129));
  NOR4_X1   g0929(.A1(new_n1116), .A2(new_n1122), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1131), .A2(KEYINPUT121), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n301), .B1(new_n746), .B2(new_n581), .C1(new_n217), .C2(new_n750), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n772), .B2(G116), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n754), .A2(G97), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n765), .A2(G283), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n756), .A2(new_n202), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1137), .B(new_n1058), .C1(G107), .C2(new_n777), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1131), .A2(KEYINPUT121), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1132), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1114), .B1(new_n1141), .B2(new_n734), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT122), .Z(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n911), .B2(new_n783), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1113), .A2(KEYINPUT123), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT123), .B1(new_n1113), .B2(new_n1144), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1112), .B1(new_n1146), .B2(new_n1147), .ZN(G378));
  NAND2_X1  g0948(.A1(new_n858), .A2(new_n268), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n297), .B(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1084), .B1(new_n899), .B2(new_n881), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n888), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT105), .B1(new_n882), .B2(new_n883), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n885), .B(KEYINPUT40), .C1(new_n874), .C2(new_n881), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1153), .B(new_n1152), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n920), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1153), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1152), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n920), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1163), .A3(new_n1157), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n729), .B1(new_n1159), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1161), .A2(new_n782), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n731), .B1(new_n843), .B2(G50), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n756), .A2(new_n201), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G77), .B2(new_n1123), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n533), .B2(new_n758), .C1(new_n764), .C2(new_n792), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n484), .A2(new_n753), .B1(new_n742), .B2(new_n223), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n274), .B1(new_n746), .B2(new_n769), .C1(new_n737), .C2(new_n202), .ZN(new_n1172));
  OR4_X1    g0972(.A1(new_n412), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n274), .B1(new_n827), .B2(new_n245), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1173), .A2(new_n1174), .B1(new_n830), .B2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G150), .A2(new_n828), .B1(new_n777), .B2(G132), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n753), .B2(new_n818), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n742), .A2(new_n1180), .B1(new_n750), .B2(new_n1128), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT124), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1179), .B(new_n1182), .C1(G125), .C2(new_n765), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT59), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1177), .B1(new_n822), .B2(new_n756), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1176), .B1(new_n1174), .B2(new_n1173), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1167), .B1(new_n1187), .B2(new_n734), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1166), .A2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT125), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1165), .A2(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1159), .A2(new_n1164), .B1(new_n1111), .B2(new_n1096), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n681), .B1(new_n1192), .B2(KEYINPUT57), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1105), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1096), .B1(new_n1088), .B2(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1162), .A2(new_n1163), .A3(new_n1157), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1163), .B1(new_n1162), .B2(new_n1157), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(KEYINPUT57), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1191), .B1(new_n1193), .B2(new_n1199), .ZN(G375));
  INV_X1    g1000(.A(new_n1096), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1194), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(new_n985), .A3(new_n1106), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1099), .A2(new_n782), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n754), .A2(G107), .B1(new_n464), .B2(new_n777), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n581), .B2(new_n764), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT126), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n282), .B1(new_n747), .B2(G303), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n221), .B2(new_n756), .C1(new_n533), .C2(new_n750), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1017), .B(new_n1209), .C1(G283), .C2(new_n772), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G137), .A2(new_n772), .B1(new_n754), .B2(G150), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1168), .B(new_n827), .C1(G128), .C2(new_n747), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n765), .A2(G132), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n758), .A2(new_n1128), .B1(new_n750), .B2(new_n822), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G50), .B2(new_n828), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n735), .B1(new_n1211), .B2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n796), .B(new_n1218), .C1(new_n202), .C2(new_n842), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1105), .A2(new_n730), .B1(new_n1204), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1203), .A2(new_n1220), .ZN(G381));
  AND3_X1   g1021(.A1(new_n1042), .A2(new_n1043), .A3(new_n1064), .ZN(new_n1222));
  INV_X1    g1022(.A(G384), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  OR2_X1    g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  OR4_X1    g1025(.A1(G387), .A2(new_n1224), .A3(G381), .A4(new_n1225), .ZN(new_n1226));
  OR3_X1    g1026(.A1(new_n1226), .A2(G378), .A3(G375), .ZN(G407));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n661), .A2(G213), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(G407), .B(G213), .C1(G375), .C2(new_n1231), .ZN(G409));
  NAND2_X1  g1032(.A1(new_n1106), .A2(KEYINPUT60), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1202), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1201), .A2(new_n1194), .A3(KEYINPUT60), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n681), .A3(new_n1235), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1236), .A2(G384), .A3(new_n1220), .ZN(new_n1237));
  AOI21_X1  g1037(.A(G384), .B1(new_n1236), .B2(new_n1220), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G2897), .B(new_n1230), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1220), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1223), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1236), .A2(G384), .A3(new_n1220), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1230), .A2(G2897), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1189), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT127), .B1(new_n1165), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n730), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT127), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1189), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1192), .A2(new_n985), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1248), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1228), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G378), .B(new_n1191), .C1(new_n1193), .C2(new_n1199), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1229), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT61), .B1(new_n1246), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT63), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1259), .B1(new_n1257), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1222), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(G393), .B(new_n800), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G390), .B(new_n967), .C1(new_n986), .C2(new_n998), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1230), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(KEYINPUT63), .A3(new_n1260), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1258), .A2(new_n1262), .A3(new_n1268), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1269), .A2(new_n1272), .A3(new_n1260), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1269), .B2(new_n1245), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1272), .B1(new_n1269), .B2(new_n1260), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1273), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1271), .B1(new_n1277), .B2(new_n1268), .ZN(G405));
  AND2_X1   g1078(.A1(G375), .A2(new_n1228), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1255), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1261), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1260), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1282), .A2(new_n1268), .A3(new_n1283), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(G402));
endmodule


