//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  INV_X1    g001(.A(G469), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G227), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n189), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI211_X1 g011(.A(KEYINPUT76), .B(KEYINPUT1), .C1(new_n194), .C2(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(G128), .A3(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n205), .A3(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n199), .A2(KEYINPUT77), .A3(new_n201), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G107), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G104), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n212), .A3(G104), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n215), .A2(new_n217), .A3(new_n209), .A4(new_n211), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n219));
  OR2_X1    g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n214), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n208), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n214), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n218), .A2(new_n219), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n218), .A2(new_n219), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n195), .A2(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n201), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n229), .A3(new_n206), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT11), .ZN(new_n232));
  INV_X1    g046(.A(G134), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(G137), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(G137), .ZN(new_n235));
  INV_X1    g049(.A(G137), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT11), .A3(G134), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G131), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT64), .B(G131), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n240), .A2(new_n235), .A3(new_n234), .A4(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT12), .B1(new_n231), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT12), .ZN(new_n244));
  INV_X1    g058(.A(new_n242), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n244), .B(new_n245), .C1(new_n223), .C2(new_n230), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n215), .A2(new_n217), .A3(new_n211), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G101), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n225), .B2(new_n226), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n200), .A2(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT0), .B(G128), .Z(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n200), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n248), .A3(G101), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n256), .A2(KEYINPUT75), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(KEYINPUT75), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n251), .A2(new_n255), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n229), .A2(new_n206), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n222), .A2(KEYINPUT10), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT10), .B1(new_n208), .B2(new_n222), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n242), .B(KEYINPUT78), .Z(new_n264));
  NOR3_X1   g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n193), .B1(new_n247), .B2(new_n265), .ZN(new_n266));
  OR3_X1    g080(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n192), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT10), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n199), .A2(KEYINPUT77), .A3(new_n201), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT77), .B1(new_n199), .B2(new_n201), .ZN(new_n271));
  INV_X1    g085(.A(new_n206), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n269), .B1(new_n273), .B2(new_n227), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n274), .A2(KEYINPUT79), .A3(new_n259), .A4(new_n261), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT79), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n262), .B2(new_n263), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n245), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n266), .B1(new_n268), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n188), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n259), .A2(new_n261), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT79), .B1(new_n282), .B2(new_n274), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n262), .A2(new_n263), .A3(new_n276), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n242), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n192), .B1(new_n285), .B2(new_n267), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n267), .B(new_n192), .C1(new_n243), .C2(new_n246), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n188), .B(new_n280), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT80), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n193), .B1(new_n278), .B2(new_n265), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n292), .B2(new_n287), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT80), .A3(new_n188), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n281), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(KEYINPUT9), .B(G234), .Z(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n187), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n279), .A2(new_n280), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G469), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n292), .A2(new_n287), .ZN(new_n303));
  AND4_X1   g117(.A1(KEYINPUT80), .A2(new_n303), .A3(new_n188), .A4(new_n280), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT80), .B1(new_n293), .B2(new_n188), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT81), .A3(new_n298), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G214), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT2), .B(G113), .Z(new_n311));
  XNOR2_X1  g125(.A(G116), .B(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT65), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n312), .B2(new_n311), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(new_n251), .A3(new_n258), .A4(new_n257), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n320), .A2(KEYINPUT5), .A3(G119), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n312), .B2(KEYINPUT5), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G113), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n222), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(G110), .B(G122), .Z(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n326), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n319), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(KEYINPUT6), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n255), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(G125), .B2(new_n260), .ZN(new_n333));
  INV_X1    g147(.A(G953), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G224), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n333), .B(new_n335), .Z(new_n336));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n325), .A2(new_n337), .A3(new_n326), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n330), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n332), .A2(KEYINPUT82), .B1(KEYINPUT7), .B2(new_n335), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n340), .B(new_n333), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n317), .A2(new_n323), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(new_n222), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n326), .B(KEYINPUT8), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n341), .B(new_n329), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n280), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G210), .B1(G237), .B2(G902), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT83), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n339), .A2(new_n280), .A3(new_n345), .A4(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n310), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G125), .B(G140), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT16), .ZN(new_n354));
  OR3_X1    g168(.A1(new_n331), .A2(KEYINPUT16), .A3(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G146), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(G146), .A3(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G237), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n334), .A3(G214), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(new_n194), .ZN(new_n364));
  INV_X1    g178(.A(new_n240), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(KEYINPUT17), .A3(new_n365), .ZN(new_n366));
  OR3_X1    g180(.A1(new_n364), .A2(KEYINPUT86), .A3(new_n365), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n365), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT86), .B1(new_n364), .B2(new_n365), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n361), .B(new_n366), .C1(new_n370), .C2(KEYINPUT17), .ZN(new_n371));
  XNOR2_X1  g185(.A(G113), .B(G122), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(new_n210), .ZN(new_n373));
  NAND3_X1  g187(.A1(KEYINPUT85), .A2(KEYINPUT18), .A3(G131), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n364), .B(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n353), .B(new_n357), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n353), .B(KEYINPUT19), .Z(new_n380));
  OAI21_X1  g194(.A(new_n359), .B1(new_n380), .B2(G146), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT87), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n383), .B(new_n359), .C1(new_n380), .C2(G146), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n370), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT88), .B1(new_n385), .B2(new_n377), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(new_n373), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(KEYINPUT88), .A3(new_n377), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n379), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n391));
  INV_X1    g205(.A(G475), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .A4(new_n280), .ZN(new_n393));
  INV_X1    g207(.A(new_n388), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n394), .A2(new_n386), .A3(new_n373), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n392), .B(new_n280), .C1(new_n395), .C2(new_n379), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n373), .B1(new_n371), .B2(new_n377), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n280), .B1(new_n379), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT89), .B(G475), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(G234), .A2(G237), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(G952), .A3(new_n334), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT21), .B(G898), .Z(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(G902), .A3(G953), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G128), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT13), .B1(new_n412), .B2(G143), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n233), .ZN(new_n414));
  XNOR2_X1  g228(.A(G128), .B(G143), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G116), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT90), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n418), .A2(new_n212), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n212), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n212), .ZN(new_n422));
  INV_X1    g236(.A(G122), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT14), .B1(new_n423), .B2(G116), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n320), .B2(G122), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n423), .A2(KEYINPUT14), .A3(G116), .ZN(new_n426));
  OAI21_X1  g240(.A(G107), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n415), .B(new_n233), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n422), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G217), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n297), .A2(new_n431), .A3(G953), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n421), .A2(new_n429), .A3(new_n432), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n280), .ZN(new_n437));
  INV_X1    g251(.A(G478), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT15), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n439), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n405), .A2(new_n411), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n308), .A2(new_n352), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT91), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n412), .A2(G119), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT23), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n446), .B1(KEYINPUT72), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G119), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G128), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT72), .B(KEYINPUT23), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n448), .B(new_n450), .C1(new_n451), .C2(new_n446), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G110), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT73), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n450), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT71), .ZN(new_n457));
  MUX2_X1   g271(.A(KEYINPUT71), .B(new_n457), .S(new_n446), .Z(new_n458));
  XOR2_X1   g272(.A(KEYINPUT24), .B(G110), .Z(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n360), .A3(new_n460), .ZN(new_n461));
  OAI22_X1  g275(.A1(new_n458), .A2(new_n459), .B1(new_n452), .B2(G110), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n353), .A2(new_n357), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n359), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n334), .A2(G221), .A3(G234), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT22), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(G137), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n465), .B(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n431), .B1(G234), .B2(new_n280), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(G902), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n280), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT25), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(KEYINPUT25), .A3(new_n280), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n472), .B1(new_n477), .B2(new_n470), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(G472), .A2(G902), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT67), .ZN(new_n481));
  INV_X1    g295(.A(new_n235), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n233), .A2(G137), .ZN(new_n483));
  OAI21_X1  g297(.A(G131), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n241), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n241), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n260), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n242), .A2(new_n255), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT66), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT66), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n242), .A2(new_n490), .A3(new_n255), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT68), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n260), .A2(new_n241), .A3(new_n484), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n488), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n493), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n242), .A2(new_n490), .A3(new_n255), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n490), .B1(new_n242), .B2(new_n255), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT68), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT30), .A4(new_n487), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n494), .A2(new_n318), .A3(new_n497), .A4(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n318), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n504), .A3(new_n487), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT26), .B(G101), .Z(new_n506));
  NAND3_X1  g320(.A1(new_n362), .A2(new_n334), .A3(G210), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n503), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n511), .A2(KEYINPUT31), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT31), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n503), .A2(new_n513), .A3(new_n505), .A4(new_n510), .ZN(new_n514));
  INV_X1    g328(.A(new_n510), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n496), .A2(new_n318), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n487), .A2(new_n488), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT28), .B1(new_n519), .B2(new_n504), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n515), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n480), .B1(new_n512), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT32), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n511), .A2(KEYINPUT31), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n514), .A3(new_n521), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(KEYINPUT32), .A3(new_n480), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(KEYINPUT70), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n530), .A3(new_n524), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n503), .A2(new_n505), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n515), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n510), .B1(new_n518), .B2(new_n520), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT29), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n492), .A2(new_n318), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n505), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n520), .B1(new_n539), .B2(KEYINPUT28), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT29), .A3(new_n510), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n280), .ZN(new_n542));
  OAI21_X1  g356(.A(G472), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n479), .B1(new_n532), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n352), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n300), .B2(new_n307), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n443), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n445), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(G101), .ZN(G3));
  INV_X1    g364(.A(new_n523), .ZN(new_n551));
  INV_X1    g365(.A(G472), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n527), .B2(new_n280), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI211_X1 g369(.A(new_n479), .B(new_n555), .C1(new_n300), .C2(new_n307), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n436), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n434), .A2(KEYINPUT33), .A3(new_n435), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n558), .A2(G478), .A3(new_n280), .A4(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT93), .B(G478), .Z(new_n565));
  NAND2_X1  g379(.A1(new_n437), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n405), .A2(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n310), .B(new_n411), .C1(new_n349), .C2(new_n351), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n556), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT34), .B(G104), .Z(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(G6));
  INV_X1    g388(.A(new_n397), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n390), .A2(new_n392), .A3(new_n280), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n398), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n442), .A2(new_n404), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n352), .A2(new_n577), .A3(new_n578), .A4(new_n410), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n569), .A2(new_n581), .A3(new_n577), .A4(new_n578), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n556), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(new_n212), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT95), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n586), .B(KEYINPUT35), .Z(G9));
  NAND2_X1  g401(.A1(new_n477), .A2(new_n470), .ZN(new_n588));
  INV_X1    g402(.A(new_n468), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(KEYINPUT36), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n465), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n471), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n554), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT96), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n445), .A2(new_n548), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT97), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT37), .B(G110), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G12));
  NAND2_X1  g413(.A1(new_n532), .A2(new_n543), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n334), .A2(G900), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n406), .A2(G902), .ZN(new_n603));
  OR3_X1    g417(.A1(new_n602), .A2(KEYINPUT98), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT98), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n407), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n398), .B2(new_n576), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n578), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n546), .A2(new_n600), .A3(new_n593), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G128), .ZN(G30));
  NAND2_X1  g426(.A1(new_n349), .A2(new_n351), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n613), .B(KEYINPUT38), .Z(new_n614));
  NAND2_X1  g428(.A1(new_n405), .A2(new_n442), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n310), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n606), .B(KEYINPUT39), .Z(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n308), .A2(new_n619), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n614), .B(new_n617), .C1(new_n620), .C2(KEYINPUT40), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n539), .A2(KEYINPUT99), .A3(new_n515), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n511), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT99), .B1(new_n539), .B2(new_n515), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n280), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(G472), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n593), .B1(new_n532), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n621), .B(new_n627), .C1(KEYINPUT40), .C2(new_n620), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G143), .ZN(G45));
  NAND4_X1  g443(.A1(new_n405), .A2(new_n593), .A3(new_n567), .A4(new_n606), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n308), .A2(new_n631), .A3(new_n600), .A4(new_n352), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n546), .A2(KEYINPUT100), .A3(new_n600), .A4(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G146), .ZN(G48));
  NAND2_X1  g451(.A1(new_n303), .A2(new_n280), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n639), .A3(G469), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT101), .B1(new_n293), .B2(new_n188), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n291), .A2(new_n294), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n298), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n641), .A2(new_n640), .B1(new_n291), .B2(new_n294), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n298), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n544), .A3(new_n571), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT41), .B(G113), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G15));
  AOI21_X1  g466(.A(KEYINPUT102), .B1(new_n647), .B2(new_n298), .ZN(new_n653));
  AND4_X1   g467(.A1(KEYINPUT102), .A2(new_n642), .A3(new_n643), .A4(new_n298), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n544), .B(new_n583), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n649), .A2(KEYINPUT103), .A3(new_n544), .A4(new_n583), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G116), .ZN(G18));
  NOR2_X1   g474(.A1(new_n644), .A2(new_n545), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n661), .A2(new_n600), .A3(new_n443), .A4(new_n593), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G119), .ZN(G21));
  OAI21_X1  g477(.A(new_n514), .B1(new_n510), .B2(new_n540), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n480), .B1(new_n512), .B2(new_n664), .ZN(new_n665));
  AOI211_X1 g479(.A(KEYINPUT104), .B(new_n552), .C1(new_n527), .C2(new_n280), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n280), .B1(new_n512), .B2(new_n522), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n668), .B2(G472), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n478), .B(new_n665), .C1(new_n666), .C2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n615), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n671), .B(new_n569), .C1(new_n653), .C2(new_n654), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G122), .ZN(G24));
  OAI21_X1  g487(.A(new_n665), .B1(new_n666), .B2(new_n669), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n630), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n661), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G125), .ZN(G27));
  NOR2_X1   g491(.A1(new_n568), .A2(new_n607), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n295), .A2(new_n299), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n613), .A2(new_n310), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AND4_X1   g496(.A1(new_n679), .A2(new_n306), .A3(new_n298), .A4(new_n681), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n678), .B(new_n544), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n680), .A2(new_n679), .A3(new_n681), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n306), .A2(new_n298), .A3(new_n681), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT105), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n525), .A2(KEYINPUT106), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n528), .A3(new_n543), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n525), .A2(KEYINPUT106), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n479), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n690), .A2(new_n695), .A3(KEYINPUT42), .A4(new_n678), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n686), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G131), .ZN(G33));
  OAI211_X1 g512(.A(new_n544), .B(new_n610), .C1(new_n682), .C2(new_n683), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT107), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n690), .A2(new_n701), .A3(new_n544), .A4(new_n610), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G134), .ZN(G36));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n705));
  INV_X1    g519(.A(new_n567), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n405), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT43), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n555), .A3(new_n593), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n705), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n710), .A2(KEYINPUT109), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(KEYINPUT109), .ZN(new_n712));
  OAI221_X1 g526(.A(new_n681), .B1(new_n705), .B2(new_n709), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT110), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n279), .B(KEYINPUT45), .ZN(new_n715));
  OAI21_X1  g529(.A(G469), .B1(new_n715), .B2(G902), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT46), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n643), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT108), .Z(new_n719));
  NOR2_X1   g533(.A1(new_n716), .A2(KEYINPUT46), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n298), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n618), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n714), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT111), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G137), .ZN(G39));
  XNOR2_X1  g539(.A(new_n721), .B(KEYINPUT47), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n600), .A2(new_n478), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n678), .A3(new_n681), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G140), .ZN(G42));
  INV_X1    g544(.A(new_n407), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n708), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n647), .A2(new_n298), .A3(new_n681), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n734), .A2(new_n479), .A3(new_n694), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT118), .Z(new_n736));
  INV_X1    g550(.A(KEYINPUT119), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT48), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n739), .A2(KEYINPUT48), .ZN(new_n741));
  NOR4_X1   g555(.A1(new_n732), .A2(new_n310), .A3(new_n613), .A4(new_n670), .ZN(new_n742));
  INV_X1    g556(.A(new_n647), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n298), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n742), .B1(new_n727), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n532), .A2(new_n626), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n733), .A2(new_n746), .A3(new_n479), .A4(new_n407), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n393), .A2(new_n398), .B1(new_n401), .B2(new_n403), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n747), .A2(new_n748), .A3(new_n706), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n674), .B(new_n734), .C1(new_n588), .C2(new_n592), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n732), .A2(new_n644), .A3(new_n670), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n751), .A2(new_n310), .A3(new_n614), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT50), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(KEYINPUT50), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n749), .B(new_n750), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n745), .A2(new_n755), .A3(KEYINPUT51), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n334), .A2(G952), .ZN(new_n757));
  INV_X1    g571(.A(new_n568), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n757), .B1(new_n747), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n740), .A2(new_n741), .A3(new_n756), .A4(new_n759), .ZN(new_n760));
  OAI22_X1  g574(.A1(new_n726), .A2(KEYINPUT117), .B1(new_n298), .B2(new_n743), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n726), .A2(KEYINPUT117), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n742), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n763), .B2(new_n755), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n751), .A2(new_n352), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n690), .A2(new_n675), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n697), .A2(new_n703), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n549), .A2(new_n659), .A3(new_n650), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n748), .A2(new_n442), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n570), .B1(new_n568), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n308), .A2(new_n478), .A3(new_n554), .A4(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n772), .A2(new_n672), .A3(new_n662), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n596), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n442), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n600), .A2(new_n775), .A3(new_n404), .A4(new_n593), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n681), .A2(new_n608), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n300), .B2(new_n307), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n777), .B1(new_n776), .B2(new_n779), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n768), .A2(new_n769), .A3(new_n774), .A4(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n308), .A2(new_n600), .A3(new_n352), .A4(new_n593), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n676), .B1(new_n784), .B2(new_n609), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n616), .A2(new_n613), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n680), .A3(new_n606), .A4(new_n627), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n636), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n636), .A3(KEYINPUT114), .A4(new_n788), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n783), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n785), .B1(new_n634), .B2(new_n635), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT114), .B1(new_n799), .B2(new_n788), .ZN(new_n800));
  INV_X1    g614(.A(new_n793), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT52), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n794), .A3(new_n783), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT53), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n798), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n783), .A2(new_n794), .A3(KEYINPUT53), .A4(new_n797), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT116), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n803), .A2(new_n809), .A3(new_n796), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n803), .B2(new_n796), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n807), .B(new_n808), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n765), .A2(new_n766), .A3(new_n805), .A4(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(G952), .B2(G953), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n478), .A2(new_n309), .A3(new_n298), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n743), .B2(KEYINPUT49), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n743), .A2(KEYINPUT49), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n816), .B1(new_n817), .B2(KEYINPUT112), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(KEYINPUT112), .B2(new_n817), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n614), .A3(new_n707), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n814), .B1(new_n746), .B2(new_n820), .ZN(G75));
  OR2_X1    g635(.A1(new_n810), .A2(new_n811), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n280), .B1(new_n822), .B2(new_n807), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT56), .B1(new_n823), .B2(new_n348), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n330), .A2(new_n338), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(new_n336), .Z(new_n826));
  XNOR2_X1  g640(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  AOI211_X1 g644(.A(KEYINPUT56), .B(new_n828), .C1(new_n823), .C2(new_n348), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n334), .A2(G952), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(G51));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n806), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n806), .A2(new_n834), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n835), .B(new_n836), .C1(new_n810), .C2(new_n811), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n812), .ZN(new_n839));
  NAND2_X1  g653(.A1(G469), .A2(G902), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT57), .Z(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n303), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n823), .A2(G469), .A3(new_n715), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n832), .B1(new_n843), .B2(new_n844), .ZN(G54));
  NAND3_X1  g659(.A1(new_n823), .A2(KEYINPUT58), .A3(G475), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(new_n389), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n389), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n847), .A2(new_n848), .A3(new_n832), .ZN(G60));
  OAI21_X1  g663(.A(new_n805), .B1(new_n837), .B2(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(G478), .A2(G902), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT59), .Z(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n558), .A2(new_n559), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n852), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT121), .B1(new_n839), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n861));
  INV_X1    g675(.A(new_n859), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n861), .B(new_n862), .C1(new_n838), .C2(new_n812), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n858), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n832), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n856), .B1(new_n850), .B2(new_n853), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n855), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n867), .ZN(G63));
  NAND2_X1  g682(.A1(G217), .A2(G902), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT60), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n837), .A2(new_n591), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n822), .B2(new_n807), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n865), .B(new_n872), .C1(new_n873), .C2(new_n469), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT61), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n874), .B(new_n876), .ZN(G66));
  NOR2_X1   g691(.A1(new_n769), .A2(new_n774), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(G953), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n334), .B1(new_n408), .B2(G224), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n825), .B1(G898), .B2(new_n334), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(G69));
  AOI21_X1  g699(.A(new_n601), .B1(new_n190), .B2(G953), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n601), .B(KEYINPUT126), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n494), .A2(new_n497), .A3(new_n502), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(new_n380), .Z(new_n889));
  AND2_X1   g703(.A1(new_n723), .A2(new_n729), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n697), .A2(new_n703), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n799), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n722), .A2(new_n695), .A3(new_n787), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(KEYINPUT127), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n894), .A2(KEYINPUT127), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n890), .A2(new_n892), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n887), .B(new_n889), .C1(new_n897), .C2(new_n334), .ZN(new_n898));
  INV_X1    g712(.A(new_n544), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n308), .A2(new_n619), .A3(new_n681), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n899), .B(new_n900), .C1(new_n568), .C2(new_n770), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n723), .A2(new_n729), .A3(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n901), .A2(new_n902), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n628), .A2(new_n799), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT62), .Z(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n334), .A3(new_n889), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n886), .B1(new_n898), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n889), .B1(new_n897), .B2(new_n334), .ZN(new_n912));
  INV_X1    g726(.A(new_n887), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n886), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n915), .A3(new_n909), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n916), .ZN(G72));
  NOR2_X1   g731(.A1(new_n534), .A2(new_n515), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n904), .A2(new_n905), .A3(new_n907), .A4(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n897), .B2(new_n535), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n832), .B1(new_n920), .B2(new_n878), .ZN(new_n921));
  INV_X1    g735(.A(new_n535), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n918), .ZN(new_n923));
  NAND2_X1  g737(.A1(G472), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT63), .Z(new_n925));
  OR2_X1    g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n798), .A2(new_n804), .A3(new_n925), .A4(new_n923), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n921), .A2(new_n926), .A3(new_n927), .ZN(G57));
endmodule


