

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U552 ( .A1(G299), .A2(n730), .ZN(n728) );
  INV_X1 U553 ( .A(KEYINPUT27), .ZN(n707) );
  XOR2_X1 U554 ( .A(KEYINPUT95), .B(n699), .Z(n709) );
  NAND2_X1 U555 ( .A1(n692), .A2(n796), .ZN(n694) );
  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n796) );
  INV_X1 U557 ( .A(G2105), .ZN(n533) );
  OR2_X1 U558 ( .A1(n775), .A2(n774), .ZN(n820) );
  NOR2_X1 U559 ( .A1(G651), .A2(n646), .ZN(n654) );
  NOR2_X2 U560 ( .A1(n557), .A2(n556), .ZN(G160) );
  INV_X1 U561 ( .A(G651), .ZN(n523) );
  NOR2_X1 U562 ( .A1(G543), .A2(n523), .ZN(n520) );
  XOR2_X1 U563 ( .A(KEYINPUT1), .B(n520), .Z(n657) );
  NAND2_X1 U564 ( .A1(G65), .A2(n657), .ZN(n522) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n646) );
  NAND2_X1 U566 ( .A1(G53), .A2(n654), .ZN(n521) );
  NAND2_X1 U567 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U569 ( .A1(G91), .A2(n653), .ZN(n526) );
  OR2_X1 U570 ( .A1(n523), .A2(n646), .ZN(n524) );
  XOR2_X1 U571 ( .A(KEYINPUT68), .B(n524), .Z(n661) );
  NAND2_X1 U572 ( .A1(G78), .A2(n661), .ZN(n525) );
  NAND2_X1 U573 ( .A1(n526), .A2(n525), .ZN(n527) );
  OR2_X1 U574 ( .A1(n528), .A2(n527), .ZN(G299) );
  INV_X1 U575 ( .A(G2104), .ZN(n532) );
  NOR2_X4 U576 ( .A1(G2105), .A2(n532), .ZN(n886) );
  NAND2_X1 U577 ( .A1(G102), .A2(n886), .ZN(n531) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X2 U579 ( .A(KEYINPUT17), .B(n529), .Z(n887) );
  NAND2_X1 U580 ( .A1(G138), .A2(n887), .ZN(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n538) );
  NOR2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n882) );
  NAND2_X1 U583 ( .A1(G114), .A2(n882), .ZN(n536) );
  NOR2_X1 U584 ( .A1(n533), .A2(G2104), .ZN(n534) );
  XNOR2_X1 U585 ( .A(n534), .B(KEYINPUT66), .ZN(n883) );
  NAND2_X1 U586 ( .A1(G126), .A2(n883), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U588 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U589 ( .A1(n653), .A2(G89), .ZN(n539) );
  XNOR2_X1 U590 ( .A(n539), .B(KEYINPUT4), .ZN(n541) );
  NAND2_X1 U591 ( .A1(G76), .A2(n661), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U593 ( .A(KEYINPUT5), .B(n542), .ZN(n548) );
  NAND2_X1 U594 ( .A1(n657), .A2(G63), .ZN(n543) );
  XOR2_X1 U595 ( .A(KEYINPUT75), .B(n543), .Z(n545) );
  NAND2_X1 U596 ( .A1(n654), .A2(G51), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U598 ( .A(KEYINPUT6), .B(n546), .Z(n547) );
  NAND2_X1 U599 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U600 ( .A(KEYINPUT7), .B(n549), .ZN(G168) );
  XOR2_X1 U601 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U602 ( .A1(G101), .A2(n886), .ZN(n550) );
  XNOR2_X1 U603 ( .A(n550), .B(KEYINPUT23), .ZN(n551) );
  XNOR2_X1 U604 ( .A(n551), .B(KEYINPUT67), .ZN(n553) );
  NAND2_X1 U605 ( .A1(G113), .A2(n882), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U607 ( .A1(G137), .A2(n887), .ZN(n555) );
  NAND2_X1 U608 ( .A1(G125), .A2(n883), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U610 ( .A(G2443), .B(G2446), .Z(n559) );
  XNOR2_X1 U611 ( .A(G2427), .B(G2451), .ZN(n558) );
  XNOR2_X1 U612 ( .A(n559), .B(n558), .ZN(n565) );
  XOR2_X1 U613 ( .A(G2430), .B(G2454), .Z(n561) );
  XNOR2_X1 U614 ( .A(G1341), .B(G1348), .ZN(n560) );
  XNOR2_X1 U615 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U616 ( .A(G2435), .B(G2438), .Z(n562) );
  XNOR2_X1 U617 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U618 ( .A(n565), .B(n564), .Z(n566) );
  AND2_X1 U619 ( .A1(G14), .A2(n566), .ZN(G401) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U623 ( .A(n567), .B(KEYINPUT72), .ZN(n568) );
  XOR2_X1 U624 ( .A(KEYINPUT10), .B(n568), .Z(n913) );
  NAND2_X1 U625 ( .A1(n913), .A2(G567), .ZN(n569) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U627 ( .A1(n657), .A2(G56), .ZN(n570) );
  XNOR2_X1 U628 ( .A(KEYINPUT14), .B(n570), .ZN(n576) );
  NAND2_X1 U629 ( .A1(n653), .A2(G81), .ZN(n571) );
  XNOR2_X1 U630 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G68), .A2(n661), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U633 ( .A(KEYINPUT13), .B(n574), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U635 ( .A(n577), .B(KEYINPUT73), .ZN(n579) );
  NAND2_X1 U636 ( .A1(n654), .A2(G43), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n579), .A2(n578), .ZN(n915) );
  INV_X1 U638 ( .A(G860), .ZN(n601) );
  OR2_X1 U639 ( .A1(n915), .A2(n601), .ZN(G153) );
  NAND2_X1 U640 ( .A1(G64), .A2(n657), .ZN(n581) );
  NAND2_X1 U641 ( .A1(G52), .A2(n654), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n587) );
  NAND2_X1 U643 ( .A1(G90), .A2(n653), .ZN(n583) );
  NAND2_X1 U644 ( .A1(G77), .A2(n661), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U646 ( .A(KEYINPUT9), .B(n584), .Z(n585) );
  XNOR2_X1 U647 ( .A(KEYINPUT70), .B(n585), .ZN(n586) );
  NOR2_X1 U648 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U649 ( .A(KEYINPUT71), .B(n588), .Z(G171) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G301), .A2(G868), .ZN(n589) );
  XNOR2_X1 U652 ( .A(n589), .B(KEYINPUT74), .ZN(n598) );
  INV_X1 U653 ( .A(G868), .ZN(n674) );
  NAND2_X1 U654 ( .A1(G66), .A2(n657), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G92), .A2(n653), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U657 ( .A1(n654), .A2(G54), .ZN(n593) );
  NAND2_X1 U658 ( .A1(G79), .A2(n661), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U661 ( .A(KEYINPUT15), .B(n596), .ZN(n914) );
  NAND2_X1 U662 ( .A1(n674), .A2(n914), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n598), .A2(n597), .ZN(G284) );
  NOR2_X1 U664 ( .A1(G286), .A2(n674), .ZN(n600) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n599) );
  NOR2_X1 U666 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n601), .A2(G559), .ZN(n602) );
  INV_X1 U668 ( .A(n914), .ZN(n719) );
  NAND2_X1 U669 ( .A1(n602), .A2(n719), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n603), .B(KEYINPUT16), .ZN(n604) );
  XNOR2_X1 U671 ( .A(KEYINPUT76), .B(n604), .ZN(G148) );
  NOR2_X1 U672 ( .A1(n914), .A2(n674), .ZN(n605) );
  XNOR2_X1 U673 ( .A(n605), .B(KEYINPUT77), .ZN(n606) );
  NOR2_X1 U674 ( .A1(G559), .A2(n606), .ZN(n608) );
  NOR2_X1 U675 ( .A1(G868), .A2(n915), .ZN(n607) );
  NOR2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U677 ( .A(KEYINPUT78), .B(n609), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G99), .A2(n886), .ZN(n611) );
  NAND2_X1 U679 ( .A1(G111), .A2(n882), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n611), .A2(n610), .ZN(n618) );
  NAND2_X1 U681 ( .A1(n883), .A2(G123), .ZN(n612) );
  XOR2_X1 U682 ( .A(KEYINPUT79), .B(n612), .Z(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT18), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G135), .A2(n887), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U686 ( .A(KEYINPUT80), .B(n616), .ZN(n617) );
  NOR2_X1 U687 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U688 ( .A(n619), .B(KEYINPUT81), .ZN(n999) );
  XOR2_X1 U689 ( .A(G2096), .B(KEYINPUT82), .Z(n620) );
  XNOR2_X1 U690 ( .A(n999), .B(n620), .ZN(n621) );
  INV_X1 U691 ( .A(G2100), .ZN(n851) );
  NAND2_X1 U692 ( .A1(n621), .A2(n851), .ZN(G156) );
  NAND2_X1 U693 ( .A1(n719), .A2(G559), .ZN(n671) );
  XNOR2_X1 U694 ( .A(n915), .B(n671), .ZN(n622) );
  NOR2_X1 U695 ( .A1(n622), .A2(G860), .ZN(n629) );
  NAND2_X1 U696 ( .A1(G67), .A2(n657), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G93), .A2(n653), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n654), .A2(G55), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G80), .A2(n661), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n627) );
  OR2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n673) );
  XOR2_X1 U703 ( .A(n629), .B(n673), .Z(G145) );
  NAND2_X1 U704 ( .A1(G48), .A2(n654), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT84), .ZN(n637) );
  NAND2_X1 U706 ( .A1(G61), .A2(n657), .ZN(n632) );
  NAND2_X1 U707 ( .A1(G86), .A2(n653), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n661), .A2(G73), .ZN(n633) );
  XOR2_X1 U710 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U713 ( .A(KEYINPUT85), .B(n638), .Z(G305) );
  NAND2_X1 U714 ( .A1(G62), .A2(n657), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G75), .A2(n661), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n653), .A2(G88), .ZN(n641) );
  XOR2_X1 U718 ( .A(KEYINPUT86), .B(n641), .Z(n642) );
  NOR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n654), .A2(G50), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(G303) );
  INV_X1 U722 ( .A(G303), .ZN(G166) );
  NAND2_X1 U723 ( .A1(G49), .A2(n654), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G87), .A2(n646), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n657), .A2(n649), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n650) );
  XOR2_X1 U728 ( .A(KEYINPUT83), .B(n650), .Z(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U730 ( .A1(G85), .A2(n653), .ZN(n656) );
  NAND2_X1 U731 ( .A1(G47), .A2(n654), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U733 ( .A1(G60), .A2(n657), .ZN(n658) );
  XNOR2_X1 U734 ( .A(KEYINPUT69), .B(n658), .ZN(n659) );
  NOR2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U736 ( .A1(G72), .A2(n661), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n663), .A2(n662), .ZN(G290) );
  XNOR2_X1 U738 ( .A(n915), .B(G305), .ZN(n670) );
  XOR2_X1 U739 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n665) );
  XOR2_X1 U740 ( .A(G299), .B(G166), .Z(n664) );
  XNOR2_X1 U741 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n666), .B(G288), .ZN(n667) );
  XOR2_X1 U743 ( .A(n673), .B(n667), .Z(n668) );
  XNOR2_X1 U744 ( .A(n668), .B(G290), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n670), .B(n669), .ZN(n902) );
  XNOR2_X1 U746 ( .A(n671), .B(n902), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n672), .A2(G868), .ZN(n676) );
  NAND2_X1 U748 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U749 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U754 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n682) );
  NAND2_X1 U757 ( .A1(G132), .A2(G82), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U759 ( .A1(n683), .A2(G96), .ZN(n684) );
  NOR2_X1 U760 ( .A1(n684), .A2(G218), .ZN(n685) );
  XNOR2_X1 U761 ( .A(n685), .B(KEYINPUT89), .ZN(n838) );
  NAND2_X1 U762 ( .A1(n838), .A2(G2106), .ZN(n689) );
  NAND2_X1 U763 ( .A1(G69), .A2(G120), .ZN(n686) );
  NOR2_X1 U764 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U765 ( .A1(G108), .A2(n687), .ZN(n839) );
  NAND2_X1 U766 ( .A1(n839), .A2(G567), .ZN(n688) );
  NAND2_X1 U767 ( .A1(n689), .A2(n688), .ZN(n840) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n690) );
  NOR2_X1 U769 ( .A1(n840), .A2(n690), .ZN(n837) );
  NAND2_X1 U770 ( .A1(n837), .A2(G36), .ZN(G176) );
  NOR2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n759) );
  NOR2_X1 U772 ( .A1(G1971), .A2(G303), .ZN(n691) );
  NOR2_X1 U773 ( .A1(n759), .A2(n691), .ZN(n923) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n795) );
  INV_X1 U775 ( .A(n795), .ZN(n692) );
  INV_X1 U776 ( .A(KEYINPUT64), .ZN(n693) );
  XNOR2_X2 U777 ( .A(n694), .B(n693), .ZN(n712) );
  INV_X1 U778 ( .A(n712), .ZN(n742) );
  NAND2_X1 U779 ( .A1(n742), .A2(G8), .ZN(n778) );
  NOR2_X1 U780 ( .A1(G1966), .A2(n778), .ZN(n751) );
  NOR2_X1 U781 ( .A1(n742), .A2(G2084), .ZN(n752) );
  NOR2_X1 U782 ( .A1(n751), .A2(n752), .ZN(n695) );
  NAND2_X1 U783 ( .A1(G8), .A2(n695), .ZN(n696) );
  XNOR2_X1 U784 ( .A(KEYINPUT30), .B(n696), .ZN(n697) );
  NOR2_X1 U785 ( .A1(G168), .A2(n697), .ZN(n698) );
  XNOR2_X1 U786 ( .A(n698), .B(KEYINPUT99), .ZN(n704) );
  NOR2_X1 U787 ( .A1(G1961), .A2(n712), .ZN(n702) );
  XOR2_X1 U788 ( .A(G2078), .B(KEYINPUT25), .Z(n975) );
  INV_X1 U789 ( .A(n712), .ZN(n699) );
  NOR2_X1 U790 ( .A1(n975), .A2(n709), .ZN(n700) );
  XNOR2_X1 U791 ( .A(n700), .B(KEYINPUT96), .ZN(n701) );
  NOR2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n735) );
  NAND2_X1 U793 ( .A1(n735), .A2(G301), .ZN(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n706) );
  XOR2_X1 U795 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n705) );
  XNOR2_X1 U796 ( .A(n706), .B(n705), .ZN(n739) );
  INV_X1 U797 ( .A(n709), .ZN(n720) );
  NAND2_X1 U798 ( .A1(G2072), .A2(n720), .ZN(n708) );
  XNOR2_X1 U799 ( .A(n708), .B(n707), .ZN(n711) );
  XOR2_X1 U800 ( .A(G1956), .B(KEYINPUT97), .Z(n945) );
  NAND2_X1 U801 ( .A1(n709), .A2(n945), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n730) );
  AND2_X1 U803 ( .A1(n712), .A2(G1996), .ZN(n714) );
  XNOR2_X1 U804 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n713) );
  XNOR2_X1 U805 ( .A(n714), .B(n713), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n742), .A2(G1341), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U808 ( .A1(n915), .A2(n717), .ZN(n718) );
  OR2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n726) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n724) );
  NAND2_X1 U811 ( .A1(G2067), .A2(n720), .ZN(n722) );
  NAND2_X1 U812 ( .A1(n742), .A2(G1348), .ZN(n721) );
  NAND2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U817 ( .A(n729), .B(KEYINPUT98), .ZN(n733) );
  NAND2_X1 U818 ( .A1(G299), .A2(n730), .ZN(n731) );
  XNOR2_X1 U819 ( .A(KEYINPUT28), .B(n731), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U821 ( .A(n734), .B(KEYINPUT29), .ZN(n737) );
  NOR2_X1 U822 ( .A1(G301), .A2(n735), .ZN(n736) );
  NOR2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n750) );
  INV_X1 U825 ( .A(n750), .ZN(n740) );
  NAND2_X1 U826 ( .A1(n740), .A2(G286), .ZN(n747) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n778), .ZN(n741) );
  XNOR2_X1 U828 ( .A(n741), .B(KEYINPUT102), .ZN(n744) );
  NOR2_X1 U829 ( .A1(n742), .A2(G2090), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U831 ( .A1(n745), .A2(G303), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U833 ( .A1(G8), .A2(n748), .ZN(n749) );
  XNOR2_X1 U834 ( .A(KEYINPUT32), .B(n749), .ZN(n757) );
  NOR2_X1 U835 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U836 ( .A1(G8), .A2(n752), .ZN(n753) );
  NAND2_X1 U837 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U838 ( .A(n755), .B(KEYINPUT101), .Z(n756) );
  NAND2_X1 U839 ( .A1(n757), .A2(n756), .ZN(n767) );
  NAND2_X1 U840 ( .A1(n923), .A2(n767), .ZN(n758) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n922) );
  NAND2_X1 U842 ( .A1(n758), .A2(n922), .ZN(n764) );
  XOR2_X1 U843 ( .A(G1981), .B(G305), .Z(n933) );
  INV_X1 U844 ( .A(n933), .ZN(n762) );
  NAND2_X1 U845 ( .A1(n759), .A2(KEYINPUT33), .ZN(n760) );
  NOR2_X1 U846 ( .A1(n778), .A2(n760), .ZN(n761) );
  OR2_X1 U847 ( .A1(n762), .A2(n761), .ZN(n770) );
  OR2_X1 U848 ( .A1(n778), .A2(n770), .ZN(n763) );
  NOR2_X1 U849 ( .A1(n764), .A2(n763), .ZN(n775) );
  NAND2_X1 U850 ( .A1(G8), .A2(G166), .ZN(n765) );
  NOR2_X1 U851 ( .A1(G2090), .A2(n765), .ZN(n766) );
  XNOR2_X1 U852 ( .A(n766), .B(KEYINPUT103), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n769), .A2(n778), .ZN(n773) );
  INV_X1 U855 ( .A(n770), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n771), .A2(KEYINPUT33), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U859 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U860 ( .A1(n778), .A2(n777), .ZN(n818) );
  NAND2_X1 U861 ( .A1(G117), .A2(n882), .ZN(n780) );
  NAND2_X1 U862 ( .A1(G129), .A2(n883), .ZN(n779) );
  NAND2_X1 U863 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U864 ( .A1(n886), .A2(G105), .ZN(n781) );
  XOR2_X1 U865 ( .A(KEYINPUT38), .B(n781), .Z(n782) );
  NOR2_X1 U866 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U867 ( .A1(n887), .A2(G141), .ZN(n784) );
  NAND2_X1 U868 ( .A1(n785), .A2(n784), .ZN(n893) );
  NOR2_X1 U869 ( .A1(G1996), .A2(n893), .ZN(n997) );
  XOR2_X1 U870 ( .A(KEYINPUT92), .B(G1991), .Z(n974) );
  NAND2_X1 U871 ( .A1(G95), .A2(n886), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G107), .A2(n882), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U874 ( .A1(G119), .A2(n883), .ZN(n788) );
  XNOR2_X1 U875 ( .A(KEYINPUT91), .B(n788), .ZN(n789) );
  NOR2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n887), .A2(G131), .ZN(n791) );
  AND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n877) );
  NOR2_X1 U879 ( .A1(n974), .A2(n877), .ZN(n794) );
  AND2_X1 U880 ( .A1(n893), .A2(G1996), .ZN(n793) );
  NOR2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n1013) );
  NOR2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n821) );
  XNOR2_X1 U883 ( .A(KEYINPUT93), .B(n821), .ZN(n797) );
  NOR2_X1 U884 ( .A1(n1013), .A2(n797), .ZN(n822) );
  AND2_X1 U885 ( .A1(n974), .A2(n877), .ZN(n1011) );
  NOR2_X1 U886 ( .A1(G1986), .A2(G290), .ZN(n798) );
  NOR2_X1 U887 ( .A1(n1011), .A2(n798), .ZN(n799) );
  NOR2_X1 U888 ( .A1(n822), .A2(n799), .ZN(n800) );
  NOR2_X1 U889 ( .A1(n997), .A2(n800), .ZN(n801) );
  XNOR2_X1 U890 ( .A(KEYINPUT39), .B(n801), .ZN(n812) );
  XNOR2_X1 U891 ( .A(KEYINPUT37), .B(G2067), .ZN(n813) );
  NAND2_X1 U892 ( .A1(G116), .A2(n882), .ZN(n803) );
  NAND2_X1 U893 ( .A1(G128), .A2(n883), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U895 ( .A(n804), .B(KEYINPUT35), .ZN(n809) );
  NAND2_X1 U896 ( .A1(G104), .A2(n886), .ZN(n806) );
  NAND2_X1 U897 ( .A1(G140), .A2(n887), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U899 ( .A(KEYINPUT34), .B(n807), .Z(n808) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U901 ( .A(n810), .B(KEYINPUT36), .Z(n897) );
  NOR2_X1 U902 ( .A1(n813), .A2(n897), .ZN(n1014) );
  NAND2_X1 U903 ( .A1(n1014), .A2(n821), .ZN(n811) );
  XNOR2_X1 U904 ( .A(n811), .B(KEYINPUT90), .ZN(n824) );
  NAND2_X1 U905 ( .A1(n812), .A2(n824), .ZN(n815) );
  AND2_X1 U906 ( .A1(n813), .A2(n897), .ZN(n814) );
  XOR2_X1 U907 ( .A(KEYINPUT104), .B(n814), .Z(n1005) );
  NAND2_X1 U908 ( .A1(n815), .A2(n1005), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n816), .A2(n821), .ZN(n829) );
  INV_X1 U910 ( .A(n829), .ZN(n817) );
  OR2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n831) );
  XNOR2_X1 U913 ( .A(G1986), .B(G290), .ZN(n928) );
  AND2_X1 U914 ( .A1(n928), .A2(n821), .ZN(n827) );
  INV_X1 U915 ( .A(n822), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U917 ( .A(n825), .B(KEYINPUT94), .ZN(n826) );
  OR2_X1 U918 ( .A1(n827), .A2(n826), .ZN(n828) );
  AND2_X1 U919 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U920 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U921 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n913), .ZN(G217) );
  NAND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n834) );
  INV_X1 U924 ( .A(G661), .ZN(n833) );
  NOR2_X1 U925 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U926 ( .A(n835), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U928 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U930 ( .A(G132), .ZN(G219) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G82), .ZN(G220) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n840), .ZN(G319) );
  XNOR2_X1 U938 ( .A(G1981), .B(KEYINPUT41), .ZN(n850) );
  XOR2_X1 U939 ( .A(G1956), .B(G1961), .Z(n842) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1966), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U942 ( .A(G1976), .B(G1971), .Z(n844) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U945 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U946 ( .A(KEYINPUT106), .B(G2474), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(G229) );
  XNOR2_X1 U949 ( .A(n851), .B(G2096), .ZN(n853) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(G2678), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U952 ( .A(KEYINPUT43), .B(G2090), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U958 ( .A1(G136), .A2(n887), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G112), .A2(n882), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n868) );
  NAND2_X1 U961 ( .A1(G100), .A2(n886), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(KEYINPUT108), .ZN(n866) );
  XOR2_X1 U963 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n864) );
  NAND2_X1 U964 ( .A1(G124), .A2(n883), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U967 ( .A1(n868), .A2(n867), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G103), .A2(n886), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G139), .A2(n887), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U971 ( .A1(G115), .A2(n882), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G127), .A2(n883), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U974 ( .A(KEYINPUT47), .B(n873), .ZN(n874) );
  XNOR2_X1 U975 ( .A(KEYINPUT109), .B(n874), .ZN(n875) );
  NOR2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n1001) );
  XNOR2_X1 U977 ( .A(n877), .B(n1001), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n878), .B(G162), .ZN(n879) );
  XOR2_X1 U979 ( .A(n879), .B(KEYINPUT48), .Z(n881) );
  XNOR2_X1 U980 ( .A(G164), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n896) );
  NAND2_X1 U982 ( .A1(G118), .A2(n882), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G130), .A2(n883), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n892) );
  NAND2_X1 U985 ( .A1(G106), .A2(n886), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G142), .A2(n887), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U988 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U989 ( .A1(n892), .A2(n891), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U991 ( .A(n896), .B(n895), .Z(n899) );
  XOR2_X1 U992 ( .A(G160), .B(n897), .Z(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U994 ( .A(n900), .B(n999), .Z(n901) );
  NOR2_X1 U995 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U996 ( .A(n902), .B(KEYINPUT110), .ZN(n904) );
  XOR2_X1 U997 ( .A(n914), .B(G286), .Z(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U999 ( .A(n905), .B(G171), .Z(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n907), .B(KEYINPUT49), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n908), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n909), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(KEYINPUT111), .B(n910), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  INV_X1 U1010 ( .A(n913), .ZN(G223) );
  XNOR2_X1 U1011 ( .A(G16), .B(KEYINPUT56), .ZN(n939) );
  XOR2_X1 U1012 ( .A(n914), .B(G1348), .Z(n919) );
  XOR2_X1 U1013 ( .A(G171), .B(G1961), .Z(n917) );
  XNOR2_X1 U1014 ( .A(n915), .B(G1341), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n931) );
  XOR2_X1 U1017 ( .A(G299), .B(G1956), .Z(n921) );
  NAND2_X1 U1018 ( .A1(G1971), .A2(G303), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n925) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1022 ( .A(KEYINPUT120), .B(n926), .Z(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(n929), .B(KEYINPUT121), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(KEYINPUT122), .B(n932), .ZN(n937) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G168), .ZN(n934) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(KEYINPUT57), .B(n935), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1031 ( .A1(n939), .A2(n938), .ZN(n967) );
  XNOR2_X1 U1032 ( .A(G16), .B(KEYINPUT123), .ZN(n965) );
  XOR2_X1 U1033 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n963) );
  XOR2_X1 U1034 ( .A(G1966), .B(G21), .Z(n950) );
  XNOR2_X1 U1035 ( .A(G1348), .B(KEYINPUT59), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(n940), .B(G4), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G1341), .B(G19), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(G6), .B(G1981), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(G20), .B(n945), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT60), .B(n948), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(KEYINPUT124), .B(G1961), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(G5), .B(n951), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n961) );
  XNOR2_X1 U1048 ( .A(G1986), .B(G24), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G22), .B(G1971), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G1976), .B(KEYINPUT125), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n956), .B(G23), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1054 ( .A(KEYINPUT58), .B(n959), .Z(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n963), .B(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n994) );
  XNOR2_X1 U1059 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n989) );
  XNOR2_X1 U1060 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G32), .B(G1996), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(G28), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(KEYINPUT116), .B(G2072), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(G33), .B(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n979) );
  XOR2_X1 U1067 ( .A(n974), .B(G25), .Z(n977) );
  XNOR2_X1 U1068 ( .A(G27), .B(n975), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(KEYINPUT53), .B(n980), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G2090), .B(G35), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(n981), .B(KEYINPUT115), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n984), .B(KEYINPUT117), .ZN(n987) );
  XOR2_X1 U1076 ( .A(G2084), .B(G34), .Z(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT54), .B(n985), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(n989), .B(n988), .ZN(n990) );
  OR2_X1 U1080 ( .A1(G29), .A2(n990), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n991), .ZN(n992) );
  XOR2_X1 U1082 ( .A(KEYINPUT119), .B(n992), .Z(n993) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(KEYINPUT127), .ZN(n1025) );
  INV_X1 U1085 ( .A(G29), .ZN(n1023) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1088 ( .A(KEYINPUT51), .B(n998), .Z(n1000) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1008) );
  XOR2_X1 U1090 ( .A(G2072), .B(n1001), .Z(n1003) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1017) );
  XOR2_X1 U1096 ( .A(G160), .B(G2084), .Z(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT112), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(KEYINPUT114), .B(n1018), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(KEYINPUT52), .B(KEYINPUT113), .Z(n1019) );
  XNOR2_X1 U1104 ( .A(n1020), .B(n1019), .ZN(n1021) );
  NOR2_X1 U1105 ( .A1(KEYINPUT55), .A2(n1021), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1026), .Z(G150) );
  INV_X1 U1109 ( .A(G150), .ZN(G311) );
endmodule

