//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n211));
  AOI21_X1  g010(.A(G36gat), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n209), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT15), .B1(new_n212), .B2(new_n213), .ZN(new_n215));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n215), .A2(new_n216), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT17), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n221), .B1(new_n217), .B2(new_n218), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n207), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n219), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(new_n207), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT18), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n207), .B(new_n219), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n224), .B(KEYINPUT13), .Z(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n223), .A2(new_n226), .A3(KEYINPUT18), .A4(new_n224), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT11), .B(G169gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n237), .B(new_n238), .Z(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n229), .A2(new_n233), .A3(new_n241), .A4(new_n234), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  OR2_X1    g045(.A1(G141gat), .A2(G148gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(G141gat), .A2(G148gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT75), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT75), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(new_n251), .A3(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253));
  OR2_X1    g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(KEYINPUT2), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n250), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT2), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n247), .A2(new_n257), .A3(new_n248), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(KEYINPUT74), .ZN(new_n259));
  OR3_X1    g058(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .A4(new_n253), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G211gat), .A2(G218gat), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n267), .A2(KEYINPUT22), .ZN(new_n268));
  XNOR2_X1  g067(.A(G197gat), .B(G204gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n266), .A2(new_n271), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n263), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n262), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n272), .A2(new_n273), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n256), .A2(new_n275), .A3(new_n261), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n263), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G228gat), .ZN(new_n282));
  INV_X1    g081(.A(G233gat), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n276), .A2(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n266), .B(new_n271), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT3), .B1(new_n286), .B2(new_n263), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n285), .B(new_n280), .C1(new_n287), .C2(new_n262), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT82), .B(G22gat), .Z(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G78gat), .B(G106gat), .Z(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT81), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT31), .B(G50gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n284), .A2(new_n288), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(G22gat), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT83), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n290), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT84), .ZN(new_n300));
  INV_X1    g099(.A(new_n289), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  AOI211_X1 g101(.A(KEYINPUT84), .B(new_n289), .C1(new_n284), .C2(new_n288), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n294), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n297), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G183gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(G190gat), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT24), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(new_n308), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  XOR2_X1   g115(.A(KEYINPUT65), .B(KEYINPUT23), .Z(new_n317));
  OAI211_X1 g116(.A(new_n312), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G169gat), .ZN(new_n319));
  INV_X1    g118(.A(G176gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n316), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n316), .B(KEYINPUT66), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT23), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(KEYINPUT25), .A3(new_n322), .ZN(new_n329));
  OAI22_X1  g128(.A1(new_n326), .A2(KEYINPUT25), .B1(new_n329), .B2(new_n318), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n321), .B1(KEYINPUT26), .B2(new_n323), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n313), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT27), .B(G183gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n308), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT68), .B1(new_n336), .B2(KEYINPUT67), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT28), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n334), .B(new_n339), .C1(new_n337), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n330), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT29), .B1(new_n330), .B2(new_n342), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n277), .ZN(new_n348));
  XOR2_X1   g147(.A(G8gat), .B(G36gat), .Z(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT72), .ZN(new_n350));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n345), .B(new_n286), .C1(new_n344), .C2(new_n346), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n348), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT30), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT30), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n348), .A2(new_n354), .A3(new_n357), .A4(new_n353), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n348), .A2(new_n354), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n352), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n360), .A2(KEYINPUT73), .A3(new_n352), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n359), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G113gat), .ZN(new_n367));
  INV_X1    g166(.A(G120gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G113gat), .A2(G120gat), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT1), .ZN(new_n372));
  XOR2_X1   g171(.A(G127gat), .B(G134gat), .Z(new_n373));
  OAI211_X1 g172(.A(new_n371), .B(new_n372), .C1(new_n373), .C2(KEYINPUT69), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(new_n372), .A3(new_n370), .ZN(new_n375));
  XNOR2_X1  g174(.A(G127gat), .B(G134gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n370), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT69), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n375), .B(new_n376), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n256), .A2(new_n261), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT4), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n374), .A2(new_n379), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n262), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n278), .A3(new_n380), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n262), .A2(KEYINPUT77), .A3(new_n383), .A4(new_n384), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n392), .B(KEYINPUT76), .Z(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(KEYINPUT39), .ZN(new_n395));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT0), .ZN(new_n397));
  XNOR2_X1  g196(.A(G57gat), .B(G85gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n262), .A2(new_n384), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n380), .A2(new_n381), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n394), .B(KEYINPUT39), .C1(new_n393), .C2(new_n404), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n401), .A2(KEYINPUT40), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT40), .B1(new_n401), .B2(new_n405), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n390), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n409));
  INV_X1    g208(.A(new_n393), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n389), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT78), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n389), .A2(new_n409), .A3(new_n410), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n390), .A4(new_n387), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n382), .A2(new_n385), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(new_n410), .A3(new_n389), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n409), .B1(new_n404), .B2(new_n393), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n412), .A2(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(new_n399), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n406), .A2(new_n407), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n307), .B1(new_n366), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT37), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n348), .B2(new_n354), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT86), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n352), .B1(new_n360), .B2(KEYINPUT37), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(KEYINPUT38), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n426), .A2(KEYINPUT87), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT87), .B1(new_n426), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n419), .B2(new_n399), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n415), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n418), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n434), .A2(new_n399), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(KEYINPUT6), .B2(new_n420), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT38), .B1(new_n427), .B2(new_n424), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n355), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n422), .B1(new_n431), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n343), .A2(new_n384), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n330), .A2(new_n342), .A3(new_n380), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n445), .B(KEYINPUT64), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n446), .A3(new_n443), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT32), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT32), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n451), .A3(new_n447), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(G15gat), .B(G43gat), .Z(new_n458));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n455), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n457), .B1(new_n455), .B2(new_n460), .ZN(new_n462));
  OR3_X1    g261(.A1(new_n453), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n453), .B1(new_n461), .B2(new_n462), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT36), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT79), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n433), .B2(new_n436), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n434), .A2(new_n435), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n400), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n419), .A2(new_n399), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n471), .A2(KEYINPUT79), .A3(new_n432), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n420), .A2(KEYINPUT6), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n475), .A2(new_n365), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n475), .B2(new_n365), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n307), .B(KEYINPUT85), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n441), .B(new_n467), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n294), .B1(new_n299), .B2(new_n304), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n463), .B(new_n464), .C1(new_n482), .C2(new_n297), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT35), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n359), .A2(new_n363), .A3(new_n484), .A4(new_n364), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n483), .A2(new_n485), .A3(new_n438), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n477), .A2(new_n478), .A3(new_n483), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(new_n484), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n246), .B1(new_n481), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(G57gat), .A2(G64gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(G57gat), .A2(G64gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(KEYINPUT9), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G71gat), .A2(G78gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(G71gat), .A2(G78gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(KEYINPUT89), .A3(new_n492), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n499));
  AND2_X1   g298(.A1(G57gat), .A2(G64gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(G57gat), .A2(G64gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n494), .B1(new_n496), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n503), .A2(KEYINPUT90), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT90), .B1(new_n503), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n497), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT21), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT91), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(G183gat), .B(G211gat), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT92), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n513), .B(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n207), .B1(new_n509), .B2(new_n508), .ZN(new_n517));
  XNOR2_X1  g316(.A(G127gat), .B(G155gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n517), .B(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n521), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT8), .ZN(new_n526));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G85gat), .ZN(new_n530));
  INV_X1    g329(.A(G92gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n526), .A2(new_n529), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G99gat), .B(G106gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n538));
  AND3_X1   g337(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g340(.A1(KEYINPUT8), .A2(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n535), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n534), .A2(new_n536), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT94), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n220), .B2(new_n222), .ZN(new_n549));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT93), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n219), .A2(new_n547), .B1(KEYINPUT41), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT95), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n554), .A2(new_n556), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n552), .A2(KEYINPUT41), .ZN(new_n560));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n557), .B2(new_n558), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n524), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n545), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n570), .B(new_n497), .C1(new_n506), .C2(new_n507), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT96), .B(KEYINPUT10), .ZN(new_n572));
  INV_X1    g371(.A(new_n497), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n500), .A2(new_n501), .A3(new_n499), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT89), .B1(new_n491), .B2(new_n492), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n505), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT90), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n503), .A2(KEYINPUT90), .A3(new_n505), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n573), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n571), .B(new_n572), .C1(new_n580), .C2(new_n547), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT97), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n548), .A2(new_n508), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n571), .A4(new_n572), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(KEYINPUT10), .A3(new_n547), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n580), .A2(KEYINPUT98), .A3(KEYINPUT10), .A4(new_n547), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n582), .A2(new_n585), .B1(new_n589), .B2(new_n590), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT99), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n583), .B2(new_n571), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT100), .ZN(new_n600));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  NAND3_X1  g402(.A1(new_n598), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n586), .A2(new_n591), .B1(G230gat), .B2(G233gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  INV_X1    g406(.A(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n490), .A2(new_n568), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(new_n475), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n365), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT16), .B(G8gat), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n206), .B2(new_n615), .ZN(new_n618));
  MUX2_X1   g417(.A(new_n617), .B(new_n618), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g418(.A(G15gat), .B1(new_n612), .B2(new_n467), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n465), .A2(G15gat), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n612), .B2(new_n621), .ZN(G1326gat));
  NOR2_X1   g421(.A1(new_n612), .A2(new_n480), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT43), .B(G22gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(G1327gat));
  INV_X1    g424(.A(KEYINPUT44), .ZN(new_n626));
  AOI211_X1 g425(.A(new_n626), .B(new_n566), .C1(new_n481), .C2(new_n489), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n522), .A2(new_n523), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n610), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n245), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n475), .A2(new_n365), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT80), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n475), .A2(new_n365), .A3(new_n476), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n307), .A2(new_n465), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n486), .B1(new_n635), .B2(KEYINPUT35), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI211_X1 g437(.A(KEYINPUT101), .B(new_n486), .C1(new_n635), .C2(KEYINPUT35), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n481), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n567), .ZN(new_n641));
  AOI211_X1 g440(.A(new_n627), .B(new_n630), .C1(new_n641), .C2(new_n626), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(G29gat), .B1(new_n643), .B2(new_n475), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n628), .A2(new_n566), .A3(new_n610), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n490), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n475), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n209), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT45), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(new_n650), .ZN(G1328gat));
  OAI21_X1  g450(.A(G36gat), .B1(new_n643), .B2(new_n365), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n646), .A2(G36gat), .A3(new_n365), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT46), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(G1329gat));
  INV_X1    g454(.A(new_n465), .ZN(new_n656));
  AOI21_X1  g455(.A(G43gat), .B1(new_n647), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n466), .A2(G43gat), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n642), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT47), .Z(G1330gat));
  NAND2_X1  g459(.A1(new_n441), .A2(new_n467), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n479), .A2(new_n480), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n489), .A2(KEYINPUT101), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n636), .A2(new_n637), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n626), .B1(new_n666), .B2(new_n566), .ZN(new_n667));
  INV_X1    g466(.A(new_n627), .ZN(new_n668));
  INV_X1    g467(.A(new_n630), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n667), .A2(new_n307), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n627), .B1(new_n641), .B2(new_n626), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n673), .A2(KEYINPUT104), .A3(new_n307), .A4(new_n669), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n674), .A3(G50gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n480), .ZN(new_n676));
  INV_X1    g475(.A(G50gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT102), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n647), .A2(KEYINPUT103), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n678), .B(KEYINPUT102), .Z(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n646), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT48), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n675), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n667), .A2(new_n676), .A3(new_n668), .A4(new_n669), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G50gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n647), .A2(new_n679), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT48), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n687), .A2(KEYINPUT105), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n677), .B1(new_n670), .B2(new_n671), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n685), .B1(new_n696), .B2(new_n674), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT48), .B1(new_n689), .B2(new_n690), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n699), .ZN(G1331gat));
  NOR4_X1   g499(.A1(new_n524), .A2(new_n245), .A3(new_n567), .A4(new_n611), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n640), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n475), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g503(.A(new_n702), .B(KEYINPUT106), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n365), .B(KEYINPUT107), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT49), .B(G64gat), .Z(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n708), .B2(new_n710), .ZN(G1333gat));
  NAND3_X1  g510(.A1(new_n705), .A2(G71gat), .A3(new_n466), .ZN(new_n712));
  INV_X1    g511(.A(G71gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n702), .B2(new_n465), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g515(.A1(new_n705), .A2(new_n676), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g517(.A1(new_n628), .A2(new_n245), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n640), .A2(KEYINPUT51), .A3(new_n567), .A4(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724));
  INV_X1    g523(.A(new_n719), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n641), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n727), .A2(new_n530), .A3(new_n648), .A4(new_n610), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n725), .A2(new_n611), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n673), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G85gat), .B1(new_n730), .B2(new_n475), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(G1336gat));
  NOR3_X1   g531(.A1(new_n706), .A2(G92gat), .A3(new_n611), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G92gat), .B1(new_n730), .B2(new_n706), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n673), .A2(new_n366), .A3(new_n729), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n726), .A2(new_n720), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n738), .A2(G92gat), .B1(new_n739), .B2(new_n733), .ZN(new_n740));
  OAI22_X1  g539(.A1(new_n734), .A2(new_n737), .B1(new_n736), .B2(new_n740), .ZN(G1337gat));
  NOR3_X1   g540(.A1(new_n465), .A2(new_n611), .A3(G99gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G99gat), .B1(new_n730), .B2(new_n467), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n743), .A2(KEYINPUT109), .A3(new_n744), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1338gat));
  INV_X1    g548(.A(new_n307), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n750), .A2(G106gat), .A3(new_n611), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n727), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G106gat), .B1(new_n730), .B2(new_n750), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n673), .A2(new_n676), .A3(new_n729), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n756), .A2(G106gat), .B1(new_n739), .B2(new_n751), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n752), .A2(new_n755), .B1(new_n754), .B2(new_n757), .ZN(G1339gat));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n603), .B1(new_n605), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n595), .B1(new_n596), .B2(KEYINPUT99), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n586), .A2(new_n591), .A3(KEYINPUT99), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n595), .B1(new_n589), .B2(new_n590), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n586), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT110), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n586), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(KEYINPUT54), .A3(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(KEYINPUT55), .B(new_n760), .C1(new_n763), .C2(new_n769), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n770), .A2(new_n245), .A3(new_n604), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n760), .B1(new_n763), .B2(new_n769), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n773), .B1(new_n772), .B2(new_n774), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n771), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n230), .A2(new_n232), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n224), .B1(new_n223), .B2(new_n226), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI211_X1 g580(.A(KEYINPUT112), .B(new_n224), .C1(new_n223), .C2(new_n226), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n239), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(new_n244), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n610), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n567), .B1(new_n777), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n783), .A2(new_n787), .A3(new_n244), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n783), .B2(new_n244), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n788), .A2(new_n789), .A3(new_n566), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n770), .A2(new_n604), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n790), .B(new_n791), .C1(new_n775), .C2(new_n776), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n524), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  NOR4_X1   g593(.A1(new_n524), .A2(new_n245), .A3(new_n567), .A4(new_n610), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  AOI211_X1 g595(.A(new_n475), .B(new_n483), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n706), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n367), .A3(new_n245), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n676), .B1(new_n794), .B2(new_n796), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n707), .A2(new_n475), .A3(new_n465), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n245), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n805), .A3(G113gat), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n805), .B1(new_n804), .B2(G113gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n799), .B1(new_n807), .B2(new_n808), .ZN(G1340gat));
  NAND2_X1  g608(.A1(new_n610), .A2(new_n368), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT115), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n798), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G120gat), .B1(new_n802), .B2(new_n611), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1341gat));
  INV_X1    g613(.A(G127gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n815), .A3(new_n628), .ZN(new_n816));
  OAI21_X1  g615(.A(G127gat), .B1(new_n802), .B2(new_n524), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1342gat));
  NAND2_X1  g617(.A1(new_n365), .A2(new_n567), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(G134gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n797), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(KEYINPUT56), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT116), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n803), .A2(new_n567), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n824), .A2(G134gat), .B1(KEYINPUT56), .B2(new_n821), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1343gat));
  AOI21_X1  g625(.A(new_n750), .B1(new_n794), .B2(new_n796), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n648), .A3(new_n467), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n828), .A2(KEYINPUT120), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(KEYINPUT120), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n707), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(G141gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n245), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n480), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n770), .A2(new_n245), .A3(new_n604), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n598), .A2(KEYINPUT54), .A3(new_n766), .A4(new_n768), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n838), .B2(new_n760), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n785), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n566), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n628), .B1(new_n841), .B2(new_n792), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n836), .B1(new_n842), .B2(new_n795), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(new_n836), .C1(new_n842), .C2(new_n795), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n844), .B(new_n846), .C1(new_n827), .C2(KEYINPUT57), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n707), .A2(new_n466), .A3(new_n475), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n245), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G141gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  NOR4_X1   g651(.A1(new_n828), .A2(G141gat), .A3(new_n246), .A4(new_n707), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(KEYINPUT118), .A3(G141gat), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n852), .B(new_n834), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n850), .A2(new_n854), .ZN(new_n858));
  INV_X1    g657(.A(new_n853), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT119), .B1(new_n860), .B2(KEYINPUT58), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n851), .B1(new_n857), .B2(new_n861), .ZN(G1344gat));
  INV_X1    g661(.A(G148gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n831), .A2(new_n863), .A3(new_n610), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n842), .A2(new_n795), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT121), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n480), .B1(new_n866), .B2(KEYINPUT121), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n827), .A2(KEYINPUT57), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n872), .B1(new_n869), .B2(new_n870), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n610), .B(new_n848), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n865), .B1(new_n874), .B2(G148gat), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n847), .A2(new_n848), .ZN(new_n876));
  AOI211_X1 g675(.A(KEYINPUT59), .B(new_n863), .C1(new_n876), .C2(new_n610), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n864), .B1(new_n875), .B2(new_n877), .ZN(G1345gat));
  AOI21_X1  g677(.A(G155gat), .B1(new_n831), .B2(new_n628), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n628), .A2(G155gat), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT123), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n879), .B1(new_n876), .B2(new_n881), .ZN(G1346gat));
  AOI211_X1 g681(.A(G162gat), .B(new_n819), .C1(new_n829), .C2(new_n830), .ZN(new_n883));
  INV_X1    g682(.A(G162gat), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n876), .B2(new_n567), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n883), .A2(new_n885), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n648), .A2(new_n365), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n800), .A2(new_n656), .A3(new_n887), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(new_n246), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(KEYINPUT125), .A3(G169gat), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT125), .B1(new_n889), .B2(G169gat), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n648), .B1(new_n794), .B2(new_n796), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n706), .A2(new_n483), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT124), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n245), .A2(new_n319), .ZN(new_n897));
  OAI22_X1  g696(.A1(new_n891), .A2(new_n892), .B1(new_n896), .B2(new_n897), .ZN(G1348gat));
  OAI21_X1  g697(.A(G176gat), .B1(new_n888), .B2(new_n611), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n610), .A2(new_n320), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n896), .B2(new_n900), .ZN(G1349gat));
  OAI21_X1  g700(.A(G183gat), .B1(new_n888), .B2(new_n524), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n628), .A2(new_n335), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n895), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g703(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n904), .B(new_n905), .Z(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n888), .B2(new_n566), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n907), .A2(KEYINPUT61), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n567), .A2(new_n308), .ZN(new_n911));
  OAI22_X1  g710(.A1(new_n909), .A2(new_n910), .B1(new_n896), .B2(new_n911), .ZN(G1351gat));
  XOR2_X1   g711(.A(KEYINPUT127), .B(G197gat), .Z(new_n913));
  NOR3_X1   g712(.A1(new_n466), .A2(new_n648), .A3(new_n365), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n871), .B2(new_n873), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n913), .B1(new_n915), .B2(new_n246), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n466), .A2(new_n706), .A3(new_n750), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n893), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n246), .A2(new_n913), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(G1352gat));
  OAI21_X1  g719(.A(G204gat), .B1(new_n915), .B2(new_n611), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n918), .A2(G204gat), .A3(new_n611), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT62), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1353gat));
  OR3_X1    g723(.A1(new_n918), .A2(G211gat), .A3(new_n524), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n628), .B(new_n914), .C1(new_n871), .C2(new_n873), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT63), .B1(new_n926), .B2(G211gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1354gat));
  OAI21_X1  g728(.A(G218gat), .B1(new_n915), .B2(new_n566), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n566), .A2(G218gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n918), .B2(new_n931), .ZN(G1355gat));
endmodule


