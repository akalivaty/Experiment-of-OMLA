

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X2 U553 ( .A(KEYINPUT72), .B(n617), .ZN(n1011) );
  AND2_X1 U554 ( .A1(n746), .A2(n679), .ZN(n685) );
  BUF_X1 U555 ( .A(n698), .Z(n699) );
  INV_X1 U556 ( .A(KEYINPUT28), .ZN(n604) );
  NOR2_X2 U557 ( .A1(G2105), .A2(n521), .ZN(n579) );
  XNOR2_X2 U558 ( .A(n522), .B(KEYINPUT65), .ZN(n692) );
  NOR2_X1 U559 ( .A1(n621), .A2(n620), .ZN(n636) );
  NAND2_X1 U560 ( .A1(n600), .A2(n599), .ZN(n646) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n644) );
  INV_X1 U562 ( .A(KEYINPUT91), .ZN(n660) );
  XNOR2_X1 U563 ( .A(n661), .B(n660), .ZN(n667) );
  NAND2_X1 U564 ( .A1(n596), .A2(n595), .ZN(n662) );
  NOR2_X1 U565 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  AND2_X1 U567 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U568 ( .A(KEYINPUT17), .B(n518), .Z(n698) );
  NOR2_X1 U569 ( .A1(n565), .A2(n531), .ZN(n792) );
  NOR2_X1 U570 ( .A1(G651), .A2(n565), .ZN(n795) );
  XNOR2_X1 U571 ( .A(KEYINPUT40), .B(KEYINPUT98), .ZN(n764) );
  INV_X1 U572 ( .A(G2104), .ZN(n521) );
  NAND2_X1 U573 ( .A1(G102), .A2(n579), .ZN(n520) );
  NAND2_X1 U574 ( .A1(G138), .A2(n698), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n520), .A2(n519), .ZN(n526) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U577 ( .A1(G114), .A2(n881), .ZN(n524) );
  NAND2_X1 U578 ( .A1(n521), .A2(G2105), .ZN(n522) );
  NAND2_X1 U579 ( .A1(G126), .A2(n692), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U581 ( .A1(n526), .A2(n525), .ZN(G164) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n565) );
  NAND2_X1 U583 ( .A1(G53), .A2(n795), .ZN(n529) );
  INV_X1 U584 ( .A(G651), .ZN(n531) );
  NOR2_X1 U585 ( .A1(G543), .A2(n531), .ZN(n527) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n527), .Z(n613) );
  NAND2_X1 U587 ( .A1(G65), .A2(n613), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U589 ( .A(KEYINPUT70), .B(n530), .Z(n535) );
  NOR2_X1 U590 ( .A1(G543), .A2(G651), .ZN(n791) );
  NAND2_X1 U591 ( .A1(G91), .A2(n791), .ZN(n533) );
  NAND2_X1 U592 ( .A1(G78), .A2(n792), .ZN(n532) );
  AND2_X1 U593 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U594 ( .A1(n535), .A2(n534), .ZN(G299) );
  NAND2_X1 U595 ( .A1(G52), .A2(n795), .ZN(n537) );
  NAND2_X1 U596 ( .A1(G64), .A2(n613), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n542) );
  NAND2_X1 U598 ( .A1(G90), .A2(n791), .ZN(n539) );
  NAND2_X1 U599 ( .A1(G77), .A2(n792), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U602 ( .A1(n542), .A2(n541), .ZN(G171) );
  NAND2_X1 U603 ( .A1(G89), .A2(n791), .ZN(n543) );
  XOR2_X1 U604 ( .A(KEYINPUT75), .B(n543), .Z(n544) );
  XNOR2_X1 U605 ( .A(n544), .B(KEYINPUT4), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G76), .A2(n792), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U608 ( .A(n547), .B(KEYINPUT5), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G51), .A2(n795), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G63), .A2(n613), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT6), .B(n550), .Z(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U614 ( .A(n553), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U615 ( .A(G168), .B(KEYINPUT8), .Z(n554) );
  XNOR2_X1 U616 ( .A(KEYINPUT76), .B(n554), .ZN(G286) );
  NAND2_X1 U617 ( .A1(G88), .A2(n791), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G75), .A2(n792), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G50), .A2(n795), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G62), .A2(n613), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U623 ( .A1(n560), .A2(n559), .ZN(G166) );
  INV_X1 U624 ( .A(G166), .ZN(G303) );
  NAND2_X1 U625 ( .A1(G49), .A2(n795), .ZN(n562) );
  NAND2_X1 U626 ( .A1(G74), .A2(G651), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n613), .A2(n563), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(KEYINPUT80), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G87), .A2(n565), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(G288) );
  NAND2_X1 U632 ( .A1(G86), .A2(n791), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G61), .A2(n613), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n792), .A2(G73), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT2), .B(n570), .Z(n571) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT81), .B(n573), .Z(n575) );
  NAND2_X1 U639 ( .A1(n795), .A2(G48), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(G305) );
  NAND2_X1 U641 ( .A1(G137), .A2(n698), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(KEYINPUT66), .ZN(n584) );
  NAND2_X1 U643 ( .A1(G113), .A2(n881), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G125), .A2(n692), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G101), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(KEYINPUT23), .B(n580), .ZN(n581) );
  NOR2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(KEYINPUT64), .B(n585), .Z(n596) );
  BUF_X1 U651 ( .A(n596), .Z(G160) );
  NAND2_X1 U652 ( .A1(G60), .A2(n613), .ZN(n586) );
  XOR2_X1 U653 ( .A(KEYINPUT68), .B(n586), .Z(n591) );
  NAND2_X1 U654 ( .A1(G85), .A2(n791), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G72), .A2(n792), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U657 ( .A(KEYINPUT67), .B(n589), .Z(n590) );
  NOR2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n795), .A2(G47), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n593), .A2(n592), .ZN(G290) );
  NOR2_X1 U661 ( .A1(G164), .A2(G1384), .ZN(n712) );
  AND2_X1 U662 ( .A1(G40), .A2(n712), .ZN(n595) );
  INV_X1 U663 ( .A(n662), .ZN(n598) );
  INV_X1 U664 ( .A(KEYINPUT87), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U666 ( .A1(KEYINPUT87), .A2(n662), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n646), .A2(G2072), .ZN(n601) );
  XNOR2_X1 U668 ( .A(n601), .B(KEYINPUT27), .ZN(n603) );
  INV_X1 U669 ( .A(G1956), .ZN(n939) );
  NOR2_X1 U670 ( .A1(n646), .A2(n939), .ZN(n602) );
  NOR2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n639) );
  INV_X1 U672 ( .A(G299), .ZN(n1004) );
  NOR2_X1 U673 ( .A1(n639), .A2(n1004), .ZN(n605) );
  XNOR2_X1 U674 ( .A(n605), .B(n604), .ZN(n643) );
  NAND2_X1 U675 ( .A1(n662), .A2(G1341), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(KEYINPUT88), .ZN(n618) );
  NAND2_X1 U677 ( .A1(G68), .A2(n792), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n791), .A2(G81), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT12), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT13), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G43), .A2(n795), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U684 ( .A1(n613), .A2(G56), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT14), .B(n614), .Z(n615) );
  NAND2_X1 U686 ( .A1(n618), .A2(n1011), .ZN(n621) );
  NAND2_X1 U687 ( .A1(n598), .A2(G1996), .ZN(n619) );
  XOR2_X1 U688 ( .A(KEYINPUT26), .B(n619), .Z(n620) );
  NAND2_X1 U689 ( .A1(G92), .A2(n791), .ZN(n623) );
  NAND2_X1 U690 ( .A1(G66), .A2(n613), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U692 ( .A(KEYINPUT74), .B(n624), .ZN(n628) );
  NAND2_X1 U693 ( .A1(G79), .A2(n792), .ZN(n626) );
  NAND2_X1 U694 ( .A1(G54), .A2(n795), .ZN(n625) );
  NAND2_X1 U695 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U697 ( .A(KEYINPUT15), .B(n629), .Z(n904) );
  NAND2_X1 U698 ( .A1(n636), .A2(n904), .ZN(n635) );
  NAND2_X1 U699 ( .A1(n646), .A2(G2067), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(KEYINPUT90), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n662), .A2(G1348), .ZN(n631) );
  XOR2_X1 U702 ( .A(KEYINPUT89), .B(n631), .Z(n632) );
  NAND2_X1 U703 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n638) );
  OR2_X1 U705 ( .A1(n904), .A2(n636), .ZN(n637) );
  NAND2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n639), .A2(n1004), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U709 ( .A1(n643), .A2(n642), .ZN(n645) );
  XNOR2_X1 U710 ( .A(n645), .B(n644), .ZN(n650) );
  INV_X1 U711 ( .A(G1961), .ZN(n952) );
  NAND2_X1 U712 ( .A1(n952), .A2(n662), .ZN(n648) );
  XNOR2_X1 U713 ( .A(G2078), .B(KEYINPUT25), .ZN(n924) );
  NAND2_X1 U714 ( .A1(n646), .A2(n924), .ZN(n647) );
  NAND2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n654) );
  NAND2_X1 U716 ( .A1(G171), .A2(n654), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n659) );
  NAND2_X1 U718 ( .A1(G8), .A2(n662), .ZN(n753) );
  NOR2_X1 U719 ( .A1(G1966), .A2(n753), .ZN(n674) );
  NOR2_X1 U720 ( .A1(G2084), .A2(n662), .ZN(n671) );
  NOR2_X1 U721 ( .A1(n674), .A2(n671), .ZN(n651) );
  NAND2_X1 U722 ( .A1(G8), .A2(n651), .ZN(n652) );
  XNOR2_X1 U723 ( .A(KEYINPUT30), .B(n652), .ZN(n653) );
  NOR2_X1 U724 ( .A1(G168), .A2(n653), .ZN(n656) );
  NOR2_X1 U725 ( .A1(G171), .A2(n654), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT31), .B(n657), .Z(n658) );
  NAND2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n672) );
  NAND2_X1 U729 ( .A1(n672), .A2(G286), .ZN(n661) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n753), .ZN(n664) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n662), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U733 ( .A1(n665), .A2(G303), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U735 ( .A(KEYINPUT92), .B(n668), .ZN(n669) );
  NAND2_X1 U736 ( .A1(n669), .A2(G8), .ZN(n670) );
  XNOR2_X1 U737 ( .A(KEYINPUT32), .B(n670), .ZN(n746) );
  NAND2_X1 U738 ( .A1(G8), .A2(n671), .ZN(n676) );
  INV_X1 U739 ( .A(n672), .ZN(n673) );
  NOR2_X1 U740 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n747) );
  NAND2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n1009) );
  INV_X1 U743 ( .A(n753), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n1009), .A2(n677), .ZN(n681) );
  INV_X1 U745 ( .A(n681), .ZN(n678) );
  AND2_X1 U746 ( .A1(n747), .A2(n678), .ZN(n679) );
  NOR2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n687), .A2(n680), .ZN(n1000) );
  OR2_X1 U750 ( .A1(n681), .A2(n1000), .ZN(n683) );
  INV_X1 U751 ( .A(KEYINPUT33), .ZN(n682) );
  NAND2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n686), .B(KEYINPUT93), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n687), .A2(KEYINPUT33), .ZN(n688) );
  OR2_X1 U755 ( .A1(n753), .A2(n688), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n691), .B(KEYINPUT94), .ZN(n743) );
  XOR2_X1 U757 ( .A(G1981), .B(G305), .Z(n1001) );
  NAND2_X1 U758 ( .A1(G117), .A2(n881), .ZN(n694) );
  NAND2_X1 U759 ( .A1(G129), .A2(n692), .ZN(n693) );
  NAND2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U761 ( .A1(n579), .A2(G105), .ZN(n695) );
  XOR2_X1 U762 ( .A(KEYINPUT38), .B(n695), .Z(n696) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n701) );
  NAND2_X1 U764 ( .A1(n699), .A2(G141), .ZN(n700) );
  NAND2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n891) );
  NAND2_X1 U766 ( .A1(G1996), .A2(n891), .ZN(n709) );
  NAND2_X1 U767 ( .A1(G95), .A2(n579), .ZN(n703) );
  NAND2_X1 U768 ( .A1(G107), .A2(n881), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U770 ( .A1(G131), .A2(n699), .ZN(n705) );
  NAND2_X1 U771 ( .A1(G119), .A2(n692), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  OR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n890) );
  NAND2_X1 U774 ( .A1(G1991), .A2(n890), .ZN(n708) );
  NAND2_X1 U775 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U776 ( .A(KEYINPUT84), .B(n710), .ZN(n988) );
  NAND2_X1 U777 ( .A1(G40), .A2(G160), .ZN(n711) );
  NOR2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n739) );
  NAND2_X1 U779 ( .A1(n988), .A2(n739), .ZN(n713) );
  XOR2_X1 U780 ( .A(KEYINPUT85), .B(n713), .Z(n726) );
  NAND2_X1 U781 ( .A1(n579), .A2(G104), .ZN(n714) );
  XNOR2_X1 U782 ( .A(n714), .B(KEYINPUT82), .ZN(n716) );
  NAND2_X1 U783 ( .A1(G140), .A2(n699), .ZN(n715) );
  NAND2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n718) );
  XOR2_X1 U785 ( .A(KEYINPUT83), .B(KEYINPUT34), .Z(n717) );
  XNOR2_X1 U786 ( .A(n718), .B(n717), .ZN(n723) );
  NAND2_X1 U787 ( .A1(G116), .A2(n881), .ZN(n720) );
  NAND2_X1 U788 ( .A1(G128), .A2(n692), .ZN(n719) );
  NAND2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U790 ( .A(KEYINPUT35), .B(n721), .Z(n722) );
  NOR2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U792 ( .A(KEYINPUT36), .B(n724), .ZN(n901) );
  XNOR2_X1 U793 ( .A(G2067), .B(KEYINPUT37), .ZN(n735) );
  NOR2_X1 U794 ( .A1(n901), .A2(n735), .ZN(n981) );
  NAND2_X1 U795 ( .A1(n739), .A2(n981), .ZN(n733) );
  NAND2_X1 U796 ( .A1(n726), .A2(n733), .ZN(n725) );
  XOR2_X1 U797 ( .A(n725), .B(KEYINPUT86), .Z(n757) );
  AND2_X1 U798 ( .A1(n1001), .A2(n757), .ZN(n741) );
  NOR2_X1 U799 ( .A1(G1996), .A2(n891), .ZN(n973) );
  INV_X1 U800 ( .A(n726), .ZN(n729) );
  NOR2_X1 U801 ( .A1(G1986), .A2(G290), .ZN(n727) );
  NOR2_X1 U802 ( .A1(G1991), .A2(n890), .ZN(n978) );
  NOR2_X1 U803 ( .A1(n727), .A2(n978), .ZN(n728) );
  NOR2_X1 U804 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U805 ( .A(n730), .B(KEYINPUT96), .ZN(n731) );
  NOR2_X1 U806 ( .A1(n973), .A2(n731), .ZN(n732) );
  XNOR2_X1 U807 ( .A(n732), .B(KEYINPUT39), .ZN(n734) );
  NAND2_X1 U808 ( .A1(n734), .A2(n733), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n901), .A2(n735), .ZN(n986) );
  NAND2_X1 U810 ( .A1(n736), .A2(n986), .ZN(n737) );
  NAND2_X1 U811 ( .A1(n739), .A2(n737), .ZN(n738) );
  XNOR2_X1 U812 ( .A(KEYINPUT97), .B(n738), .ZN(n758) );
  XNOR2_X1 U813 ( .A(G1986), .B(G290), .ZN(n998) );
  NAND2_X1 U814 ( .A1(n739), .A2(n998), .ZN(n740) );
  OR2_X1 U815 ( .A1(n758), .A2(n740), .ZN(n761) );
  AND2_X1 U816 ( .A1(n741), .A2(n761), .ZN(n742) );
  NAND2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n763) );
  NOR2_X1 U818 ( .A1(G2090), .A2(G303), .ZN(n744) );
  XOR2_X1 U819 ( .A(KEYINPUT95), .B(n744), .Z(n745) );
  NAND2_X1 U820 ( .A1(G8), .A2(n745), .ZN(n749) );
  NAND2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n750), .A2(n753), .ZN(n755) );
  NOR2_X1 U824 ( .A1(G1981), .A2(G305), .ZN(n751) );
  XOR2_X1 U825 ( .A(n751), .B(KEYINPUT24), .Z(n752) );
  OR2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  AND2_X1 U828 ( .A1(n757), .A2(n756), .ZN(n759) );
  OR2_X1 U829 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U830 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U831 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U832 ( .A(n765), .B(n764), .ZN(G329) );
  INV_X1 U833 ( .A(G57), .ZN(G237) );
  INV_X1 U834 ( .A(G132), .ZN(G219) );
  INV_X1 U835 ( .A(G82), .ZN(G220) );
  NAND2_X1 U836 ( .A1(G94), .A2(G452), .ZN(n766) );
  XNOR2_X1 U837 ( .A(n766), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U839 ( .A(n767), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U840 ( .A(G223), .ZN(n826) );
  NAND2_X1 U841 ( .A1(n826), .A2(G567), .ZN(n768) );
  XNOR2_X1 U842 ( .A(n768), .B(KEYINPUT71), .ZN(n769) );
  XNOR2_X1 U843 ( .A(KEYINPUT11), .B(n769), .ZN(G234) );
  NAND2_X1 U844 ( .A1(G860), .A2(n1011), .ZN(G153) );
  XNOR2_X1 U845 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U846 ( .A1(G868), .A2(G301), .ZN(n771) );
  INV_X1 U847 ( .A(n904), .ZN(n996) );
  INV_X1 U848 ( .A(G868), .ZN(n811) );
  NAND2_X1 U849 ( .A1(n996), .A2(n811), .ZN(n770) );
  NAND2_X1 U850 ( .A1(n771), .A2(n770), .ZN(G284) );
  XNOR2_X1 U851 ( .A(KEYINPUT77), .B(G868), .ZN(n772) );
  NOR2_X1 U852 ( .A1(G286), .A2(n772), .ZN(n774) );
  NOR2_X1 U853 ( .A1(G868), .A2(G299), .ZN(n773) );
  NOR2_X1 U854 ( .A1(n774), .A2(n773), .ZN(G297) );
  INV_X1 U855 ( .A(G860), .ZN(n775) );
  NAND2_X1 U856 ( .A1(n775), .A2(G559), .ZN(n776) );
  NAND2_X1 U857 ( .A1(n776), .A2(n904), .ZN(n777) );
  XNOR2_X1 U858 ( .A(n777), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U859 ( .A1(n904), .A2(G868), .ZN(n778) );
  NOR2_X1 U860 ( .A1(G559), .A2(n778), .ZN(n780) );
  AND2_X1 U861 ( .A1(n1011), .A2(n811), .ZN(n779) );
  NOR2_X1 U862 ( .A1(n780), .A2(n779), .ZN(G282) );
  NAND2_X1 U863 ( .A1(G99), .A2(n579), .ZN(n782) );
  NAND2_X1 U864 ( .A1(G111), .A2(n881), .ZN(n781) );
  NAND2_X1 U865 ( .A1(n782), .A2(n781), .ZN(n788) );
  NAND2_X1 U866 ( .A1(G123), .A2(n692), .ZN(n783) );
  XNOR2_X1 U867 ( .A(n783), .B(KEYINPUT78), .ZN(n784) );
  XNOR2_X1 U868 ( .A(n784), .B(KEYINPUT18), .ZN(n786) );
  NAND2_X1 U869 ( .A1(G135), .A2(n699), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U871 ( .A1(n788), .A2(n787), .ZN(n977) );
  XNOR2_X1 U872 ( .A(n977), .B(G2096), .ZN(n790) );
  INV_X1 U873 ( .A(G2100), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(G156) );
  NAND2_X1 U875 ( .A1(G93), .A2(n791), .ZN(n794) );
  NAND2_X1 U876 ( .A1(G80), .A2(n792), .ZN(n793) );
  NAND2_X1 U877 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U878 ( .A1(G55), .A2(n795), .ZN(n796) );
  XNOR2_X1 U879 ( .A(KEYINPUT79), .B(n796), .ZN(n797) );
  NOR2_X1 U880 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U881 ( .A1(n613), .A2(G67), .ZN(n799) );
  NAND2_X1 U882 ( .A1(n800), .A2(n799), .ZN(n810) );
  NAND2_X1 U883 ( .A1(G559), .A2(n904), .ZN(n801) );
  XOR2_X1 U884 ( .A(n1011), .B(n801), .Z(n808) );
  NOR2_X1 U885 ( .A1(n808), .A2(G860), .ZN(n802) );
  XOR2_X1 U886 ( .A(n810), .B(n802), .Z(G145) );
  XNOR2_X1 U887 ( .A(KEYINPUT19), .B(G303), .ZN(n803) );
  XNOR2_X1 U888 ( .A(n803), .B(n810), .ZN(n804) );
  XNOR2_X1 U889 ( .A(n804), .B(G288), .ZN(n805) );
  XNOR2_X1 U890 ( .A(n805), .B(G290), .ZN(n806) );
  XNOR2_X1 U891 ( .A(n1004), .B(n806), .ZN(n807) );
  XNOR2_X1 U892 ( .A(n807), .B(G305), .ZN(n908) );
  XNOR2_X1 U893 ( .A(n908), .B(n808), .ZN(n809) );
  NAND2_X1 U894 ( .A1(n809), .A2(G868), .ZN(n813) );
  NAND2_X1 U895 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U896 ( .A1(n813), .A2(n812), .ZN(G295) );
  NAND2_X1 U897 ( .A1(G2078), .A2(G2084), .ZN(n814) );
  XOR2_X1 U898 ( .A(KEYINPUT20), .B(n814), .Z(n815) );
  NAND2_X1 U899 ( .A1(G2090), .A2(n815), .ZN(n816) );
  XNOR2_X1 U900 ( .A(KEYINPUT21), .B(n816), .ZN(n817) );
  NAND2_X1 U901 ( .A1(n817), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U903 ( .A1(G220), .A2(G219), .ZN(n818) );
  XOR2_X1 U904 ( .A(KEYINPUT22), .B(n818), .Z(n819) );
  NOR2_X1 U905 ( .A1(G218), .A2(n819), .ZN(n820) );
  NAND2_X1 U906 ( .A1(G96), .A2(n820), .ZN(n832) );
  NAND2_X1 U907 ( .A1(n832), .A2(G2106), .ZN(n824) );
  NAND2_X1 U908 ( .A1(G120), .A2(G69), .ZN(n821) );
  NOR2_X1 U909 ( .A1(G237), .A2(n821), .ZN(n822) );
  NAND2_X1 U910 ( .A1(G108), .A2(n822), .ZN(n833) );
  NAND2_X1 U911 ( .A1(n833), .A2(G567), .ZN(n823) );
  NAND2_X1 U912 ( .A1(n824), .A2(n823), .ZN(n846) );
  NAND2_X1 U913 ( .A1(G661), .A2(G483), .ZN(n825) );
  NOR2_X1 U914 ( .A1(n846), .A2(n825), .ZN(n830) );
  NAND2_X1 U915 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n826), .ZN(G217) );
  NAND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n827) );
  XNOR2_X1 U918 ( .A(KEYINPUT103), .B(n827), .ZN(n828) );
  NAND2_X1 U919 ( .A1(n828), .A2(G661), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT104), .B(n829), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(G188) );
  XNOR2_X1 U923 ( .A(G69), .B(KEYINPUT105), .ZN(G235) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  NOR2_X1 U927 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U929 ( .A(G2443), .B(G2438), .ZN(n843) );
  XOR2_X1 U930 ( .A(G2454), .B(G2430), .Z(n835) );
  XNOR2_X1 U931 ( .A(G2446), .B(KEYINPUT99), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U933 ( .A(G2451), .B(G2427), .Z(n837) );
  XNOR2_X1 U934 ( .A(G1341), .B(G1348), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U936 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U937 ( .A(KEYINPUT100), .B(G2435), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n844), .A2(G14), .ZN(n845) );
  XNOR2_X1 U941 ( .A(KEYINPUT101), .B(n845), .ZN(n915) );
  XNOR2_X1 U942 ( .A(n915), .B(KEYINPUT102), .ZN(G401) );
  INV_X1 U943 ( .A(n846), .ZN(G319) );
  XNOR2_X1 U944 ( .A(G1996), .B(G2474), .ZN(n856) );
  XOR2_X1 U945 ( .A(G1991), .B(G1986), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1961), .B(G1956), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U948 ( .A(G1976), .B(G1981), .Z(n850) );
  XNOR2_X1 U949 ( .A(G1966), .B(G1971), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U951 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U952 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U955 ( .A(G2100), .B(G2096), .Z(n858) );
  XNOR2_X1 U956 ( .A(KEYINPUT42), .B(G2678), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U958 ( .A(KEYINPUT43), .B(G2090), .Z(n860) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U962 ( .A(G2078), .B(G2084), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(G227) );
  NAND2_X1 U964 ( .A1(G136), .A2(n699), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G112), .A2(n881), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G124), .A2(n692), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n867), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G100), .A2(n579), .ZN(n868) );
  XOR2_X1 U970 ( .A(KEYINPUT107), .B(n868), .Z(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U972 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G115), .A2(n881), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G127), .A2(n692), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n875), .B(KEYINPUT47), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G139), .A2(n699), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G103), .A2(n579), .ZN(n878) );
  XNOR2_X1 U980 ( .A(KEYINPUT109), .B(n878), .ZN(n879) );
  NOR2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n967) );
  NAND2_X1 U982 ( .A1(G118), .A2(n881), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G130), .A2(n692), .ZN(n882) );
  NAND2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U985 ( .A1(G106), .A2(n579), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G142), .A2(n699), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U988 ( .A(KEYINPUT45), .B(n886), .Z(n887) );
  NOR2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n967), .B(n889), .ZN(n900) );
  XNOR2_X1 U991 ( .A(G164), .B(n890), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U993 ( .A(n893), .B(KEYINPUT48), .Z(n895) );
  XNOR2_X1 U994 ( .A(KEYINPUT108), .B(KEYINPUT46), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n977), .B(n896), .ZN(n898) );
  XNOR2_X1 U997 ( .A(G160), .B(G162), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n902), .B(n901), .Z(n903) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n903), .ZN(G395) );
  XOR2_X1 U1002 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n906) );
  XNOR2_X1 U1003 ( .A(G171), .B(n904), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n907), .B(G286), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n910), .B(n1011), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n911), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n912) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n912), .Z(n913) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n913), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1017 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1030) );
  XNOR2_X1 U1018 ( .A(KEYINPUT55), .B(KEYINPUT115), .ZN(n994) );
  XOR2_X1 U1019 ( .A(G2090), .B(G35), .Z(n920) );
  XOR2_X1 U1020 ( .A(G34), .B(KEYINPUT54), .Z(n918) );
  XNOR2_X1 U1021 ( .A(n918), .B(G2084), .ZN(n919) );
  NAND2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n934) );
  XOR2_X1 U1023 ( .A(G1991), .B(G25), .Z(n921) );
  NAND2_X1 U1024 ( .A1(n921), .A2(G28), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(G1996), .B(G32), .ZN(n923) );
  XNOR2_X1 U1026 ( .A(G33), .B(G2072), .ZN(n922) );
  NOR2_X1 U1027 ( .A1(n923), .A2(n922), .ZN(n928) );
  XOR2_X1 U1028 ( .A(n924), .B(G27), .Z(n926) );
  XNOR2_X1 U1029 ( .A(G2067), .B(G26), .ZN(n925) );
  NOR2_X1 U1030 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1033 ( .A(KEYINPUT116), .B(n931), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(KEYINPUT53), .B(n932), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1036 ( .A(n994), .B(n935), .Z(n936) );
  XNOR2_X1 U1037 ( .A(KEYINPUT117), .B(n936), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(G29), .A2(n937), .ZN(n1028) );
  XNOR2_X1 U1039 ( .A(G1348), .B(KEYINPUT59), .ZN(n938) );
  XNOR2_X1 U1040 ( .A(n938), .B(G4), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(KEYINPUT120), .B(G20), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(n940), .B(n939), .ZN(n941) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(G6), .B(G1981), .ZN(n943) );
  NOR2_X1 U1046 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1047 ( .A(n945), .B(KEYINPUT121), .ZN(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1049 ( .A(KEYINPUT60), .B(n948), .Z(n950) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(KEYINPUT122), .B(n951), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(n952), .B(G5), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n964) );
  XOR2_X1 U1055 ( .A(G1986), .B(G24), .Z(n960) );
  XOR2_X1 U1056 ( .A(G1976), .B(G23), .Z(n955) );
  XNOR2_X1 U1057 ( .A(KEYINPUT123), .B(n955), .ZN(n957) );
  XNOR2_X1 U1058 ( .A(G22), .B(G1971), .ZN(n956) );
  NOR2_X1 U1059 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1060 ( .A(n958), .B(KEYINPUT124), .ZN(n959) );
  NAND2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1062 ( .A(KEYINPUT58), .B(n961), .Z(n962) );
  XNOR2_X1 U1063 ( .A(KEYINPUT125), .B(n962), .ZN(n963) );
  NOR2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1065 ( .A(KEYINPUT61), .B(n965), .Z(n966) );
  NOR2_X1 U1066 ( .A1(G16), .A2(n966), .ZN(n1025) );
  XNOR2_X1 U1067 ( .A(G2072), .B(n967), .ZN(n969) );
  XNOR2_X1 U1068 ( .A(G164), .B(G2078), .ZN(n968) );
  NAND2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1070 ( .A(n970), .B(KEYINPUT50), .ZN(n971) );
  XNOR2_X1 U1071 ( .A(n971), .B(KEYINPUT113), .ZN(n976) );
  XOR2_X1 U1072 ( .A(G2090), .B(G162), .Z(n972) );
  NOR2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1074 ( .A(KEYINPUT51), .B(n974), .Z(n975) );
  NAND2_X1 U1075 ( .A1(n976), .A2(n975), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(G2084), .B(G160), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n982) );
  NOR2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1080 ( .A(KEYINPUT112), .B(n983), .Z(n984) );
  NOR2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n990) );
  INV_X1 U1082 ( .A(n986), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(KEYINPUT52), .B(n991), .ZN(n992) );
  XOR2_X1 U1086 ( .A(KEYINPUT114), .B(n992), .Z(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n995), .A2(G29), .ZN(n1023) );
  XNOR2_X1 U1089 ( .A(KEYINPUT56), .B(G16), .ZN(n1021) );
  XNOR2_X1 U1090 ( .A(G1348), .B(n996), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1018) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G168), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(n1003), .B(KEYINPUT57), .ZN(n1016) );
  XNOR2_X1 U1096 ( .A(n1004), .B(G1956), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(G1971), .A2(G303), .ZN(n1005) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(G171), .B(G1961), .Z(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(G1341), .B(n1011), .Z(n1012) );
  XNOR2_X1 U1103 ( .A(KEYINPUT118), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT119), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(G11), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(n1030), .B(n1029), .ZN(G311) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

