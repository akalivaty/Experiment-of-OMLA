//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G250), .ZN(new_n203));
  INV_X1    g0003(.A(G1), .ZN(new_n204));
  INV_X1    g0004(.A(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n203), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n205), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT64), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n223), .B1(new_n216), .B2(new_n224), .C1(new_n225), .C2(new_n203), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n211), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n207), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n222), .A2(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(new_n204), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G50), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n213), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(new_n204), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n256), .B1(new_n260), .B2(new_n255), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n215), .A2(KEYINPUT8), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G58), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT68), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n205), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G50), .A2(G58), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n205), .B1(new_n270), .B2(new_n216), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n205), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n271), .B1(new_n276), .B2(G150), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n269), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n261), .B1(new_n278), .B2(new_n258), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT9), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G223), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n284), .B1(new_n228), .B2(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(new_n289), .A3(G274), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n204), .B1(G41), .B2(G45), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n296), .B1(G226), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n291), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(G200), .B2(new_n301), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n281), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n279), .B1(new_n307), .B2(new_n301), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT70), .B(G179), .Z(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n310), .B2(new_n301), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT7), .B1(new_n316), .B2(new_n205), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT7), .ZN(new_n318));
  AOI211_X1 g0118(.A(new_n318), .B(G20), .C1(new_n313), .C2(new_n315), .ZN(new_n319));
  OAI21_X1  g0119(.A(G68), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G58), .A2(G68), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n217), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G20), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT73), .ZN(new_n324));
  INV_X1    g0124(.A(new_n276), .ZN(new_n325));
  INV_X1    g0125(.A(G159), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n274), .B2(new_n275), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n205), .B1(new_n217), .B2(new_n321), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT73), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n320), .A2(KEYINPUT16), .A3(new_n327), .A4(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT16), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n318), .B1(new_n282), .B2(G20), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n316), .A2(KEYINPUT7), .A3(new_n205), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n216), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n328), .A2(new_n329), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n331), .A2(new_n337), .A3(new_n258), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n266), .A2(new_n260), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n254), .B2(new_n266), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT74), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n289), .A2(G232), .A3(new_n297), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n295), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G87), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT75), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n313), .A2(new_n315), .A3(G226), .A4(G1698), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n313), .A2(new_n315), .A3(G223), .A4(new_n283), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n346), .B1(new_n352), .B2(new_n290), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n309), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT76), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n354), .B(new_n355), .C1(G169), .C2(new_n353), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(KEYINPUT76), .A3(new_n309), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n343), .A2(new_n344), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT18), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT18), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n343), .A2(new_n361), .A3(new_n344), .A4(new_n358), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT77), .B(G190), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n363), .B(new_n346), .C1(new_n290), .C2(new_n352), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n352), .A2(new_n290), .ZN(new_n366));
  INV_X1    g0166(.A(new_n346), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(new_n338), .A3(new_n340), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT17), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n360), .A2(new_n362), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n282), .A2(G232), .A3(G1698), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G97), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n313), .A2(new_n315), .A3(G226), .A4(new_n283), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n290), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT13), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n289), .A2(G274), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n299), .A2(G238), .B1(new_n379), .B2(new_n294), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n377), .B2(new_n380), .ZN(new_n382));
  OAI21_X1  g0182(.A(G169), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n377), .A2(new_n380), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT72), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT71), .B(KEYINPUT13), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n386), .ZN(new_n389));
  NAND2_X1  g0189(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n377), .A2(KEYINPUT72), .A3(new_n380), .A4(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n387), .A2(new_n389), .A3(G179), .A4(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT14), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n393), .B(G169), .C1(new_n381), .C2(new_n382), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n384), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n258), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n276), .A2(G50), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n268), .A2(G77), .B1(G20), .B2(new_n216), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n399), .A2(KEYINPUT11), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(KEYINPUT11), .ZN(new_n401));
  OR3_X1    g0201(.A1(new_n253), .A2(KEYINPUT12), .A3(G68), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT12), .B1(new_n253), .B2(G68), .ZN(new_n403));
  AOI22_X1  g0203(.A1(G68), .A2(new_n259), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n395), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n385), .A2(KEYINPUT13), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n388), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n408), .B2(G200), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n387), .A2(new_n389), .A3(G190), .A4(new_n391), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n265), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n325), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n415), .A2(new_n267), .B1(new_n205), .B2(new_n228), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n258), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n253), .A2(G77), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n259), .B2(G77), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n295), .B1(new_n229), .B2(new_n298), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n282), .A2(G232), .A3(new_n283), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n422), .B1(new_n230), .B2(new_n282), .C1(new_n285), .C2(new_n224), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n421), .B1(new_n423), .B2(new_n290), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n420), .B1(new_n424), .B2(G190), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n365), .B2(new_n424), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n309), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n420), .B1(new_n424), .B2(G169), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n312), .A2(new_n372), .A3(new_n412), .A4(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT82), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n203), .A2(new_n283), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n210), .A2(G1698), .ZN(new_n434));
  AND4_X1   g0234(.A1(new_n313), .A2(new_n433), .A3(new_n315), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G294), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT81), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G294), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n273), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n432), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n313), .A2(new_n433), .A3(new_n315), .A4(new_n434), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT81), .B(G294), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n442), .B(KEYINPUT82), .C1(new_n273), .C2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n290), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n204), .A2(G45), .ZN(new_n446));
  OR2_X1    g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  NAND2_X1  g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n449), .A2(new_n290), .A3(new_n211), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n379), .A2(new_n449), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n445), .A2(new_n302), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n433), .A2(new_n434), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n455), .A2(new_n316), .B1(new_n443), .B2(new_n273), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n289), .B1(new_n456), .B2(new_n432), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n450), .B1(new_n457), .B2(new_n444), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT83), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n302), .A4(new_n452), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n445), .A2(new_n452), .A3(new_n451), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n365), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n454), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n313), .A2(new_n315), .A3(new_n205), .A4(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT22), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT22), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n282), .A2(new_n466), .A3(new_n205), .A4(G87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G116), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G20), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT23), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n205), .B2(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n230), .A2(KEYINPUT23), .A3(G20), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT24), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT24), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n468), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n396), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n253), .B1(G1), .B2(new_n273), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(new_n258), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n230), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT25), .B1(new_n254), .B2(new_n230), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n482), .A2(new_n230), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n463), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n293), .A2(G1), .ZN(new_n489));
  INV_X1    g0289(.A(new_n213), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n488), .A2(new_n489), .B1(new_n490), .B2(new_n288), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G257), .B1(new_n379), .B2(new_n449), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n313), .A2(new_n315), .A3(G250), .A4(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n313), .A2(new_n315), .A3(G244), .A4(new_n283), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n282), .A2(new_n498), .A3(G244), .A4(new_n283), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT79), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n290), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n497), .A2(new_n499), .ZN(new_n503));
  INV_X1    g0303(.A(new_n495), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n503), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n492), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n307), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n230), .A2(KEYINPUT6), .A3(G97), .ZN(new_n508));
  OR2_X1    g0308(.A1(new_n508), .A2(KEYINPUT78), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g0310(.A(G97), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n230), .ZN(new_n512));
  NOR2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n508), .A2(KEYINPUT78), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n517));
  OAI21_X1  g0317(.A(G107), .B1(new_n317), .B2(new_n319), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n396), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n254), .A2(new_n511), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n482), .B2(new_n511), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n309), .B(new_n492), .C1(new_n502), .C2(new_n505), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n507), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n519), .A2(new_n521), .ZN(new_n525));
  OAI211_X1 g0325(.A(G190), .B(new_n492), .C1(new_n502), .C2(new_n505), .ZN(new_n526));
  INV_X1    g0326(.A(new_n492), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n503), .A2(new_n504), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n289), .B1(new_n528), .B2(KEYINPUT79), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n500), .A2(new_n501), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n525), .B(new_n526), .C1(new_n531), .C2(new_n365), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n487), .A2(new_n524), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n461), .A2(new_n307), .ZN(new_n534));
  INV_X1    g0334(.A(G179), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n458), .A2(new_n535), .A3(new_n452), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n536), .C1(new_n479), .C2(new_n485), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n494), .B(new_n205), .C1(G33), .C2(new_n511), .ZN(new_n538));
  INV_X1    g0338(.A(G116), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G20), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n258), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT20), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n253), .A2(G116), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n481), .B2(G116), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n307), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n491), .A2(G270), .B1(new_n379), .B2(new_n449), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n314), .A2(G33), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n549));
  OAI21_X1  g0349(.A(G303), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n313), .A2(new_n315), .A3(G264), .A4(G1698), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n313), .A2(new_n315), .A3(G257), .A4(new_n283), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n290), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT80), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT80), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n547), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n546), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n547), .A2(new_n554), .A3(G179), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n543), .A2(new_n545), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n546), .A2(new_n556), .A3(KEYINPUT21), .A4(new_n558), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n537), .A2(new_n561), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n363), .ZN(new_n567));
  INV_X1    g0367(.A(new_n558), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n557), .B1(new_n547), .B2(new_n554), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n556), .A2(G200), .A3(new_n558), .ZN(new_n571));
  INV_X1    g0371(.A(new_n563), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n205), .B1(new_n374), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n513), .A2(new_n225), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n313), .A2(new_n315), .A3(new_n205), .A4(G68), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n574), .B1(new_n267), .B2(new_n511), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n258), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n415), .A2(new_n254), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n481), .A2(G87), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n289), .A2(G274), .A3(new_n489), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n289), .A2(G250), .A3(new_n446), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n313), .A2(new_n315), .A3(G244), .A4(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n313), .A2(new_n315), .A3(G238), .A4(new_n283), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(new_n469), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n587), .B1(new_n290), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G190), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n584), .B(new_n592), .C1(new_n365), .C2(new_n591), .ZN(new_n593));
  INV_X1    g0393(.A(new_n591), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n307), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n581), .B(new_n582), .C1(new_n415), .C2(new_n482), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(new_n309), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n573), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n533), .A2(new_n566), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n431), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g0401(.A(new_n601), .B(KEYINPUT84), .Z(G372));
  INV_X1    g0402(.A(new_n306), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n358), .A2(new_n361), .A3(new_n341), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n361), .B1(new_n358), .B2(new_n341), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT87), .B1(new_n428), .B2(new_n429), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n423), .A2(new_n290), .ZN(new_n609));
  INV_X1    g0409(.A(new_n421), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n307), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT87), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n420), .A4(new_n427), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n411), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n406), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n607), .B1(new_n616), .B2(new_n371), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n311), .B1(new_n603), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n431), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n598), .A2(new_n593), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n524), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n524), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n584), .B(KEYINPUT85), .C1(new_n365), .C2(new_n591), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n590), .A2(new_n290), .ZN(new_n627));
  INV_X1    g0427(.A(new_n587), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n365), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n625), .A2(new_n592), .A3(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n632), .A2(KEYINPUT86), .A3(new_n598), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT86), .B1(new_n632), .B2(new_n598), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n624), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n623), .B1(new_n635), .B2(new_n621), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n566), .A2(new_n487), .A3(new_n524), .A4(new_n532), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n633), .A2(new_n634), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n598), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n619), .B1(new_n620), .B2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(new_n537), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n204), .A2(new_n205), .A3(G13), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT27), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n645), .A2(new_n204), .A3(new_n205), .A4(G13), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  OR3_X1    g0448(.A1(new_n647), .A2(KEYINPUT88), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT88), .B1(new_n647), .B2(new_n648), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n486), .A2(new_n652), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n486), .B2(new_n463), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(new_n655), .B2(new_n642), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n563), .A2(new_n651), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n573), .A2(new_n658), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n657), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT89), .Z(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT90), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT90), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n665), .A3(G330), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n656), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n655), .A2(new_n657), .A3(new_n537), .A4(new_n652), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n653), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n667), .A2(new_n669), .ZN(G399));
  NOR2_X1   g0470(.A1(new_n209), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n576), .A2(G116), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n218), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n524), .A2(KEYINPUT26), .A3(new_n622), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n631), .A2(new_n592), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n629), .A2(new_n630), .A3(new_n626), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n598), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT86), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n632), .A2(KEYINPUT86), .A3(new_n598), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n524), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n678), .B1(new_n685), .B2(new_n621), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n652), .B1(new_n639), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n687), .A2(KEYINPUT92), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT92), .ZN(new_n690));
  INV_X1    g0490(.A(new_n598), .ZN(new_n691));
  INV_X1    g0491(.A(new_n566), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n533), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n683), .A2(new_n684), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n677), .B1(new_n635), .B2(KEYINPUT26), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n651), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n690), .B1(new_n697), .B2(KEYINPUT29), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n688), .B1(new_n640), .B2(new_n651), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n689), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n562), .A2(new_n458), .A3(new_n591), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n506), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n445), .A2(new_n451), .A3(new_n591), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n547), .A2(new_n554), .A3(G179), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n531), .A2(new_n708), .A3(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n506), .A2(KEYINPUT91), .A3(new_n461), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT91), .B1(new_n506), .B2(new_n461), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n556), .A2(new_n309), .A3(new_n558), .A4(new_n594), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n710), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n702), .B1(new_n716), .B2(new_n652), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT31), .B(new_n651), .C1(new_n718), .C2(new_n710), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n566), .A2(new_n599), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n487), .A2(new_n524), .A3(new_n532), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(new_n652), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n701), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n676), .B1(new_n726), .B2(G1), .ZN(G364));
  NAND2_X1  g0527(.A1(new_n664), .A2(new_n666), .ZN(new_n728));
  INV_X1    g0528(.A(G13), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n204), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n671), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n662), .A2(G330), .ZN(new_n734));
  OR3_X1    g0534(.A1(new_n728), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n205), .A2(G190), .A3(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n310), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n205), .A2(G179), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(G190), .A3(G200), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n738), .A2(G311), .B1(new_n741), .B2(G303), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n309), .A2(new_n205), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n363), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G322), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n736), .A2(new_n535), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n739), .A2(new_n302), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G329), .A2(new_n749), .B1(new_n751), .B2(G283), .ZN(new_n752));
  INV_X1    g0552(.A(new_n443), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n535), .A2(new_n365), .A3(G190), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n282), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n742), .A2(new_n747), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n743), .A2(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(KEYINPUT96), .A3(new_n302), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT96), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n758), .B2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT33), .B(G317), .Z(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n758), .A2(new_n363), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n757), .B(new_n766), .C1(G326), .C2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT95), .B(G159), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n748), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n316), .B1(new_n751), .B2(G107), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n771), .B(new_n772), .C1(new_n215), .C2(new_n745), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n738), .A2(G77), .B1(new_n741), .B2(G87), .ZN(new_n774));
  INV_X1    g0574(.A(new_n755), .ZN(new_n775));
  INV_X1    g0575(.A(new_n767), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n774), .B1(new_n511), .B2(new_n775), .C1(new_n776), .C2(new_n255), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n773), .B(new_n777), .C1(G68), .C2(new_n763), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n768), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n213), .B1(G20), .B2(new_n307), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT94), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n733), .B(KEYINPUT93), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n208), .A2(new_n282), .ZN(new_n783));
  INV_X1    g0583(.A(G355), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n783), .A2(new_n784), .B1(G116), .B2(new_n208), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n248), .A2(G45), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n209), .A2(new_n282), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n293), .B2(new_n219), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n785), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n780), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n782), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n793), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n797), .B1(new_n781), .B2(new_n796), .C1(new_n662), .C2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n735), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n420), .A2(new_n651), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n608), .B2(new_n614), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT99), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n428), .B2(new_n429), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n612), .A2(KEYINPUT99), .A3(new_n420), .A4(new_n427), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n805), .A2(new_n426), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n803), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n792), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n780), .A2(new_n791), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n782), .B1(G77), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT97), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n769), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n746), .A2(G143), .B1(new_n738), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  INV_X1    g0617(.A(G150), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n816), .B1(new_n817), .B2(new_n776), .C1(new_n764), .C2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT34), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n751), .A2(G68), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n255), .B2(new_n740), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT98), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n316), .B1(new_n755), .B2(G58), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n748), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n764), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G303), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n776), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n738), .A2(G116), .B1(new_n751), .B2(G87), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n230), .B2(new_n740), .C1(new_n832), .C2(new_n748), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n316), .B1(new_n511), .B2(new_n775), .C1(new_n745), .C2(new_n436), .ZN(new_n834));
  OR3_X1    g0634(.A1(new_n830), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n820), .A2(new_n826), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n809), .B(new_n814), .C1(new_n836), .C2(new_n780), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n807), .A2(new_n802), .ZN(new_n838));
  INV_X1    g0638(.A(new_n803), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n640), .B2(new_n651), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n807), .A2(new_n651), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n636), .B2(new_n639), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(new_n724), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n733), .B1(new_n844), .B2(new_n724), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n837), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  NOR2_X1   g0649(.A1(new_n730), .A2(new_n204), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT40), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n327), .A2(new_n330), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n332), .B1(new_n852), .B2(new_n335), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n258), .A3(new_n331), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n647), .B1(new_n854), .B2(new_n340), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n372), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n340), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n356), .A2(new_n357), .A3(new_n647), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n369), .A2(new_n338), .A3(new_n340), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n343), .A2(new_n344), .A3(new_n858), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n370), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n856), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n856), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n395), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n411), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n401), .A2(new_n404), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n399), .A2(KEYINPUT11), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n651), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(KEYINPUT100), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT100), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n405), .A2(new_n878), .A3(new_n651), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n406), .A2(new_n411), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n840), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n723), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n851), .B1(new_n869), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n856), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n884));
  INV_X1    g0684(.A(new_n647), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n343), .A2(new_n344), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n606), .B2(new_n371), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n356), .A2(new_n357), .B1(new_n338), .B2(new_n340), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n860), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n863), .B1(new_n889), .B2(new_n886), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT101), .B1(new_n862), .B2(new_n864), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n862), .A2(KEYINPUT101), .A3(new_n864), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n884), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n877), .A2(new_n879), .ZN(new_n896));
  AOI221_X4 g0696(.A(new_n896), .B1(new_n410), .B2(new_n409), .C1(new_n395), .C2(new_n405), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n874), .B1(new_n870), .B2(new_n411), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n808), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n651), .B1(new_n718), .B2(new_n710), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n600), .A2(new_n652), .B1(new_n900), .B2(new_n702), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n901), .B2(new_n719), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n895), .A2(KEYINPUT40), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n883), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT102), .Z(new_n905));
  NAND2_X1  g0705(.A1(new_n431), .A2(new_n723), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(G330), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n619), .B1(new_n700), .B2(new_n620), .ZN(new_n910));
  INV_X1    g0710(.A(new_n869), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n897), .A2(new_n898), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n805), .A2(new_n806), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n652), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n843), .B2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n911), .A2(new_n915), .B1(new_n607), .B2(new_n647), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n895), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n406), .A2(new_n651), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n856), .A2(new_n866), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT38), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(KEYINPUT39), .A3(new_n884), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n918), .A2(new_n919), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n910), .B(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n850), .B1(new_n909), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n909), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(G116), .A3(new_n214), .A4(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n219), .A2(G77), .A3(new_n321), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(G50), .B2(new_n216), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(G1), .A3(new_n729), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n928), .A2(new_n932), .A3(new_n935), .ZN(G367));
  NAND2_X1  g0736(.A1(new_n651), .A2(new_n630), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n694), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT103), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n598), .A2(new_n937), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(KEYINPUT103), .B2(new_n938), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n793), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n243), .A2(new_n788), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n794), .B1(new_n208), .B2(new_n415), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n782), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n738), .A2(G283), .B1(G107), .B2(new_n755), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n511), .B2(new_n750), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n767), .B2(G311), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT46), .B1(new_n741), .B2(G116), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n741), .A2(KEYINPUT46), .A3(G116), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n749), .A2(G317), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(new_n316), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n950), .B(new_n953), .C1(G303), .C2(new_n746), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n949), .B(new_n954), .C1(new_n443), .C2(new_n764), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n282), .B1(new_n228), .B2(new_n750), .C1(new_n745), .C2(new_n818), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n737), .A2(new_n255), .B1(new_n216), .B2(new_n775), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n748), .A2(new_n817), .B1(new_n740), .B2(new_n215), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n767), .A2(G143), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n764), .C2(new_n769), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n955), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT47), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n946), .B1(new_n963), .B2(new_n780), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n943), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n657), .A2(new_n652), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n656), .B(new_n966), .Z(new_n967));
  AND3_X1   g0767(.A1(new_n664), .A2(KEYINPUT106), .A3(new_n666), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT106), .B1(new_n664), .B2(new_n666), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n967), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n656), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n728), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n624), .A2(new_n651), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n524), .B(new_n532), .C1(new_n525), .C2(new_n652), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n669), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n669), .A2(new_n977), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n974), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n667), .A2(new_n983), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n726), .B1(new_n972), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n671), .B(KEYINPUT41), .Z(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n732), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n977), .A2(new_n668), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT42), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n977), .B(KEYINPUT105), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n624), .B1(new_n994), .B2(new_n642), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n993), .B1(new_n995), .B2(new_n651), .ZN(new_n996));
  XNOR2_X1  g0796(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n942), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n996), .B(new_n998), .C1(new_n999), .C2(new_n942), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n996), .B2(new_n998), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n667), .A2(new_n994), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n965), .B1(new_n991), .B2(new_n1003), .ZN(G387));
  INV_X1    g0804(.A(new_n726), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n972), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n970), .A2(new_n726), .A3(new_n971), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n671), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n780), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n746), .A2(G317), .B1(new_n738), .B2(G303), .ZN(new_n1010));
  INV_X1    g0810(.A(G322), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n776), .C1(new_n764), .C2(new_n832), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT48), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n741), .A2(new_n753), .B1(new_n755), .B2(G283), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT49), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n316), .B1(new_n750), .B2(new_n539), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G326), .B2(new_n749), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n767), .A2(G159), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT107), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n763), .A2(new_n266), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n282), .B1(new_n511), .B2(new_n750), .C1(new_n745), .C2(new_n255), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n775), .A2(new_n415), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n818), .B2(new_n748), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n737), .A2(new_n216), .B1(new_n228), .B2(new_n740), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1025), .A2(new_n1026), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1009), .B1(new_n1023), .B2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n783), .A2(new_n673), .B1(G107), .B2(new_n208), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n239), .A2(new_n293), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n673), .ZN(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n1036), .C1(G68), .C2(G77), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n265), .A2(new_n255), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT50), .Z(new_n1039));
  AOI21_X1  g0839(.A(new_n788), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1034), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n782), .B1(new_n1041), .B2(new_n795), .ZN(new_n1042));
  OR3_X1    g0842(.A1(new_n1033), .A2(KEYINPUT108), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(KEYINPUT108), .B1(new_n1033), .B2(new_n1042), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n656), .A2(new_n793), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n969), .A2(new_n967), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT106), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n728), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n664), .A2(KEYINPUT106), .A3(new_n666), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1047), .B1(new_n1051), .B2(new_n967), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1046), .B1(new_n1052), .B2(new_n732), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1008), .A2(new_n1053), .ZN(G393));
  NAND2_X1  g0854(.A1(new_n1007), .A2(new_n987), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n671), .B1(new_n1007), .B2(new_n987), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n985), .A2(new_n986), .A3(new_n732), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT111), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n782), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n767), .A2(G317), .B1(new_n746), .B2(G311), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  OAI22_X1  g0862(.A1(new_n748), .A2(new_n1011), .B1(new_n740), .B2(new_n827), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(KEYINPUT109), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n737), .A2(new_n436), .B1(new_n539), .B2(new_n775), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1063), .A2(KEYINPUT109), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n316), .B1(new_n750), .B2(new_n230), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1062), .B(new_n1068), .C1(new_n829), .C2(new_n764), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n767), .A2(G150), .B1(new_n746), .B2(G159), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT51), .Z(new_n1071));
  AOI22_X1  g0871(.A1(new_n749), .A2(G143), .B1(G77), .B2(new_n755), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n216), .B2(new_n740), .C1(new_n413), .C2(new_n737), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n316), .B(new_n1073), .C1(G87), .C2(new_n751), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1071), .B(new_n1074), .C1(new_n255), .C2(new_n764), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1009), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n787), .A2(new_n251), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n795), .B1(G97), .B2(new_n209), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1060), .B(new_n1076), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT110), .Z(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n798), .B2(new_n994), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1058), .A2(new_n1059), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1059), .B1(new_n1058), .B2(new_n1081), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1056), .A2(new_n1057), .B1(new_n1083), .B2(new_n1084), .ZN(G390));
  OAI21_X1  g0885(.A(KEYINPUT112), .B1(new_n915), .B2(new_n919), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT112), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n919), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n914), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n721), .A2(new_n694), .A3(new_n566), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n685), .A2(KEYINPUT26), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n598), .C1(new_n1091), .C2(new_n623), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1089), .B1(new_n1092), .B2(new_n842), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1087), .B(new_n1088), .C1(new_n1093), .C2(new_n912), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n918), .A2(new_n923), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1086), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n912), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1097), .A2(new_n723), .A3(G330), .A4(new_n808), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1089), .B1(new_n697), .B2(new_n808), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1088), .B(new_n895), .C1(new_n1099), .C2(new_n912), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1098), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1095), .A2(new_n791), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n782), .B1(new_n266), .B2(new_n811), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT114), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n763), .A2(G107), .B1(G97), .B2(new_n738), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1107), .A2(KEYINPUT117), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(KEYINPUT117), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n821), .B1(new_n436), .B2(new_n748), .C1(new_n228), .C2(new_n775), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n316), .B1(new_n225), .B2(new_n740), .C1(new_n745), .C2(new_n539), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(G283), .C2(new_n767), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n316), .B1(new_n755), .B2(G159), .ZN(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1114), .B1(new_n255), .B2(new_n750), .C1(new_n1115), .C2(new_n748), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n818), .B2(new_n740), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n741), .A2(G150), .A3(new_n1117), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(new_n745), .C2(new_n825), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1116), .B(new_n1121), .C1(G128), .C2(new_n767), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n763), .A2(G137), .B1(new_n738), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT115), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1122), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1125), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1128), .A2(KEYINPUT115), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1113), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1106), .B1(new_n1130), .B2(new_n780), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1103), .A2(new_n732), .B1(new_n1104), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n431), .A2(new_n725), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n619), .B(new_n1134), .C1(new_n700), .C2(new_n620), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n912), .B1(new_n724), .B2(new_n840), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1136), .A2(new_n1099), .A3(new_n1098), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1093), .B1(new_n1136), .B2(new_n1098), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1101), .A2(new_n1102), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1098), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1140), .A2(new_n1146), .A3(new_n671), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT113), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1140), .A2(new_n1146), .A3(KEYINPUT113), .A4(new_n671), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1133), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(G378));
  AOI21_X1  g0952(.A(new_n882), .B1(new_n884), .B2(new_n922), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n903), .B(G330), .C1(new_n1153), .C2(KEYINPUT40), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT122), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT122), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n883), .A2(new_n1156), .A3(G330), .A4(new_n903), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n279), .A2(new_n647), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT55), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n312), .B(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n312), .B(new_n1159), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1155), .A2(new_n1157), .A3(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n904), .A2(new_n1167), .A3(new_n1156), .A4(G330), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n925), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n925), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1169), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n732), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n733), .B1(G50), .B2(new_n811), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n764), .A2(new_n511), .B1(new_n415), .B2(new_n737), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT119), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n749), .A2(G283), .B1(G68), .B2(new_n755), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n215), .B2(new_n750), .C1(new_n745), .C2(new_n230), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n292), .B(new_n316), .C1(new_n740), .C2(new_n228), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n776), .A2(new_n539), .B1(KEYINPUT118), .B2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(KEYINPUT118), .C2(new_n1181), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1178), .A2(KEYINPUT58), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G50), .B1(new_n273), .B2(new_n292), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n282), .B2(G41), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n738), .A2(G137), .B1(G150), .B2(new_n755), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n740), .B2(new_n1123), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G128), .B2(new_n746), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n1115), .B2(new_n776), .C1(new_n764), .C2(new_n825), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n751), .A2(new_n815), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G33), .B(G41), .C1(new_n749), .C2(G124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1184), .B(new_n1186), .C1(new_n1191), .C2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT58), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1176), .B1(new_n1198), .B2(new_n780), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1168), .B2(new_n792), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT121), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1175), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1172), .A2(KEYINPUT57), .A3(new_n1174), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1135), .B1(new_n1103), .B2(new_n1141), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n671), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1169), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1173), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1135), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1146), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT57), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1202), .B1(new_n1205), .B2(new_n1211), .ZN(G375));
  NOR2_X1   g1012(.A1(new_n1141), .A2(new_n989), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1139), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n282), .B1(new_n215), .B2(new_n750), .C1(new_n745), .C2(new_n817), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n738), .A2(G150), .B1(new_n749), .B2(G128), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n255), .B2(new_n775), .C1(new_n326), .C2(new_n740), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(G132), .C2(new_n767), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n763), .A2(new_n1124), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n316), .B1(new_n228), .B2(new_n750), .C1(new_n745), .C2(new_n827), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n738), .A2(G107), .B1(new_n749), .B2(G303), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n1028), .C1(new_n511), .C2(new_n740), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(G294), .C2(new_n767), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n763), .A2(G116), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1219), .A2(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n782), .B1(G68), .B2(new_n811), .C1(new_n1226), .C2(new_n1009), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n912), .B2(new_n791), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1214), .B2(new_n732), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1215), .A2(new_n1229), .ZN(G381));
  NAND3_X1  g1030(.A1(new_n1008), .A2(new_n800), .A3(new_n1053), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(G390), .A2(new_n1231), .A3(G381), .A4(G384), .ZN(new_n1232));
  INV_X1    g1032(.A(G387), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1175), .A2(new_n1201), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1206), .A2(new_n1207), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n672), .B1(new_n1236), .B2(new_n1210), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1235), .B1(new_n1238), .B2(new_n1204), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1234), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1147), .A2(new_n1132), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1232), .A2(new_n1233), .A3(new_n1240), .A4(new_n1241), .ZN(G407));
  INV_X1    g1042(.A(G213), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(G343), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1240), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT123), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(G213), .A3(G407), .ZN(G409));
  NOR3_X1   g1047(.A1(new_n1238), .A2(new_n1204), .A3(new_n989), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1175), .A2(new_n1200), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1241), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(G375), .B2(new_n1151), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1244), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1141), .A2(new_n672), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1135), .A2(new_n1139), .A3(KEYINPUT60), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(G384), .A3(new_n1229), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G384), .B1(new_n1257), .B2(new_n1229), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1251), .A2(new_n1252), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT62), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1251), .A2(new_n1265), .A3(new_n1252), .A4(new_n1261), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1244), .A2(G2897), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT124), .Z(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1260), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1268), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n1258), .A3(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1208), .A2(new_n990), .A3(new_n1210), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n1175), .A3(new_n1200), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1240), .A2(G378), .B1(new_n1241), .B2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1273), .B1(new_n1276), .B2(new_n1244), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .A4(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1057), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1084), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1280), .A2(new_n1055), .B1(new_n1281), .B2(new_n1082), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1008), .A2(new_n800), .A3(new_n1053), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n800), .B1(new_n1008), .B2(new_n1053), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(G387), .A2(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n987), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1005), .B1(new_n1286), .B2(new_n1052), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n731), .B1(new_n1287), .B2(new_n989), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1003), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G390), .B1(new_n1290), .B2(new_n965), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1279), .B1(new_n1285), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n965), .A3(G390), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1284), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1231), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G387), .A2(new_n1282), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1293), .A2(new_n1295), .A3(new_n1296), .A4(KEYINPUT126), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1292), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1295), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1290), .A2(KEYINPUT125), .A3(G390), .A4(new_n965), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1296), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT125), .B1(new_n1233), .B2(G390), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1299), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1298), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1278), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  OR2_X1    g1107(.A1(new_n1262), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1309), .B2(new_n1273), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1262), .A2(new_n1307), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1308), .A2(new_n1310), .A3(new_n1304), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1306), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(new_n1240), .A2(G378), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1261), .A2(KEYINPUT127), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G375), .A2(new_n1241), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1261), .A2(KEYINPUT127), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1298), .A2(new_n1303), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1298), .B2(new_n1303), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1317), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1304), .A2(new_n1318), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1317), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1298), .A2(new_n1303), .A3(new_n1319), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1323), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1322), .A2(new_n1326), .ZN(G402));
endmodule


