//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n646, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n456), .B1(new_n458), .B2(KEYINPUT67), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(KEYINPUT67), .B2(new_n458), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  INV_X1    g036(.A(KEYINPUT72), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(G2104), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR3_X1   g040(.A1(new_n465), .A2(KEYINPUT72), .A3(G2105), .ZN(new_n466));
  OAI21_X1  g041(.A(G101), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT69), .B(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT71), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n470), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n467), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(KEYINPUT70), .A2(G113), .A3(G2104), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n472), .A2(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n474), .A2(new_n482), .A3(G125), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n468), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n476), .A2(new_n484), .ZN(G160));
  NOR2_X1   g060(.A1(new_n475), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n475), .A2(new_n468), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT73), .Z(G162));
  NAND2_X1  g067(.A1(new_n463), .A2(KEYINPUT69), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT4), .A4(G138), .ZN(new_n496));
  NAND2_X1  g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n470), .A2(new_n473), .A3(new_n474), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n493), .A2(new_n495), .A3(G138), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n474), .A2(new_n482), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(new_n463), .B2(G114), .ZN(new_n505));
  NOR2_X1   g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT74), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(G102), .A2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(G114), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(G2104), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n500), .A2(new_n504), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  AND2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT75), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT75), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT6), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n518), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n520), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n527), .A2(new_n532), .A3(G62), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n521), .A2(new_n523), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G50), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n527), .A2(G75), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n529), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n534), .A2(new_n538), .ZN(G166));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n540), .B1(new_n516), .B2(new_n517), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n530), .A2(KEYINPUT76), .A3(new_n531), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n541), .A2(new_n542), .A3(G63), .A4(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT77), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT7), .Z(new_n546));
  INV_X1    g121(.A(KEYINPUT6), .ZN(new_n547));
  OR2_X1    g122(.A1(KEYINPUT75), .A2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(KEYINPUT75), .A2(G651), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n522), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n529), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n546), .B1(new_n552), .B2(G51), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n524), .A2(G89), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n544), .A2(new_n553), .A3(new_n554), .ZN(G168));
  AOI22_X1  g130(.A1(new_n552), .A2(G52), .B1(G90), .B2(new_n524), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n541), .A2(new_n542), .A3(G64), .ZN(new_n557));
  NAND2_X1  g132(.A1(G77), .A2(G543), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n526), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G171));
  NAND2_X1  g137(.A1(new_n552), .A2(G43), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n541), .A2(new_n542), .A3(G56), .ZN(new_n565));
  NAND2_X1  g140(.A1(G68), .A2(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n526), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n524), .A2(G81), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n563), .A2(new_n564), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n535), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G43), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT78), .B1(new_n573), .B2(new_n567), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G860), .ZN(G153));
  NAND4_X1  g152(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g153(.A1(G1), .A2(G3), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT8), .ZN(new_n580));
  NAND4_X1  g155(.A1(G319), .A2(G483), .A3(G661), .A4(new_n580), .ZN(G188));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n532), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G651), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(G65), .B1(new_n516), .B2(new_n517), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n588), .A2(KEYINPUT80), .A3(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g165(.A1(KEYINPUT79), .A2(G53), .ZN(new_n591));
  OAI211_X1 g166(.A(G543), .B(new_n591), .C1(new_n550), .C2(new_n522), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT9), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n592), .A2(new_n593), .B1(new_n524), .B2(G91), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n535), .A2(KEYINPUT9), .A3(G543), .A4(new_n591), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(G299));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n556), .B2(new_n560), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n524), .A2(G90), .ZN(new_n599));
  INV_X1    g174(.A(G52), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n571), .B2(new_n600), .ZN(new_n601));
  NOR3_X1   g176(.A1(new_n601), .A2(KEYINPUT81), .A3(new_n559), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n598), .A2(new_n602), .ZN(G301));
  NAND3_X1  g178(.A1(new_n544), .A2(new_n553), .A3(new_n554), .ZN(G286));
  INV_X1    g179(.A(G166), .ZN(G303));
  NAND3_X1  g180(.A1(new_n535), .A2(G87), .A3(new_n532), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n535), .A2(G49), .A3(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(G74), .B1(new_n541), .B2(new_n542), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(new_n584), .C2(new_n608), .ZN(G288));
  NAND2_X1  g184(.A1(G48), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT83), .B1(new_n551), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n535), .A2(new_n612), .A3(G48), .A4(G543), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n524), .A2(G86), .ZN(new_n614));
  INV_X1    g189(.A(G73), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT82), .B1(new_n615), .B2(new_n529), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n617), .A2(G73), .A3(G543), .ZN(new_n618));
  INV_X1    g193(.A(G61), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n618), .C1(new_n518), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n527), .ZN(new_n621));
  NAND4_X1  g196(.A1(new_n611), .A2(new_n613), .A3(new_n614), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT84), .ZN(G305));
  AOI22_X1  g198(.A1(new_n552), .A2(G47), .B1(G85), .B2(new_n524), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n541), .A2(new_n542), .A3(G60), .ZN(new_n625));
  INV_X1    g200(.A(G72), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n529), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n527), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(G290));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NOR2_X1   g205(.A1(G301), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n524), .A2(G92), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G79), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n635), .A2(new_n529), .A3(KEYINPUT85), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT85), .B1(new_n635), .B2(new_n529), .ZN(new_n637));
  INV_X1    g212(.A(G66), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n518), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n552), .A2(G54), .B1(G651), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT86), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n631), .B1(new_n643), .B2(new_n630), .ZN(G284));
  AOI21_X1  g219(.A(new_n631), .B1(new_n643), .B2(new_n630), .ZN(G321));
  NAND2_X1  g220(.A1(G299), .A2(new_n630), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(G168), .B2(new_n630), .ZN(G297));
  OAI21_X1  g222(.A(new_n646), .B1(G168), .B2(new_n630), .ZN(G280));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n643), .B1(new_n649), .B2(G860), .ZN(G148));
  NAND2_X1  g225(.A1(new_n643), .A2(new_n649), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n643), .A2(KEYINPUT87), .A3(new_n649), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(G868), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n576), .A2(new_n630), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT11), .Z(G282));
  INV_X1    g233(.A(new_n657), .ZN(G323));
  OR2_X1    g234(.A1(new_n464), .A2(new_n466), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT3), .B(G2104), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT13), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT89), .B(G2100), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT90), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n486), .A2(G135), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n488), .A2(G123), .ZN(new_n671));
  OAI221_X1 g246(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G2096), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(G2096), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n665), .A2(new_n667), .ZN(new_n676));
  NAND4_X1  g251(.A1(new_n669), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(G156));
  XNOR2_X1  g252(.A(G2427), .B(G2438), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2430), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT15), .B(G2435), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT14), .ZN(new_n683));
  XOR2_X1   g258(.A(G1341), .B(G1348), .Z(new_n684));
  XNOR2_X1  g259(.A(G2443), .B(G2446), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT91), .B(KEYINPUT16), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2451), .B(G2454), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G14), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(G401));
  XNOR2_X1  g269(.A(G2072), .B(G2078), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT17), .ZN(new_n696));
  XNOR2_X1  g271(.A(G2067), .B(G2678), .ZN(new_n697));
  XOR2_X1   g272(.A(G2084), .B(G2090), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT93), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n696), .A2(new_n697), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(new_n699), .C1(new_n695), .C2(new_n697), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n698), .A2(new_n695), .A3(new_n697), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n701), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G2096), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G2100), .ZN(G227));
  XOR2_X1   g284(.A(G1971), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT94), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT19), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1956), .B(G2474), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1961), .B(G1966), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n713), .A2(new_n714), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n712), .A2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n720));
  OAI221_X1 g295(.A(new_n716), .B1(new_n712), .B2(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  OR3_X1    g297(.A1(new_n721), .A2(G1986), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(G1986), .B1(new_n721), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(G1991), .B(G1996), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT96), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1981), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(G229));
  NOR2_X1   g309(.A1(G6), .A2(G16), .ZN(new_n735));
  INV_X1    g310(.A(G305), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT32), .B(G1981), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT99), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n737), .B(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT98), .B(G16), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(G22), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G166), .B2(new_n742), .ZN(new_n744));
  INV_X1    g319(.A(G1971), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G16), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G23), .ZN(new_n748));
  INV_X1    g323(.A(G288), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n747), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT33), .B(G1976), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT34), .B1(new_n740), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n742), .A2(G24), .ZN(new_n755));
  INV_X1    g330(.A(G290), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n742), .ZN(new_n757));
  INV_X1    g332(.A(G1986), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT97), .B(G29), .Z(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G25), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n486), .A2(G131), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n488), .A2(G119), .ZN(new_n764));
  OAI221_X1 g339(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(new_n761), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT35), .B(G1991), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n754), .A2(new_n759), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n740), .A2(KEYINPUT34), .A3(new_n753), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n747), .A2(G4), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n643), .B2(new_n747), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1348), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n760), .A2(G26), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT28), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n488), .A2(G128), .ZN(new_n781));
  OAI221_X1 g356(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n468), .C2(G116), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G140), .B2(new_n486), .ZN(new_n784));
  INV_X1    g359(.A(G29), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2067), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n742), .A2(G19), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n576), .B2(new_n742), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1341), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n778), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT100), .ZN(new_n792));
  NOR2_X1   g367(.A1(G286), .A2(new_n747), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT102), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G16), .B2(G21), .ZN(new_n795));
  INV_X1    g370(.A(G1966), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT103), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n795), .A2(new_n796), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n785), .A2(G33), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT25), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n486), .A2(G139), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n661), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n802), .B(new_n803), .C1(new_n468), .C2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n800), .B1(new_n805), .B2(G29), .ZN(new_n806));
  INV_X1    g381(.A(G2072), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT101), .ZN(new_n809));
  INV_X1    g384(.A(G28), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT30), .ZN(new_n811));
  AOI21_X1  g386(.A(G29), .B1(new_n810), .B2(KEYINPUT30), .ZN(new_n812));
  OR2_X1    g387(.A1(KEYINPUT31), .A2(G11), .ZN(new_n813));
  NAND2_X1  g388(.A1(KEYINPUT31), .A2(G11), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n811), .A2(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(G160), .A2(G29), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT24), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(G34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(G34), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n760), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G2084), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n815), .B1(new_n673), .B2(new_n760), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n747), .A2(G5), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G171), .B2(new_n747), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n823), .B1(G1961), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n806), .A2(new_n807), .B1(new_n822), .B2(new_n821), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n761), .A2(G27), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G164), .B2(new_n761), .ZN(new_n829));
  INV_X1    g404(.A(G2078), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n826), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  OR3_X1    g407(.A1(new_n799), .A2(new_n809), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(G162), .A2(new_n761), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G35), .B2(new_n761), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT29), .B(G2090), .Z(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT26), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n660), .A2(G105), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n486), .A2(G141), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n488), .A2(G129), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  MUX2_X1   g420(.A(G32), .B(new_n845), .S(G29), .Z(new_n846));
  XOR2_X1   g421(.A(KEYINPUT27), .B(G1996), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n825), .B2(G1961), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n846), .A2(new_n847), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n835), .A2(new_n836), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n741), .A2(G20), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT23), .ZN(new_n854));
  INV_X1    g429(.A(G299), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n747), .ZN(new_n856));
  INV_X1    g431(.A(G1956), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n837), .A2(new_n851), .A3(new_n852), .A4(new_n858), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n798), .A2(new_n833), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n775), .A2(new_n792), .A3(new_n860), .ZN(G150));
  INV_X1    g436(.A(G150), .ZN(G311));
  NAND2_X1  g437(.A1(new_n524), .A2(G93), .ZN(new_n863));
  INV_X1    g438(.A(G55), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n571), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n541), .A2(new_n542), .A3(G67), .ZN(new_n866));
  NAND2_X1  g441(.A1(G80), .A2(G543), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n526), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G860), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT37), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n869), .B1(new_n570), .B2(new_n574), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n573), .A2(new_n567), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n869), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT38), .Z(new_n880));
  AND2_X1   g455(.A1(new_n643), .A2(G559), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n880), .B(new_n881), .Z(new_n882));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n874), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n880), .B(new_n881), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(KEYINPUT104), .A3(KEYINPUT39), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G860), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n885), .B2(KEYINPUT39), .ZN(new_n889));
  OAI211_X1 g464(.A(KEYINPUT105), .B(new_n873), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n884), .B2(new_n886), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(new_n872), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(G145));
  XNOR2_X1  g469(.A(new_n784), .B(new_n514), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n805), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n766), .B(KEYINPUT107), .Z(new_n897));
  NAND2_X1  g472(.A1(new_n486), .A2(G142), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n488), .A2(G130), .ZN(new_n899));
  OAI221_X1 g474(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n897), .B(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n896), .B(new_n902), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n664), .B(new_n845), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n896), .B(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n904), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n673), .B(KEYINPUT106), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(G160), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(G162), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  INV_X1    g489(.A(new_n912), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n906), .A2(new_n915), .A3(new_n908), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g493(.A1(new_n642), .A2(G299), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n641), .A2(new_n855), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n653), .A2(new_n654), .A3(new_n879), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n879), .B1(new_n653), .B2(new_n654), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n919), .A2(KEYINPUT41), .A3(new_n920), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT41), .B1(new_n919), .B2(new_n920), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n924), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n736), .A2(G290), .ZN(new_n931));
  XNOR2_X1  g506(.A(G166), .B(new_n749), .ZN(new_n932));
  NAND2_X1  g507(.A1(G305), .A2(new_n756), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n930), .B1(new_n937), .B2(KEYINPUT42), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(KEYINPUT109), .A3(new_n939), .ZN(new_n940));
  OR3_X1    g515(.A1(new_n936), .A2(KEYINPUT108), .A3(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT108), .B1(new_n936), .B2(new_n939), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n938), .A2(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n929), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n929), .A2(new_n943), .ZN(new_n945));
  OAI21_X1  g520(.A(G868), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n870), .A2(new_n630), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(G295));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n947), .ZN(G331));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n575), .A2(new_n870), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT81), .B1(new_n601), .B2(new_n559), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n556), .A2(new_n597), .A3(new_n560), .ZN(new_n955));
  AOI21_X1  g530(.A(G286), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(G286), .A2(new_n561), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n953), .B(new_n877), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(G168), .B1(new_n598), .B2(new_n602), .ZN(new_n959));
  NAND2_X1  g534(.A1(G286), .A2(new_n561), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n959), .B(new_n960), .C1(new_n875), .C2(new_n878), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n963), .A3(new_n921), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n958), .B(new_n961), .C1(new_n926), .C2(new_n927), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n962), .B2(new_n921), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n952), .B1(new_n968), .B2(new_n937), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n936), .B1(new_n966), .B2(new_n967), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n970), .A2(new_n971), .A3(new_n914), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n970), .B2(new_n914), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n928), .A2(new_n962), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n962), .A2(new_n921), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n936), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n977), .A2(new_n914), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n968), .A2(new_n937), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n950), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n969), .A2(new_n978), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n979), .B1(new_n972), .B2(new_n973), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(new_n952), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n982), .B1(new_n950), .B2(new_n986), .ZN(G397));
  INV_X1    g562(.A(G2067), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n784), .B(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n989), .A2(new_n845), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n513), .A2(new_n504), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n475), .B1(new_n496), .B2(new_n497), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n468), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n474), .A2(new_n482), .A3(G125), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n479), .A2(new_n480), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n493), .A2(new_n495), .A3(G137), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n465), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n472), .A2(G2104), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1004), .A3(new_n470), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1000), .A2(new_n1005), .A3(G40), .A4(new_n467), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n996), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1007), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1009), .A2(G1996), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n990), .A2(new_n1007), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  XNOR2_X1  g588(.A(new_n845), .B(G1996), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n989), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n769), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1015), .A2(new_n766), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n988), .B2(new_n784), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1007), .A2(new_n758), .A3(new_n756), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT127), .Z(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT48), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n766), .B(new_n769), .Z(new_n1022));
  NOR2_X1   g597(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1009), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1020), .A2(KEYINPUT48), .ZN(new_n1025));
  OAI22_X1  g600(.A1(new_n1009), .A2(new_n1018), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1013), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(G8), .B(new_n1029), .C1(new_n534), .C2(new_n538), .ZN(new_n1030));
  INV_X1    g605(.A(G8), .ZN(new_n1031));
  INV_X1    g606(.A(new_n538), .ZN(new_n1032));
  INV_X1    g607(.A(new_n534), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(KEYINPUT113), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1030), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n1039));
  NOR2_X1   g614(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n992), .B2(new_n993), .ZN(new_n1041));
  INV_X1    g616(.A(G40), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n476), .A2(new_n484), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n468), .A2(new_n661), .A3(G138), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1044), .A2(new_n501), .B1(new_n507), .B2(new_n512), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1384), .B1(new_n1045), .B2(new_n500), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1041), .B(new_n1043), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G2090), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n995), .A2(G1384), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n992), .B2(new_n993), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1043), .B(new_n1052), .C1(new_n1046), .C2(KEYINPUT45), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1049), .A2(new_n1050), .B1(new_n1053), .B2(new_n745), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1038), .B(new_n1039), .C1(new_n1054), .C2(new_n1031), .ZN(new_n1055));
  INV_X1    g630(.A(G74), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n516), .A2(new_n517), .A3(new_n540), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT76), .B1(new_n530), .B2(new_n531), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G651), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1060), .A2(G1976), .A3(new_n606), .A4(new_n607), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1061), .B(G8), .C1(new_n994), .C2(new_n1006), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1046), .A2(new_n1043), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(G8), .A4(new_n1061), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n622), .A2(G1981), .ZN(new_n1069));
  AOI22_X1  g644(.A1(G86), .A2(new_n524), .B1(new_n620), .B2(new_n527), .ZN(new_n1070));
  INV_X1    g645(.A(G1981), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n611), .A4(new_n613), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1069), .A2(KEYINPUT49), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1066), .A2(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1068), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1052), .A2(new_n1043), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n514), .B2(new_n991), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n745), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1006), .B1(new_n514), .B2(new_n1040), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1050), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1031), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n1085), .B2(new_n1037), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(G8), .A3(new_n1037), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1055), .A2(new_n1078), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1077), .A2(new_n1073), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1068), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1088), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1094), .A2(KEYINPUT125), .A3(new_n1055), .A4(new_n1086), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1961), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1048), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1006), .B1(new_n514), .B2(new_n1051), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1099), .A2(new_n996), .A3(KEYINPUT53), .A4(new_n830), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT123), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1098), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1053), .B2(G2078), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1102), .A2(G301), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(G171), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT116), .B1(new_n1048), .B2(G2084), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1082), .A2(new_n1083), .A3(new_n1113), .A4(new_n822), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT115), .B1(new_n1116), .B2(G1966), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1053), .A2(new_n1118), .A3(new_n796), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1115), .A2(new_n1120), .A3(G168), .ZN(new_n1121));
  AOI21_X1  g696(.A(G168), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g697(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1123));
  OAI211_X1 g698(.A(G8), .B(new_n1121), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1119), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1118), .B1(new_n1053), .B2(new_n796), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1112), .B(new_n1114), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(G8), .B1(new_n1127), .B2(G286), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1111), .B1(new_n1124), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1048), .A2(new_n857), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1099), .A2(new_n996), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT80), .B1(new_n588), .B2(G651), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n582), .B(new_n584), .C1(new_n586), .C2(new_n587), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n595), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n592), .A2(new_n593), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n524), .A2(G91), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT117), .B(new_n1132), .C1(new_n1140), .C2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .A4(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1066), .A2(G2067), .ZN(new_n1146));
  AOI21_X1  g721(.A(G1348), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1145), .B(new_n642), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1136), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1053), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(G1956), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1144), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1150), .A2(new_n1151), .B1(new_n1152), .B2(new_n1133), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(KEYINPUT121), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n1156));
  OAI221_X1 g731(.A(new_n1156), .B1(new_n1152), .B2(new_n1133), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT61), .B1(new_n1158), .B2(new_n1145), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT58), .B(G1341), .Z(new_n1160));
  NAND2_X1  g735(.A1(new_n1066), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT119), .B(G1996), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1053), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n576), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1163), .B(new_n576), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1146), .ZN(new_n1171));
  INV_X1    g746(.A(G1348), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1048), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(KEYINPUT60), .A3(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1174), .A2(new_n642), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1145), .A2(new_n1153), .A3(KEYINPUT61), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(new_n1147), .B2(new_n1146), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1174), .A2(new_n1178), .A3(new_n642), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1170), .A2(new_n1175), .A3(new_n1176), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1154), .B1(new_n1159), .B2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1106), .A2(G301), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT124), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT53), .B1(new_n1116), .B2(new_n830), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(KEYINPUT123), .B2(new_n1101), .ZN(new_n1185));
  AOI21_X1  g760(.A(G301), .B1(new_n1185), .B2(new_n1104), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1108), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1096), .A2(new_n1131), .A3(new_n1181), .A4(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1078), .A2(new_n1085), .A3(new_n1037), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1072), .ZN(new_n1190));
  NOR2_X1   g765(.A1(G288), .A2(G1976), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1092), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1189), .B1(new_n1074), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1127), .A2(G8), .A3(G168), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1038), .B1(new_n1054), .B2(new_n1031), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1195), .A2(new_n1196), .A3(new_n1094), .A4(KEYINPUT63), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1089), .B2(new_n1194), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1193), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1188), .A2(KEYINPUT126), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT126), .B1(new_n1188), .B2(new_n1200), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(KEYINPUT62), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1124), .A2(new_n1130), .A3(new_n1205), .ZN(new_n1206));
  AND4_X1   g781(.A1(new_n1096), .A2(new_n1204), .A3(new_n1186), .A4(new_n1206), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1201), .A2(new_n1202), .A3(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(G290), .B(new_n758), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1009), .B1(new_n1023), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1027), .B1(new_n1208), .B2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g786(.A(new_n460), .B1(new_n692), .B2(new_n693), .ZN(new_n1213));
  OR2_X1    g787(.A1(G227), .A2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g788(.A1(G229), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n1215), .A2(new_n917), .ZN(new_n1216));
  NOR2_X1   g790(.A1(new_n1216), .A2(new_n986), .ZN(G308));
  NAND2_X1  g791(.A1(new_n985), .A2(new_n952), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1218), .A2(new_n983), .ZN(new_n1219));
  NAND3_X1  g793(.A1(new_n1219), .A2(new_n917), .A3(new_n1215), .ZN(G225));
endmodule


