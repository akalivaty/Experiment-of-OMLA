//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n209), .B1(new_n211), .B2(new_n212), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XNOR2_X1  g0032(.A(G50), .B(G58), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G351));
  INV_X1    g0041(.A(G50), .ZN(new_n242));
  INV_X1    g0042(.A(G58), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n242), .A2(new_n243), .A3(new_n214), .ZN(new_n244));
  NOR2_X1   g0044(.A1(G20), .A2(G33), .ZN(new_n245));
  AOI22_X1  g0045(.A1(new_n244), .A2(G20), .B1(G150), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT67), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n243), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n246), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G1), .A2(G13), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n259), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n257), .B1(new_n262), .B2(new_n263), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n242), .B1(new_n259), .B2(G20), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n265), .A2(new_n242), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n271), .B1(new_n210), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n210), .A2(new_n272), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n274), .ZN(new_n278));
  INV_X1    g0078(.A(G226), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(G222), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  INV_X1    g0086(.A(G223), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(G1698), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n285), .B1(new_n286), .B2(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n256), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n280), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n270), .A2(KEYINPUT9), .B1(G190), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n293), .B1(KEYINPUT9), .B2(new_n270), .C1(new_n294), .C2(new_n292), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n269), .B1(new_n292), .B2(G169), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G244), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n276), .B1(new_n278), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT3), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT3), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G107), .ZN(new_n310));
  OR2_X1    g0110(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n311));
  NAND2_X1  g0111(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n306), .A3(new_n308), .A4(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G232), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n310), .B1(new_n313), .B2(new_n314), .C1(new_n215), .C2(new_n288), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n304), .B1(new_n315), .B2(new_n291), .ZN(new_n316));
  INV_X1    g0116(.A(new_n245), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n247), .A2(new_n317), .B1(new_n252), .B2(new_n286), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n253), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n257), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n265), .A2(new_n286), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n259), .A2(G20), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n266), .A2(G77), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n316), .A2(G190), .B1(KEYINPUT69), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n315), .A2(new_n291), .ZN(new_n327));
  INV_X1    g0127(.A(new_n304), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G200), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n325), .A2(KEYINPUT69), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n326), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n316), .A2(new_n298), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n334), .B(new_n325), .C1(G169), .C2(new_n316), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n302), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n284), .B2(G20), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n309), .A2(KEYINPUT7), .A3(new_n252), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n214), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n243), .A2(new_n214), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G58), .A2(G68), .ZN(new_n344));
  OAI21_X1  g0144(.A(G20), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G159), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n317), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n338), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT72), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n257), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n340), .A2(new_n341), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(new_n352), .B2(G68), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(KEYINPUT16), .ZN(new_n354));
  OAI211_X1 g0154(.A(KEYINPUT72), .B(new_n338), .C1(new_n342), .C2(new_n347), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n350), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(G274), .B1(new_n290), .B2(new_n256), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n278), .A2(new_n314), .B1(new_n357), .B2(new_n274), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n284), .A2(G226), .A3(G1698), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G87), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n287), .C2(new_n313), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n358), .B1(new_n361), .B2(new_n291), .ZN(new_n362));
  INV_X1    g0162(.A(G190), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G200), .B2(new_n362), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n251), .B1(new_n259), .B2(G20), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n266), .B1(new_n265), .B2(new_n251), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n356), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT17), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n356), .A2(new_n365), .A3(KEYINPUT17), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT74), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n370), .A2(KEYINPUT74), .A3(new_n371), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n356), .A2(new_n367), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G169), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n362), .A2(new_n379), .ZN(new_n380));
  AOI211_X1 g0180(.A(new_n298), .B(new_n358), .C1(new_n361), .C2(new_n291), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT73), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n362), .A2(G179), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT73), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n384), .C1(new_n379), .C2(new_n362), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n378), .A2(new_n386), .A3(KEYINPUT18), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n382), .A2(new_n385), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(new_n377), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n376), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n394), .B1(new_n313), .B2(new_n279), .C1(new_n314), .C2(new_n288), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n291), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n276), .B1(new_n278), .B2(new_n215), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n393), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g0199(.A(KEYINPUT13), .B(new_n397), .C1(new_n395), .C2(new_n291), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT14), .B1(new_n401), .B2(new_n379), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(G169), .C1(new_n399), .C2(new_n400), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT71), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n401), .B2(G179), .ZN(new_n406));
  NOR4_X1   g0206(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT71), .A4(new_n298), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n402), .B(new_n404), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n253), .A2(new_n286), .B1(new_n252), .B2(G68), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT70), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n409), .A2(new_n410), .B1(new_n242), .B2(new_n317), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n409), .A2(new_n410), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n257), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT11), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n265), .A2(new_n214), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n414), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n266), .A2(G68), .A3(new_n323), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n415), .A2(new_n417), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n408), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n401), .B2(G190), .ZN(new_n422));
  OAI21_X1  g0222(.A(G200), .B1(new_n399), .B2(new_n400), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n337), .A2(new_n392), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT4), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n306), .A2(new_n308), .A3(G244), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n311), .A2(new_n312), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT4), .A4(G244), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G283), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT75), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT75), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(G33), .A3(G283), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n430), .A2(new_n431), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n291), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT5), .B(G41), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n259), .A2(G45), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT76), .B1(new_n443), .B2(new_n357), .ZN(new_n444));
  OR2_X1    g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT76), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n273), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n447), .A2(new_n291), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n444), .A2(new_n449), .B1(new_n450), .B2(G257), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n439), .A2(new_n298), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT77), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n439), .A2(new_n451), .A3(KEYINPUT77), .A4(new_n298), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n439), .A2(new_n451), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n264), .A2(G97), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n305), .A2(G1), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n265), .A2(new_n257), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n458), .B1(new_n460), .B2(G97), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n462), .A2(new_n202), .A3(G107), .ZN(new_n463));
  XNOR2_X1  g0263(.A(G97), .B(G107), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n465), .A2(new_n252), .B1(new_n286), .B2(new_n317), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n203), .B1(new_n340), .B2(new_n341), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n257), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n457), .A2(new_n379), .B1(new_n461), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n456), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n461), .A2(new_n468), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n457), .A2(G200), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n363), .C2(new_n457), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT19), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n253), .B2(new_n202), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT79), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT79), .B(new_n475), .C1(new_n253), .C2(new_n202), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n284), .A2(new_n252), .A3(G68), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n252), .B1(new_n394), .B2(new_n475), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(G87), .B2(new_n204), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n257), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n319), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n460), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n486), .B(new_n488), .C1(new_n264), .C2(new_n487), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n291), .A2(new_n442), .A3(new_n217), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n273), .B2(new_n442), .ZN(new_n491));
  INV_X1    g0291(.A(G1698), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n428), .A2(new_n492), .B1(new_n305), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT78), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n313), .B2(new_n215), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT78), .A4(G238), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n491), .B1(new_n498), .B2(new_n277), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n379), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n298), .B(new_n491), .C1(new_n498), .C2(new_n277), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n489), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n485), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n351), .B1(new_n503), .B2(new_n480), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n266), .B1(G1), .B2(new_n305), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n216), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n264), .A2(new_n487), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n499), .A2(G200), .ZN(new_n509));
  OAI211_X1 g0309(.A(G190), .B(new_n491), .C1(new_n498), .C2(new_n277), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n474), .A2(KEYINPUT80), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n470), .A2(new_n473), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(new_n512), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n443), .A2(G264), .A3(new_n277), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT84), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n450), .A2(new_n520), .A3(G264), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n444), .A2(new_n449), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n284), .A2(G257), .A3(G1698), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G294), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n525), .C1(new_n217), .C2(new_n313), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n291), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G179), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n519), .A2(new_n521), .B1(new_n526), .B2(new_n291), .ZN(new_n530));
  AOI21_X1  g0330(.A(G169), .B1(new_n530), .B2(new_n523), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n306), .A2(new_n308), .A3(new_n252), .A4(G87), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n533), .B(KEYINPUT22), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT24), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n203), .A3(G20), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT83), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n536), .B2(new_n203), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n537), .A2(KEYINPUT83), .B1(new_n540), .B2(G20), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n534), .A2(new_n535), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n535), .B1(new_n534), .B2(new_n542), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n257), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n264), .A2(G107), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT25), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n547), .A2(KEYINPUT25), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(new_n203), .B2(new_n505), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n532), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n443), .A2(G270), .A3(new_n277), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n443), .A2(KEYINPUT76), .A3(new_n357), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n448), .B1(new_n447), .B2(new_n273), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n283), .A2(new_n284), .A3(G257), .ZN(new_n559));
  AND2_X1   g0359(.A1(G264), .A2(G1698), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n306), .A2(new_n308), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G303), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n561), .B1(new_n284), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT81), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n283), .A2(new_n284), .A3(G257), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT81), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n309), .A2(G303), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n561), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n558), .B1(new_n569), .B2(new_n291), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n252), .B1(new_n202), .B2(G33), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n435), .B2(new_n433), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n257), .B1(new_n252), .B2(G116), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT20), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n571), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n436), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n255), .A2(new_n256), .B1(G20), .B2(new_n493), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT20), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n493), .B1(new_n264), .B2(new_n351), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n459), .A2(new_n493), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n262), .B2(new_n263), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n575), .A2(new_n579), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT21), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n379), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT82), .B1(new_n570), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n585), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n574), .B1(new_n572), .B2(new_n573), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n577), .A2(KEYINPUT20), .A3(new_n578), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n265), .A2(new_n581), .B1(new_n266), .B2(new_n493), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT82), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n277), .B1(new_n564), .B2(new_n568), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n558), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n587), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n379), .B1(new_n591), .B2(new_n592), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n595), .B2(new_n558), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n569), .A2(new_n291), .B1(new_n591), .B2(new_n592), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n558), .A2(new_n298), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n599), .A2(new_n584), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n554), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n528), .A2(new_n294), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n522), .A2(new_n363), .A3(new_n523), .A4(new_n527), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(KEYINPUT85), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n534), .A2(new_n542), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT24), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n543), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n551), .B1(new_n609), .B2(new_n257), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT85), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n530), .A2(new_n611), .A3(new_n363), .A4(new_n523), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n606), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n570), .A2(G190), .ZN(new_n614));
  INV_X1    g0414(.A(new_n583), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n614), .B(new_n615), .C1(new_n294), .C2(new_n570), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n603), .A2(new_n617), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n426), .A2(new_n514), .A3(new_n517), .A4(new_n618), .ZN(G372));
  INV_X1    g0419(.A(KEYINPUT89), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT88), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n456), .A2(new_n621), .A3(new_n469), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n456), .B2(new_n469), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n622), .A2(new_n623), .A3(new_n512), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n620), .B1(new_n624), .B2(KEYINPUT26), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n512), .A2(new_n470), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n470), .A2(KEYINPUT88), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n513), .ZN(new_n630));
  OAI211_X1 g0430(.A(KEYINPUT89), .B(new_n628), .C1(new_n630), .C2(new_n622), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n625), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n554), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n597), .A2(new_n602), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT86), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT86), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n597), .A2(new_n602), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n474), .A2(new_n513), .A3(new_n613), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n637), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n636), .B1(new_n597), .B2(new_n602), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n554), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n470), .A2(new_n513), .A3(new_n473), .A4(new_n613), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT87), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n632), .B(new_n502), .C1(new_n641), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n426), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n325), .B1(new_n316), .B2(G169), .ZN(new_n649));
  AOI211_X1 g0449(.A(G179), .B(new_n304), .C1(new_n315), .C2(new_n291), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n424), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n421), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n376), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n383), .B1(new_n379), .B2(new_n362), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n377), .A2(new_n388), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n388), .B1(new_n377), .B2(new_n655), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n300), .B1(new_n659), .B2(new_n296), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n648), .A2(new_n660), .ZN(G369));
  NAND3_X1  g0461(.A1(new_n259), .A2(new_n252), .A3(G13), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n615), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n635), .A2(new_n637), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT90), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n597), .A2(new_n602), .ZN(new_n672));
  INV_X1    g0472(.A(new_n669), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n616), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n671), .B1(new_n670), .B2(new_n674), .ZN(new_n677));
  OAI21_X1  g0477(.A(G330), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT91), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n642), .A2(new_n643), .A3(new_n673), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n672), .A2(new_n616), .A3(new_n673), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT90), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n675), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(KEYINPUT91), .A3(G330), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n554), .A2(new_n667), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n351), .B1(new_n608), .B2(new_n543), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n667), .B1(new_n689), .B2(new_n551), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n604), .A2(KEYINPUT85), .A3(new_n605), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n546), .A2(new_n552), .A3(new_n612), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n554), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n686), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n667), .B1(new_n597), .B2(new_n602), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n687), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n207), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n212), .B2(new_n703), .ZN(new_n706));
  XOR2_X1   g0506(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n707));
  XNOR2_X1  g0507(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n618), .A2(new_n514), .A3(new_n517), .A4(new_n668), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n457), .A2(new_n499), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n595), .A2(new_n298), .A3(new_n558), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(new_n530), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n570), .A2(G179), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(new_n457), .A3(new_n499), .A4(new_n528), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT30), .A4(new_n530), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n667), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(KEYINPUT31), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(KEYINPUT31), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n709), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n647), .A2(new_n668), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n645), .A2(new_n603), .ZN(new_n728));
  INV_X1    g0528(.A(new_n502), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n626), .B2(new_n628), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n728), .B(new_n730), .C1(new_n628), .C2(new_n624), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .A3(new_n668), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n724), .B1(new_n727), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n708), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(new_n684), .A2(G330), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT93), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G13), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n259), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n702), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n686), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n684), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n742), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n256), .B1(G20), .B2(new_n379), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n212), .A2(G45), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n309), .A2(new_n207), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT95), .ZN(new_n753));
  INV_X1    g0553(.A(G45), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n751), .B(new_n753), .C1(new_n236), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n701), .A2(new_n309), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n756), .A2(G355), .B1(new_n493), .B2(new_n701), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT94), .Z(new_n758));
  AOI211_X1 g0558(.A(new_n747), .B(new_n750), .C1(new_n755), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n252), .A2(G190), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G159), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT32), .ZN(new_n765));
  NAND3_X1  g0565(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n363), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(G50), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n252), .A2(G179), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(new_n363), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n203), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n298), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n760), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n772), .A2(G20), .A3(G190), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n284), .B1(new_n773), .B2(new_n286), .C1(new_n243), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n766), .A2(G190), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n771), .B(new_n775), .C1(G68), .C2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT96), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT96), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n216), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n252), .B1(new_n761), .B2(G190), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G97), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n768), .A2(new_n777), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n781), .A2(new_n562), .ZN(new_n788));
  INV_X1    g0588(.A(new_n784), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT33), .B(G317), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n789), .A2(G294), .B1(new_n776), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n770), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n792), .A2(G283), .B1(G326), .B2(new_n767), .ZN(new_n793));
  INV_X1    g0593(.A(new_n773), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n284), .B1(new_n794), .B2(G311), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n774), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G329), .B2(new_n763), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n791), .A2(new_n793), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n787), .B1(new_n788), .B2(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n749), .B(new_n759), .C1(new_n750), .C2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n737), .A2(new_n743), .B1(new_n748), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n325), .A2(new_n667), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n651), .B1(new_n333), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n335), .A2(new_n667), .ZN(new_n806));
  OAI21_X1  g0606(.A(KEYINPUT100), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT100), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n651), .A2(new_n668), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n331), .B1(G200), .B2(new_n329), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n810), .A2(new_n326), .B1(new_n325), .B2(new_n667), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n808), .B(new_n809), .C1(new_n811), .C2(new_n651), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n725), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT101), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n813), .A2(new_n667), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n640), .B1(new_n638), .B2(new_n639), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT87), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n729), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n817), .B1(new_n820), .B2(new_n632), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n815), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n742), .B1(new_n823), .B2(new_n723), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n723), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n750), .A2(new_n745), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT98), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n742), .B1(new_n827), .B2(G77), .ZN(new_n828));
  INV_X1    g0628(.A(new_n774), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(G143), .B1(new_n794), .B2(G159), .ZN(new_n830));
  INV_X1    g0630(.A(new_n776), .ZN(new_n831));
  INV_X1    g0631(.A(G150), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  INV_X1    g0633(.A(new_n767), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n830), .B1(new_n831), .B2(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT34), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  INV_X1    g0638(.A(new_n781), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G50), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n792), .A2(G68), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n841), .B(new_n284), .C1(new_n842), .C2(new_n762), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G58), .B2(new_n789), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n837), .A2(new_n838), .A3(new_n840), .A4(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G294), .ZN(new_n846));
  INV_X1    g0646(.A(G311), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n774), .A2(new_n846), .B1(new_n762), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n284), .B(new_n848), .C1(G116), .C2(new_n794), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n839), .A2(G107), .ZN(new_n850));
  XOR2_X1   g0650(.A(KEYINPUT99), .B(G283), .Z(new_n851));
  OAI22_X1  g0651(.A1(new_n831), .A2(new_n851), .B1(new_n834), .B2(new_n562), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n770), .A2(new_n216), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n849), .A2(new_n850), .A3(new_n786), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n845), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n828), .B1(new_n856), .B2(new_n750), .ZN(new_n857));
  INV_X1    g0657(.A(new_n813), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n746), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n825), .A2(new_n859), .ZN(G384));
  OAI21_X1  g0660(.A(G77), .B1(new_n243), .B2(new_n214), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n861), .A2(new_n212), .B1(G50), .B2(new_n214), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(G1), .A3(new_n738), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT102), .ZN(new_n864));
  INV_X1    g0664(.A(new_n465), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n493), .B(new_n211), .C1(new_n865), .C2(KEYINPUT35), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(KEYINPUT35), .B2(new_n865), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT36), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n354), .A2(new_n348), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n367), .ZN(new_n872));
  INV_X1    g0672(.A(new_n665), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n376), .B2(new_n391), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n872), .B1(new_n655), .B2(new_n873), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n877), .A2(new_n368), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n377), .A2(new_n873), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n881), .A2(new_n368), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT104), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT37), .B1(new_n389), .B2(new_n377), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n879), .B1(new_n378), .B2(new_n386), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n368), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT104), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n880), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT105), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n876), .A2(new_n890), .A3(new_n891), .A4(KEYINPUT38), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  INV_X1    g0693(.A(new_n372), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n881), .B1(new_n658), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n885), .A2(new_n888), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n377), .A2(new_n655), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT37), .B1(new_n887), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT105), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n875), .A2(new_n889), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n892), .B(new_n893), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n901), .B1(new_n875), .B2(new_n889), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(KEYINPUT39), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n421), .A2(new_n667), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n420), .A2(new_n667), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n421), .A2(new_n424), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n424), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n420), .B(new_n667), .C1(new_n913), .C2(new_n408), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n806), .B(KEYINPUT103), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n915), .B1(new_n821), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n904), .B2(new_n905), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n658), .A2(new_n873), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n910), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n727), .A2(new_n426), .A3(new_n732), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n921), .A2(new_n660), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n920), .B(new_n922), .Z(new_n923));
  AOI21_X1  g0723(.A(new_n813), .B1(new_n912), .B2(new_n914), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n722), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n904), .B2(new_n905), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n722), .A2(new_n924), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n928), .B(new_n892), .C1(new_n900), .C2(new_n902), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n927), .B1(new_n929), .B2(KEYINPUT40), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n426), .A2(new_n722), .ZN(new_n931));
  OAI21_X1  g0731(.A(G330), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n930), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n923), .A2(new_n933), .B1(new_n259), .B2(new_n739), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n923), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n870), .B1(new_n934), .B2(new_n935), .ZN(G367));
  NOR2_X1   g0736(.A1(new_n747), .A2(new_n750), .ZN(new_n937));
  INV_X1    g0737(.A(new_n753), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n937), .B1(new_n207), .B2(new_n319), .C1(new_n938), .C2(new_n231), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n742), .ZN(new_n940));
  INV_X1    g0740(.A(G143), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n834), .A2(new_n941), .B1(new_n770), .B2(new_n286), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n284), .B1(new_n773), .B2(new_n242), .C1(new_n832), .C2(new_n774), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n942), .B(new_n943), .C1(G159), .C2(new_n776), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n781), .A2(new_n243), .B1(new_n833), .B2(new_n762), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT109), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n785), .A2(G68), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n851), .A2(new_n773), .B1(new_n774), .B2(new_n562), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n284), .B(new_n951), .C1(G317), .C2(new_n763), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n839), .A2(KEYINPUT46), .A3(G116), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n792), .A2(G97), .B1(G311), .B2(new_n767), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n789), .A2(G107), .B1(G294), .B2(new_n776), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT46), .B1(new_n839), .B2(G116), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n949), .A2(new_n950), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n940), .B1(new_n959), .B2(new_n750), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n508), .A2(new_n668), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n513), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(new_n502), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n747), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n733), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n695), .B1(new_n672), .B2(new_n667), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n668), .B1(new_n546), .B2(new_n552), .ZN(new_n968));
  INV_X1    g0768(.A(new_n692), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(new_n969), .B2(new_n606), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n970), .A2(new_n634), .A3(new_n554), .A4(new_n668), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT91), .B1(new_n684), .B2(G330), .ZN(new_n974));
  INV_X1    g0774(.A(G330), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n679), .B(new_n975), .C1(new_n683), .C2(new_n675), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT106), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT106), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n680), .A2(new_n685), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n973), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n978), .B1(new_n680), .B2(new_n685), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n972), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n471), .A2(new_n668), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n470), .A2(new_n984), .A3(new_n473), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n470), .B2(new_n668), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n699), .A2(KEYINPUT45), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n971), .A2(new_n688), .ZN(new_n989));
  INV_X1    g0789(.A(new_n986), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(KEYINPUT44), .A3(new_n990), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n699), .B2(new_n986), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n987), .A2(new_n991), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n686), .A2(new_n696), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n996), .B1(new_n686), .B2(new_n696), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n966), .B1(new_n983), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n702), .B(KEYINPUT41), .Z(new_n1001));
  NOR3_X1   g0801(.A1(new_n1000), .A2(KEYINPUT107), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT107), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT106), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n972), .B1(new_n1004), .B2(new_n981), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n977), .A2(new_n973), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n697), .A2(new_n995), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n686), .A2(new_n696), .A3(new_n996), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n733), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1001), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1003), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n740), .B1(new_n1002), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n990), .A2(new_n971), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT42), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n633), .A2(new_n473), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n667), .B1(new_n1017), .B2(new_n470), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1015), .B2(KEYINPUT42), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n962), .A2(new_n963), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1016), .A2(new_n1019), .B1(KEYINPUT43), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n686), .A2(new_n696), .A3(new_n986), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT108), .B1(new_n1014), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(KEYINPUT107), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1011), .A2(new_n1003), .A3(new_n1012), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n741), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT108), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1025), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n965), .B1(new_n1026), .B2(new_n1032), .ZN(G387));
  NAND2_X1  g0833(.A1(new_n1007), .A2(new_n966), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n983), .A2(new_n733), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n1035), .A3(new_n702), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n704), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n756), .A2(new_n1037), .B1(new_n203), .B2(new_n701), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n228), .A2(new_n754), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n247), .A2(G50), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT50), .Z(new_n1041));
  OAI211_X1 g0841(.A(new_n704), .B(new_n754), .C1(new_n214), .C2(new_n286), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n753), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1038), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n749), .B1(new_n1044), .B2(new_n937), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n747), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n794), .A2(G68), .B1(new_n763), .B2(G150), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n792), .A2(G97), .B1(G159), .B2(new_n767), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n309), .B1(new_n829), .B2(G50), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n839), .A2(G77), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n785), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1051), .B1(new_n319), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n251), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1050), .B(new_n1053), .C1(new_n1054), .C2(new_n776), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n770), .A2(new_n493), .ZN(new_n1056));
  INV_X1    g0856(.A(G326), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n309), .B1(new_n762), .B2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n829), .A2(G317), .B1(new_n794), .B2(G303), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n831), .B2(new_n847), .C1(new_n796), .C2(new_n834), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n851), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n839), .A2(G294), .B1(new_n789), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1056), .B(new_n1058), .C1(new_n1067), .C2(KEYINPUT49), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1055), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n750), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1045), .B1(new_n696), .B2(new_n1046), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1036), .B(new_n1072), .C1(new_n740), .C2(new_n1007), .ZN(G393));
  INV_X1    g0873(.A(KEYINPUT110), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n740), .B1(new_n1010), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n1074), .B2(new_n1010), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n937), .B1(new_n202), .B2(new_n207), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n240), .B2(new_n753), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n749), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT111), .Z(new_n1080));
  AOI22_X1  g0880(.A1(new_n829), .A2(G311), .B1(G317), .B2(new_n767), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT52), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n839), .A2(new_n1064), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n309), .B1(new_n773), .B2(new_n846), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G322), .B2(new_n763), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n784), .A2(new_n493), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1086), .B(new_n771), .C1(G303), .C2(new_n776), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n284), .B1(new_n762), .B2(new_n941), .C1(new_n247), .C2(new_n773), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n853), .B(new_n1089), .C1(G50), .C2(new_n776), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n834), .A2(new_n832), .B1(new_n774), .B2(new_n346), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n785), .A2(G77), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n839), .A2(G68), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1088), .A2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1080), .B1(new_n1071), .B2(new_n1096), .C1(new_n986), .C2(new_n1046), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1076), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1035), .A2(new_n1010), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1035), .A2(new_n1010), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(new_n703), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1098), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(G390));
  NOR2_X1   g0903(.A1(new_n723), .A2(new_n813), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n915), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n903), .A2(new_n906), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n916), .B1(new_n647), .B2(new_n816), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n915), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n909), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT112), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(KEYINPUT112), .B(new_n909), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1107), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  MUX2_X1   g0914(.A(new_n900), .B(KEYINPUT105), .S(new_n902), .Z(new_n1115));
  NAND3_X1  g0915(.A1(new_n731), .A2(new_n668), .A3(new_n858), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n916), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n915), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n909), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1106), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1113), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT112), .B1(new_n917), .B2(new_n909), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n907), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(new_n1105), .A3(new_n1120), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n426), .A2(new_n724), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n921), .A2(new_n660), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT114), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n858), .B1(new_n724), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n723), .A2(KEYINPUT114), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1109), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1118), .B1(new_n1104), .B2(new_n915), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT113), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1109), .B1(new_n723), .B2(new_n813), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1105), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1108), .ZN(new_n1138));
  OAI211_X1 g0938(.A(KEYINPUT113), .B(new_n1109), .C1(new_n723), .C2(new_n813), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1128), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1122), .A2(new_n1126), .A3(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1142), .A2(new_n702), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT115), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1141), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(KEYINPUT115), .B(new_n1141), .C1(new_n1122), .C2(new_n1126), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1143), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1145), .A2(new_n740), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n907), .A2(new_n745), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n742), .B1(new_n827), .B2(new_n1054), .ZN(new_n1152));
  INV_X1    g0952(.A(G128), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1153), .A2(new_n834), .B1(new_n831), .B2(new_n833), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n829), .A2(G132), .B1(new_n794), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n309), .B1(new_n763), .B2(G125), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1154), .B(new_n1159), .C1(G50), .C2(new_n792), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n346), .B2(new_n1052), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n839), .A2(G150), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1093), .B1(new_n493), .B2(new_n774), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT116), .Z(new_n1165));
  INV_X1    g0965(.A(G283), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n841), .B1(new_n831), .B2(new_n203), .C1(new_n1166), .C2(new_n834), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n309), .B1(new_n762), .B2(new_n846), .C1(new_n202), .C2(new_n773), .ZN(new_n1168));
  OR3_X1    g0968(.A1(new_n782), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1161), .A2(new_n1163), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1152), .B1(new_n1170), .B2(new_n750), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1150), .B1(new_n1151), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1149), .A2(new_n1172), .ZN(G378));
  INV_X1    g0973(.A(KEYINPUT119), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n929), .A2(KEYINPUT40), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(G330), .C1(new_n1175), .C2(new_n927), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT119), .B1(new_n930), .B2(new_n975), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n269), .A2(new_n873), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n302), .B(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1179), .B(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1176), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1181), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(KEYINPUT119), .C1(new_n975), .C2(new_n930), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1182), .A2(new_n920), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n920), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n741), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1181), .A2(new_n745), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n750), .A2(G50), .A3(new_n745), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n284), .A2(G41), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(G33), .A2(G41), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1191), .A2(G50), .A3(new_n1192), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n774), .A2(KEYINPUT117), .A3(new_n203), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT117), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n829), .B2(G107), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(G58), .C2(new_n792), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1191), .B1(new_n1166), .B2(new_n762), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n831), .A2(new_n202), .B1(new_n834), .B2(new_n493), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n487), .C2(new_n794), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1200), .A3(new_n948), .A4(new_n1051), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT58), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1193), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT118), .ZN(new_n1204));
  INV_X1    g1004(.A(G124), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1192), .B1(new_n762), .B2(new_n1205), .C1(new_n346), .C2(new_n770), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n831), .A2(new_n842), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n774), .A2(new_n1153), .B1(new_n773), .B2(new_n833), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(G125), .C2(new_n767), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n832), .B2(new_n1052), .C1(new_n781), .C2(new_n1155), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1206), .B1(new_n1210), .B2(KEYINPUT59), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(KEYINPUT59), .B2(new_n1210), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1204), .B(new_n1212), .C1(new_n1202), .C2(new_n1201), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n749), .B(new_n1190), .C1(new_n1213), .C2(new_n750), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1189), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1188), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1128), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1142), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT120), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT120), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1142), .A2(new_n1220), .A3(new_n1217), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1185), .A2(new_n1186), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n703), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1142), .A2(new_n1220), .A3(new_n1217), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1220), .B1(new_n1142), .B2(new_n1217), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1187), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1223), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1216), .B1(new_n1225), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(G375));
  NAND2_X1  g1031(.A1(new_n1134), .A2(new_n1140), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1109), .A2(new_n745), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n742), .B1(new_n827), .B2(G68), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n839), .A2(G97), .B1(new_n487), .B2(new_n785), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n773), .A2(new_n203), .B1(new_n762), .B2(new_n562), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n284), .B(new_n1236), .C1(G283), .C2(new_n829), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n834), .A2(new_n846), .B1(new_n770), .B2(new_n286), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G116), .B2(new_n776), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n794), .A2(G150), .B1(new_n763), .B2(G128), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n833), .B2(new_n774), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n767), .A2(G132), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT121), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1242), .B(new_n1244), .C1(new_n776), .C2(new_n1156), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n242), .B2(new_n1052), .C1(new_n346), .C2(new_n781), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n284), .B1(new_n770), .B2(new_n243), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT122), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1240), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1234), .B1(new_n1249), .B2(new_n750), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1232), .A2(new_n741), .B1(new_n1233), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1146), .A2(new_n1012), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1232), .A2(new_n1217), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(G381));
  INV_X1    g1054(.A(G384), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1102), .A2(new_n1255), .ZN(new_n1256));
  OR2_X1    g1056(.A1(G393), .A2(G396), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(G378), .A2(G381), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1014), .A2(KEYINPUT108), .A3(new_n1025), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1030), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1258), .A2(new_n1230), .A3(new_n1261), .A4(new_n965), .ZN(G407));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n666), .A2(G213), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT123), .Z(new_n1265));
  NAND3_X1  g1065(.A1(new_n1230), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(G407), .A2(G213), .A3(new_n1266), .ZN(G409));
  XNOR2_X1  g1067(.A(G393), .B(new_n802), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G390), .B1(new_n1261), .B2(new_n965), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n965), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1271), .B(new_n1102), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1269), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(new_n1102), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1261), .A2(new_n965), .A3(G390), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1268), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1277), .B(KEYINPUT127), .Z(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1188), .A2(new_n1215), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1187), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1224), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n702), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G378), .B(new_n1280), .C1(new_n1281), .C2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1012), .B(new_n1187), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1263), .B1(new_n1286), .B2(new_n1216), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1265), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1265), .A2(G2897), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1134), .A2(new_n1140), .A3(new_n1128), .A4(KEYINPUT60), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1291), .A2(new_n702), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1141), .A2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1294), .B2(new_n1253), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1251), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1255), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(G384), .A2(new_n1295), .A3(new_n1251), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT124), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1290), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AOI211_X1 g1103(.A(KEYINPUT124), .B(new_n1289), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1299), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1288), .A2(new_n1307), .ZN(new_n1308));
  OAI221_X1 g1108(.A(new_n1279), .B1(new_n1288), .B2(new_n1306), .C1(new_n1308), .C2(KEYINPUT62), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1278), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1307), .A2(KEYINPUT63), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1288), .A2(new_n1312), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1273), .A2(new_n1276), .A3(new_n1279), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT63), .B1(new_n1288), .B2(new_n1307), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT125), .B1(new_n1288), .B2(new_n1306), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT125), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1304), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G378), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1230), .B2(G378), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1319), .B(new_n1320), .C1(new_n1322), .C2(new_n1265), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1318), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT126), .B1(new_n1317), .B2(new_n1324), .ZN(new_n1325));
  AOI211_X1 g1125(.A(new_n1265), .B(new_n1299), .C1(new_n1284), .C2(new_n1287), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1313), .B(new_n1314), .C1(new_n1326), .C2(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1318), .A2(new_n1323), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT126), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1327), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1311), .B1(new_n1325), .B2(new_n1330), .ZN(G405));
  XNOR2_X1  g1131(.A(new_n1230), .B(G378), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(new_n1307), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1277), .ZN(G402));
endmodule


