

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U555 ( .A1(n581), .A2(G2105), .ZN(n917) );
  NAND2_X1 U556 ( .A1(n670), .A2(n669), .ZN(n735) );
  XNOR2_X1 U557 ( .A(n668), .B(KEYINPUT93), .ZN(n669) );
  INV_X1 U558 ( .A(KEYINPUT30), .ZN(n547) );
  NAND2_X1 U559 ( .A1(n539), .A2(n547), .ZN(n538) );
  INV_X1 U560 ( .A(G1966), .ZN(n539) );
  AND2_X1 U561 ( .A1(n545), .A2(n541), .ZN(n540) );
  XNOR2_X1 U562 ( .A(n733), .B(KEYINPUT105), .ZN(n743) );
  NOR2_X1 U563 ( .A1(n732), .A2(n731), .ZN(n733) );
  INV_X1 U564 ( .A(n557), .ZN(n551) );
  NAND2_X1 U565 ( .A1(n531), .A2(n526), .ZN(n668) );
  INV_X1 U566 ( .A(G40), .ZN(n534) );
  XNOR2_X1 U567 ( .A(n536), .B(G2104), .ZN(n581) );
  INV_X1 U568 ( .A(KEYINPUT64), .ZN(n536) );
  NOR2_X1 U569 ( .A1(n724), .A2(n547), .ZN(n546) );
  NAND2_X1 U570 ( .A1(G1966), .A2(KEYINPUT30), .ZN(n544) );
  AND2_X1 U571 ( .A1(n549), .A2(n548), .ZN(n726) );
  XNOR2_X1 U572 ( .A(n529), .B(KEYINPUT32), .ZN(n770) );
  NAND2_X1 U573 ( .A1(n530), .A2(n740), .ZN(n529) );
  NAND2_X1 U574 ( .A1(n743), .A2(n734), .ZN(n530) );
  AND2_X1 U575 ( .A1(n558), .A2(n777), .ZN(n557) );
  NAND2_X1 U576 ( .A1(n559), .A2(KEYINPUT108), .ZN(n558) );
  INV_X1 U577 ( .A(n522), .ZN(n559) );
  XNOR2_X1 U578 ( .A(n591), .B(KEYINPUT23), .ZN(n535) );
  NAND2_X1 U579 ( .A1(n556), .A2(n555), .ZN(n792) );
  AND2_X1 U580 ( .A1(n526), .A2(n533), .ZN(G160) );
  NOR2_X1 U581 ( .A1(n593), .A2(n535), .ZN(n533) );
  NOR2_X2 U582 ( .A1(n581), .A2(G2105), .ZN(n590) );
  XOR2_X1 U583 ( .A(KEYINPUT98), .B(n661), .Z(n522) );
  XOR2_X1 U584 ( .A(KEYINPUT99), .B(n722), .Z(n756) );
  NOR2_X1 U585 ( .A1(n775), .A2(n774), .ZN(n523) );
  OR2_X1 U586 ( .A1(n756), .A2(n538), .ZN(n524) );
  NOR2_X1 U587 ( .A1(n768), .A2(n764), .ZN(n525) );
  XOR2_X1 U588 ( .A(n592), .B(KEYINPUT65), .Z(n526) );
  NOR2_X1 U589 ( .A1(n756), .A2(n755), .ZN(n527) );
  NAND2_X1 U590 ( .A1(n522), .A2(n560), .ZN(n528) );
  INV_X1 U591 ( .A(KEYINPUT108), .ZN(n560) );
  NOR2_X1 U592 ( .A1(n532), .A2(n535), .ZN(n531) );
  OR2_X1 U593 ( .A1(n593), .A2(n534), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n537), .A2(n544), .ZN(n543) );
  INV_X1 U595 ( .A(n724), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n756), .A2(G1966), .ZN(n745) );
  NAND2_X1 U597 ( .A1(n540), .A2(n524), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n724), .A2(KEYINPUT30), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n756), .A2(n546), .ZN(n545) );
  INV_X1 U601 ( .A(G168), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n550), .A2(n523), .ZN(n554) );
  NOR2_X1 U603 ( .A1(n776), .A2(n551), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n552), .A2(n523), .ZN(n555) );
  NOR2_X1 U605 ( .A1(n776), .A2(n560), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n554), .A2(n553), .ZN(n556) );
  NAND2_X1 U607 ( .A1(n557), .A2(n528), .ZN(n553) );
  NOR2_X1 U608 ( .A1(n735), .A2(n970), .ZN(n673) );
  INV_X1 U609 ( .A(KEYINPUT28), .ZN(n677) );
  INV_X1 U610 ( .A(KEYINPUT104), .ZN(n725) );
  NOR2_X1 U611 ( .A1(G164), .A2(G1384), .ZN(n670) );
  NOR2_X1 U612 ( .A1(G651), .A2(n617), .ZN(n823) );
  XNOR2_X1 U613 ( .A(G543), .B(KEYINPUT0), .ZN(n561) );
  XNOR2_X1 U614 ( .A(n561), .B(KEYINPUT67), .ZN(n617) );
  INV_X1 U615 ( .A(G651), .ZN(n568) );
  NOR2_X1 U616 ( .A1(n617), .A2(n568), .ZN(n828) );
  NAND2_X1 U617 ( .A1(G76), .A2(n828), .ZN(n565) );
  XOR2_X1 U618 ( .A(KEYINPUT4), .B(KEYINPUT79), .Z(n563) );
  NOR2_X1 U619 ( .A1(G651), .A2(G543), .ZN(n827) );
  NAND2_X1 U620 ( .A1(G89), .A2(n827), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U623 ( .A(n566), .B(KEYINPUT80), .ZN(n567) );
  XNOR2_X1 U624 ( .A(KEYINPUT5), .B(n567), .ZN(n576) );
  XNOR2_X1 U625 ( .A(KEYINPUT6), .B(KEYINPUT81), .ZN(n574) );
  NAND2_X1 U626 ( .A1(G51), .A2(n823), .ZN(n572) );
  NOR2_X1 U627 ( .A1(G543), .A2(n568), .ZN(n570) );
  XNOR2_X1 U628 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n570), .B(n569), .ZN(n824) );
  NAND2_X1 U630 ( .A1(G63), .A2(n824), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U632 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U634 ( .A(n577), .B(KEYINPUT7), .ZN(G168) );
  AND2_X1 U635 ( .A1(G2104), .A2(G2105), .ZN(n916) );
  NAND2_X1 U636 ( .A1(G114), .A2(n916), .ZN(n579) );
  NAND2_X1 U637 ( .A1(G126), .A2(n917), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U639 ( .A(KEYINPUT92), .B(n580), .ZN(n586) );
  NAND2_X1 U640 ( .A1(n590), .A2(G102), .ZN(n584) );
  NOR2_X1 U641 ( .A1(G2104), .A2(G2105), .ZN(n582) );
  XOR2_X1 U642 ( .A(KEYINPUT17), .B(n582), .Z(n587) );
  BUF_X1 U643 ( .A(n587), .Z(n902) );
  NAND2_X1 U644 ( .A1(n902), .A2(G138), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U646 ( .A1(n586), .A2(n585), .ZN(G164) );
  NAND2_X1 U647 ( .A1(G113), .A2(n916), .ZN(n589) );
  NAND2_X1 U648 ( .A1(G137), .A2(n587), .ZN(n588) );
  NAND2_X1 U649 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U650 ( .A1(G101), .A2(n590), .ZN(n591) );
  NAND2_X1 U651 ( .A1(G125), .A2(n917), .ZN(n592) );
  NAND2_X1 U652 ( .A1(G52), .A2(n823), .ZN(n595) );
  NAND2_X1 U653 ( .A1(G64), .A2(n824), .ZN(n594) );
  NAND2_X1 U654 ( .A1(n595), .A2(n594), .ZN(n601) );
  NAND2_X1 U655 ( .A1(G90), .A2(n827), .ZN(n597) );
  NAND2_X1 U656 ( .A1(G77), .A2(n828), .ZN(n596) );
  NAND2_X1 U657 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U658 ( .A(KEYINPUT71), .B(n598), .ZN(n599) );
  XNOR2_X1 U659 ( .A(KEYINPUT9), .B(n599), .ZN(n600) );
  NOR2_X1 U660 ( .A1(n601), .A2(n600), .ZN(G171) );
  INV_X1 U661 ( .A(G171), .ZN(G301) );
  XOR2_X1 U662 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U663 ( .A1(G88), .A2(n827), .ZN(n603) );
  NAND2_X1 U664 ( .A1(G75), .A2(n828), .ZN(n602) );
  NAND2_X1 U665 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U666 ( .A1(n824), .A2(G62), .ZN(n604) );
  XOR2_X1 U667 ( .A(KEYINPUT86), .B(n604), .Z(n605) );
  NOR2_X1 U668 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U669 ( .A1(n823), .A2(G50), .ZN(n607) );
  NAND2_X1 U670 ( .A1(n608), .A2(n607), .ZN(G303) );
  NAND2_X1 U671 ( .A1(G86), .A2(n827), .ZN(n610) );
  NAND2_X1 U672 ( .A1(G61), .A2(n824), .ZN(n609) );
  NAND2_X1 U673 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U674 ( .A1(G73), .A2(n828), .ZN(n611) );
  XNOR2_X1 U675 ( .A(n611), .B(KEYINPUT2), .ZN(n612) );
  XNOR2_X1 U676 ( .A(n612), .B(KEYINPUT85), .ZN(n613) );
  NOR2_X1 U677 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U678 ( .A1(n823), .A2(G48), .ZN(n615) );
  NAND2_X1 U679 ( .A1(n616), .A2(n615), .ZN(G305) );
  NAND2_X1 U680 ( .A1(G49), .A2(n823), .ZN(n619) );
  NAND2_X1 U681 ( .A1(G87), .A2(n617), .ZN(n618) );
  NAND2_X1 U682 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U683 ( .A1(n824), .A2(n620), .ZN(n622) );
  NAND2_X1 U684 ( .A1(G651), .A2(G74), .ZN(n621) );
  NAND2_X1 U685 ( .A1(n622), .A2(n621), .ZN(G288) );
  INV_X1 U686 ( .A(G303), .ZN(G166) );
  NAND2_X1 U687 ( .A1(n827), .A2(G85), .ZN(n623) );
  XNOR2_X1 U688 ( .A(n623), .B(KEYINPUT66), .ZN(n625) );
  NAND2_X1 U689 ( .A1(G72), .A2(n828), .ZN(n624) );
  NAND2_X1 U690 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U691 ( .A(KEYINPUT68), .B(n626), .ZN(n629) );
  NAND2_X1 U692 ( .A1(G47), .A2(n823), .ZN(n627) );
  XOR2_X1 U693 ( .A(KEYINPUT70), .B(n627), .Z(n628) );
  NOR2_X1 U694 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U695 ( .A1(n824), .A2(G60), .ZN(n630) );
  NAND2_X1 U696 ( .A1(n631), .A2(n630), .ZN(G290) );
  XOR2_X1 U697 ( .A(KEYINPUT93), .B(n668), .Z(n632) );
  NOR2_X1 U698 ( .A1(n670), .A2(n632), .ZN(n789) );
  XNOR2_X1 U699 ( .A(G2067), .B(KEYINPUT37), .ZN(n787) );
  NAND2_X1 U700 ( .A1(G116), .A2(n916), .ZN(n634) );
  NAND2_X1 U701 ( .A1(G128), .A2(n917), .ZN(n633) );
  NAND2_X1 U702 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U703 ( .A(n635), .B(KEYINPUT35), .ZN(n640) );
  NAND2_X1 U704 ( .A1(G140), .A2(n902), .ZN(n637) );
  NAND2_X1 U705 ( .A1(G104), .A2(n590), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U707 ( .A(KEYINPUT34), .B(n638), .Z(n639) );
  NAND2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U709 ( .A(n641), .B(KEYINPUT36), .Z(n929) );
  OR2_X1 U710 ( .A1(n787), .A2(n929), .ZN(n642) );
  XOR2_X1 U711 ( .A(KEYINPUT94), .B(n642), .Z(n963) );
  NAND2_X1 U712 ( .A1(n789), .A2(n963), .ZN(n785) );
  NAND2_X1 U713 ( .A1(G131), .A2(n902), .ZN(n644) );
  NAND2_X1 U714 ( .A1(G95), .A2(n590), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n649) );
  NAND2_X1 U716 ( .A1(G107), .A2(n916), .ZN(n646) );
  NAND2_X1 U717 ( .A1(G119), .A2(n917), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U719 ( .A(KEYINPUT95), .B(n647), .Z(n648) );
  NOR2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n927) );
  INV_X1 U721 ( .A(G1991), .ZN(n989) );
  NOR2_X1 U722 ( .A1(n927), .A2(n989), .ZN(n660) );
  NAND2_X1 U723 ( .A1(G141), .A2(n902), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n650), .B(KEYINPUT96), .ZN(n657) );
  NAND2_X1 U725 ( .A1(G117), .A2(n916), .ZN(n652) );
  NAND2_X1 U726 ( .A1(G129), .A2(n917), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n590), .A2(G105), .ZN(n653) );
  XOR2_X1 U729 ( .A(KEYINPUT38), .B(n653), .Z(n654) );
  NOR2_X1 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U732 ( .A(KEYINPUT97), .B(n658), .ZN(n924) );
  INV_X1 U733 ( .A(G1996), .ZN(n981) );
  NOR2_X1 U734 ( .A1(n924), .A2(n981), .ZN(n659) );
  OR2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n956) );
  NAND2_X1 U736 ( .A1(n956), .A2(n789), .ZN(n778) );
  NAND2_X1 U737 ( .A1(n785), .A2(n778), .ZN(n661) );
  NAND2_X1 U738 ( .A1(G53), .A2(n823), .ZN(n663) );
  NAND2_X1 U739 ( .A1(G65), .A2(n824), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U741 ( .A1(G91), .A2(n827), .ZN(n665) );
  NAND2_X1 U742 ( .A1(G78), .A2(n828), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U744 ( .A1(n667), .A2(n666), .ZN(n1018) );
  INV_X1 U745 ( .A(G2072), .ZN(n970) );
  XOR2_X1 U746 ( .A(KEYINPUT101), .B(KEYINPUT27), .Z(n671) );
  XNOR2_X1 U747 ( .A(KEYINPUT100), .B(n671), .ZN(n672) );
  XNOR2_X1 U748 ( .A(n673), .B(n672), .ZN(n675) );
  NAND2_X1 U749 ( .A1(n735), .A2(G1956), .ZN(n674) );
  NAND2_X1 U750 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U751 ( .A(KEYINPUT102), .B(n676), .Z(n679) );
  NOR2_X1 U752 ( .A1(n1018), .A2(n679), .ZN(n678) );
  XNOR2_X1 U753 ( .A(n678), .B(n677), .ZN(n715) );
  NAND2_X1 U754 ( .A1(n1018), .A2(n679), .ZN(n713) );
  NAND2_X1 U755 ( .A1(G92), .A2(n827), .ZN(n681) );
  NAND2_X1 U756 ( .A1(G66), .A2(n824), .ZN(n680) );
  NAND2_X1 U757 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U758 ( .A(KEYINPUT78), .B(n682), .ZN(n686) );
  NAND2_X1 U759 ( .A1(G79), .A2(n828), .ZN(n684) );
  NAND2_X1 U760 ( .A1(G54), .A2(n823), .ZN(n683) );
  NAND2_X1 U761 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U762 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U763 ( .A(KEYINPUT15), .B(n687), .Z(n821) );
  NAND2_X1 U764 ( .A1(G1348), .A2(n735), .ZN(n689) );
  INV_X1 U765 ( .A(n735), .ZN(n717) );
  NAND2_X1 U766 ( .A1(G2067), .A2(n717), .ZN(n688) );
  NAND2_X1 U767 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U768 ( .A(KEYINPUT103), .B(n690), .ZN(n709) );
  OR2_X1 U769 ( .A1(n821), .A2(n709), .ZN(n708) );
  NAND2_X1 U770 ( .A1(G56), .A2(n824), .ZN(n691) );
  XNOR2_X1 U771 ( .A(n691), .B(KEYINPUT75), .ZN(n692) );
  XNOR2_X1 U772 ( .A(KEYINPUT14), .B(n692), .ZN(n700) );
  XOR2_X1 U773 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n694) );
  NAND2_X1 U774 ( .A1(G81), .A2(n827), .ZN(n693) );
  XNOR2_X1 U775 ( .A(n694), .B(n693), .ZN(n697) );
  NAND2_X1 U776 ( .A1(n828), .A2(G68), .ZN(n695) );
  XNOR2_X1 U777 ( .A(KEYINPUT77), .B(n695), .ZN(n696) );
  NOR2_X1 U778 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U779 ( .A(KEYINPUT13), .B(n698), .ZN(n699) );
  NOR2_X1 U780 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U781 ( .A1(n823), .A2(G43), .ZN(n701) );
  NAND2_X1 U782 ( .A1(n702), .A2(n701), .ZN(n1025) );
  NOR2_X1 U783 ( .A1(n735), .A2(n981), .ZN(n703) );
  XOR2_X1 U784 ( .A(n703), .B(KEYINPUT26), .Z(n705) );
  NAND2_X1 U785 ( .A1(n735), .A2(G1341), .ZN(n704) );
  NAND2_X1 U786 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U787 ( .A1(n1025), .A2(n706), .ZN(n707) );
  NAND2_X1 U788 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U789 ( .A1(n709), .A2(n821), .ZN(n710) );
  AND2_X1 U790 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U791 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U792 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U793 ( .A(n716), .B(KEYINPUT29), .ZN(n721) );
  XOR2_X1 U794 ( .A(KEYINPUT25), .B(G2078), .Z(n986) );
  NOR2_X1 U795 ( .A1(n986), .A2(n735), .ZN(n719) );
  NOR2_X1 U796 ( .A1(n717), .A2(G1961), .ZN(n718) );
  NOR2_X1 U797 ( .A1(n719), .A2(n718), .ZN(n727) );
  NOR2_X1 U798 ( .A1(G301), .A2(n727), .ZN(n720) );
  NOR2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n732) );
  NAND2_X1 U800 ( .A1(n735), .A2(G8), .ZN(n722) );
  INV_X1 U801 ( .A(G8), .ZN(n723) );
  NOR2_X1 U802 ( .A1(G2084), .A2(n735), .ZN(n741) );
  OR2_X1 U803 ( .A1(n723), .A2(n741), .ZN(n724) );
  XNOR2_X1 U804 ( .A(n726), .B(n725), .ZN(n729) );
  NAND2_X1 U805 ( .A1(n727), .A2(G301), .ZN(n728) );
  NAND2_X1 U806 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U807 ( .A(KEYINPUT31), .B(n730), .Z(n731) );
  AND2_X1 U808 ( .A1(G286), .A2(G8), .ZN(n734) );
  NOR2_X1 U809 ( .A1(G2090), .A2(n735), .ZN(n737) );
  INV_X1 U810 ( .A(n756), .ZN(n767) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n756), .ZN(n736) );
  NOR2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U813 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U814 ( .A1(n723), .A2(n739), .ZN(n740) );
  INV_X1 U815 ( .A(n770), .ZN(n759) );
  NAND2_X1 U816 ( .A1(G8), .A2(n741), .ZN(n742) );
  NAND2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n768) );
  NOR2_X1 U819 ( .A1(G1981), .A2(G305), .ZN(n746) );
  XNOR2_X1 U820 ( .A(n746), .B(KEYINPUT24), .ZN(n747) );
  AND2_X1 U821 ( .A1(n747), .A2(n767), .ZN(n752) );
  INV_X1 U822 ( .A(n752), .ZN(n751) );
  NOR2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n1007) );
  AND2_X1 U824 ( .A1(n1007), .A2(KEYINPUT33), .ZN(n748) );
  AND2_X1 U825 ( .A1(n748), .A2(n767), .ZN(n749) );
  XNOR2_X1 U826 ( .A(G1981), .B(G305), .ZN(n1027) );
  OR2_X1 U827 ( .A1(n749), .A2(n1027), .ZN(n750) );
  AND2_X1 U828 ( .A1(n751), .A2(n750), .ZN(n755) );
  INV_X1 U829 ( .A(n755), .ZN(n754) );
  OR2_X1 U830 ( .A1(KEYINPUT33), .A2(n752), .ZN(n753) );
  NAND2_X1 U831 ( .A1(n754), .A2(n753), .ZN(n761) );
  INV_X1 U832 ( .A(n761), .ZN(n758) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n1008) );
  AND2_X1 U834 ( .A1(n527), .A2(n1008), .ZN(n757) );
  NOR2_X1 U835 ( .A1(n758), .A2(n757), .ZN(n764) );
  NAND2_X1 U836 ( .A1(n759), .A2(n525), .ZN(n766) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n1020) );
  NOR2_X1 U838 ( .A1(n1007), .A2(n1020), .ZN(n760) );
  XNOR2_X1 U839 ( .A(n760), .B(KEYINPUT106), .ZN(n762) );
  AND2_X1 U840 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U841 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U842 ( .A1(n766), .A2(n765), .ZN(n776) );
  OR2_X1 U843 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U844 ( .A1(n770), .A2(n769), .ZN(n775) );
  NAND2_X1 U845 ( .A1(G8), .A2(G166), .ZN(n771) );
  NOR2_X1 U846 ( .A1(G2090), .A2(n771), .ZN(n772) );
  XOR2_X1 U847 ( .A(KEYINPUT107), .B(n772), .Z(n773) );
  AND2_X1 U848 ( .A1(n756), .A2(n773), .ZN(n774) );
  XNOR2_X1 U849 ( .A(G1986), .B(G290), .ZN(n1012) );
  NAND2_X1 U850 ( .A1(n1012), .A2(n789), .ZN(n777) );
  AND2_X1 U851 ( .A1(n981), .A2(n924), .ZN(n967) );
  INV_X1 U852 ( .A(n778), .ZN(n782) );
  NOR2_X1 U853 ( .A1(G1986), .A2(G290), .ZN(n780) );
  AND2_X1 U854 ( .A1(n989), .A2(n927), .ZN(n779) );
  XOR2_X1 U855 ( .A(KEYINPUT109), .B(n779), .Z(n957) );
  NOR2_X1 U856 ( .A1(n780), .A2(n957), .ZN(n781) );
  NOR2_X1 U857 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U858 ( .A1(n967), .A2(n783), .ZN(n784) );
  XNOR2_X1 U859 ( .A(KEYINPUT39), .B(n784), .ZN(n786) );
  NAND2_X1 U860 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U861 ( .A1(n929), .A2(n787), .ZN(n960) );
  NAND2_X1 U862 ( .A1(n788), .A2(n960), .ZN(n790) );
  NAND2_X1 U863 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U864 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U865 ( .A(n793), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U866 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U867 ( .A(G132), .ZN(G219) );
  INV_X1 U868 ( .A(G82), .ZN(G220) );
  INV_X1 U869 ( .A(G57), .ZN(G237) );
  INV_X1 U870 ( .A(G108), .ZN(G238) );
  INV_X1 U871 ( .A(G120), .ZN(G236) );
  XOR2_X1 U872 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n795) );
  NAND2_X1 U873 ( .A1(G7), .A2(G661), .ZN(n794) );
  XNOR2_X1 U874 ( .A(n795), .B(n794), .ZN(n796) );
  XNOR2_X1 U875 ( .A(KEYINPUT72), .B(n796), .ZN(G223) );
  XOR2_X1 U876 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n798) );
  INV_X1 U877 ( .A(G223), .ZN(n862) );
  NAND2_X1 U878 ( .A1(n862), .A2(G567), .ZN(n797) );
  XNOR2_X1 U879 ( .A(n798), .B(n797), .ZN(G234) );
  INV_X1 U880 ( .A(G860), .ZN(n805) );
  OR2_X1 U881 ( .A1(n1025), .A2(n805), .ZN(G153) );
  NAND2_X1 U882 ( .A1(G868), .A2(G301), .ZN(n800) );
  INV_X1 U883 ( .A(n821), .ZN(n1015) );
  INV_X1 U884 ( .A(G868), .ZN(n802) );
  NAND2_X1 U885 ( .A1(n1015), .A2(n802), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(G284) );
  INV_X1 U887 ( .A(n1018), .ZN(G299) );
  NOR2_X1 U888 ( .A1(G868), .A2(G299), .ZN(n801) );
  XNOR2_X1 U889 ( .A(n801), .B(KEYINPUT82), .ZN(n804) );
  NOR2_X1 U890 ( .A1(n802), .A2(G286), .ZN(n803) );
  NOR2_X1 U891 ( .A1(n804), .A2(n803), .ZN(G297) );
  NAND2_X1 U892 ( .A1(n805), .A2(G559), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n806), .A2(n821), .ZN(n807) );
  XNOR2_X1 U894 ( .A(n807), .B(KEYINPUT83), .ZN(n808) );
  XOR2_X1 U895 ( .A(KEYINPUT16), .B(n808), .Z(G148) );
  NOR2_X1 U896 ( .A1(G868), .A2(n1025), .ZN(n811) );
  NAND2_X1 U897 ( .A1(G868), .A2(n821), .ZN(n809) );
  NOR2_X1 U898 ( .A1(G559), .A2(n809), .ZN(n810) );
  NOR2_X1 U899 ( .A1(n811), .A2(n810), .ZN(G282) );
  XOR2_X1 U900 ( .A(G2100), .B(KEYINPUT84), .Z(n820) );
  NAND2_X1 U901 ( .A1(G111), .A2(n916), .ZN(n813) );
  NAND2_X1 U902 ( .A1(G135), .A2(n902), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n818) );
  NAND2_X1 U904 ( .A1(n917), .A2(G123), .ZN(n814) );
  XNOR2_X1 U905 ( .A(n814), .B(KEYINPUT18), .ZN(n816) );
  NAND2_X1 U906 ( .A1(G99), .A2(n590), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n959) );
  XNOR2_X1 U909 ( .A(G2096), .B(n959), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(G156) );
  NAND2_X1 U911 ( .A1(n821), .A2(G559), .ZN(n840) );
  XNOR2_X1 U912 ( .A(n1025), .B(n840), .ZN(n822) );
  NOR2_X1 U913 ( .A1(n822), .A2(G860), .ZN(n833) );
  NAND2_X1 U914 ( .A1(G55), .A2(n823), .ZN(n826) );
  NAND2_X1 U915 ( .A1(G67), .A2(n824), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n826), .A2(n825), .ZN(n832) );
  NAND2_X1 U917 ( .A1(G93), .A2(n827), .ZN(n830) );
  NAND2_X1 U918 ( .A1(G80), .A2(n828), .ZN(n829) );
  NAND2_X1 U919 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U920 ( .A1(n832), .A2(n831), .ZN(n843) );
  XNOR2_X1 U921 ( .A(n833), .B(n843), .ZN(G145) );
  XOR2_X1 U922 ( .A(KEYINPUT19), .B(n843), .Z(n834) );
  XNOR2_X1 U923 ( .A(G288), .B(n834), .ZN(n835) );
  XNOR2_X1 U924 ( .A(n1018), .B(n835), .ZN(n838) );
  XNOR2_X1 U925 ( .A(n1025), .B(G303), .ZN(n836) );
  XNOR2_X1 U926 ( .A(n836), .B(G305), .ZN(n837) );
  XNOR2_X1 U927 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U928 ( .A(G290), .B(n839), .ZN(n935) );
  XNOR2_X1 U929 ( .A(n935), .B(n840), .ZN(n841) );
  NAND2_X1 U930 ( .A1(n841), .A2(G868), .ZN(n842) );
  XNOR2_X1 U931 ( .A(KEYINPUT87), .B(n842), .ZN(n846) );
  NOR2_X1 U932 ( .A1(G868), .A2(n843), .ZN(n844) );
  XNOR2_X1 U933 ( .A(n844), .B(KEYINPUT88), .ZN(n845) );
  NOR2_X1 U934 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U935 ( .A(KEYINPUT89), .B(n847), .ZN(G295) );
  NAND2_X1 U936 ( .A1(G2078), .A2(G2084), .ZN(n848) );
  XOR2_X1 U937 ( .A(KEYINPUT20), .B(n848), .Z(n849) );
  NAND2_X1 U938 ( .A1(G2090), .A2(n849), .ZN(n850) );
  XNOR2_X1 U939 ( .A(KEYINPUT21), .B(n850), .ZN(n851) );
  NAND2_X1 U940 ( .A1(n851), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U941 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U942 ( .A1(G236), .A2(G238), .ZN(n852) );
  NAND2_X1 U943 ( .A1(G69), .A2(n852), .ZN(n853) );
  NOR2_X1 U944 ( .A1(n853), .A2(G237), .ZN(n854) );
  XNOR2_X1 U945 ( .A(n854), .B(KEYINPUT91), .ZN(n868) );
  NAND2_X1 U946 ( .A1(n868), .A2(G567), .ZN(n860) );
  NOR2_X1 U947 ( .A1(G220), .A2(G219), .ZN(n855) );
  XNOR2_X1 U948 ( .A(KEYINPUT22), .B(n855), .ZN(n856) );
  NAND2_X1 U949 ( .A1(n856), .A2(G96), .ZN(n857) );
  NOR2_X1 U950 ( .A1(G218), .A2(n857), .ZN(n858) );
  XOR2_X1 U951 ( .A(KEYINPUT90), .B(n858), .Z(n869) );
  NAND2_X1 U952 ( .A1(n869), .A2(G2106), .ZN(n859) );
  NAND2_X1 U953 ( .A1(n860), .A2(n859), .ZN(n891) );
  NAND2_X1 U954 ( .A1(G483), .A2(G661), .ZN(n861) );
  NOR2_X1 U955 ( .A1(n891), .A2(n861), .ZN(n867) );
  NAND2_X1 U956 ( .A1(n867), .A2(G36), .ZN(G176) );
  NAND2_X1 U957 ( .A1(n862), .A2(G2106), .ZN(n863) );
  XNOR2_X1 U958 ( .A(n863), .B(KEYINPUT110), .ZN(G217) );
  AND2_X1 U959 ( .A1(G15), .A2(G2), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G661), .A2(n864), .ZN(G259) );
  NAND2_X1 U961 ( .A1(G3), .A2(G1), .ZN(n865) );
  XOR2_X1 U962 ( .A(KEYINPUT111), .B(n865), .Z(n866) );
  NAND2_X1 U963 ( .A1(n867), .A2(n866), .ZN(G188) );
  INV_X1 U965 ( .A(G96), .ZN(G221) );
  NOR2_X1 U966 ( .A1(n869), .A2(n868), .ZN(G325) );
  INV_X1 U967 ( .A(G325), .ZN(G261) );
  XOR2_X1 U968 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n871) );
  XNOR2_X1 U969 ( .A(G2096), .B(G2678), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U971 ( .A(n872), .B(G2100), .Z(n874) );
  XNOR2_X1 U972 ( .A(G2078), .B(G2084), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U974 ( .A(KEYINPUT42), .B(G2090), .Z(n876) );
  XNOR2_X1 U975 ( .A(G2067), .B(G2072), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U977 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U978 ( .A(KEYINPUT114), .B(KEYINPUT43), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n880), .B(n879), .ZN(G227) );
  XOR2_X1 U980 ( .A(G1976), .B(G1971), .Z(n882) );
  XNOR2_X1 U981 ( .A(G1986), .B(G1956), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n886) );
  XOR2_X1 U983 ( .A(G1981), .B(G1966), .Z(n884) );
  XNOR2_X1 U984 ( .A(G1996), .B(G1991), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U987 ( .A(KEYINPUT115), .B(G2474), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n890) );
  XOR2_X1 U989 ( .A(G1961), .B(KEYINPUT41), .Z(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(G229) );
  INV_X1 U991 ( .A(n891), .ZN(G319) );
  NAND2_X1 U992 ( .A1(n590), .A2(G100), .ZN(n898) );
  NAND2_X1 U993 ( .A1(G112), .A2(n916), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G136), .A2(n587), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n896) );
  NAND2_X1 U996 ( .A1(n917), .A2(G124), .ZN(n894) );
  XOR2_X1 U997 ( .A(KEYINPUT44), .B(n894), .Z(n895) );
  NOR2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n897) );
  NAND2_X1 U999 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U1000 ( .A(KEYINPUT116), .B(n899), .Z(G162) );
  NAND2_X1 U1001 ( .A1(G118), .A2(n916), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(G130), .A2(n917), .ZN(n900) );
  NAND2_X1 U1003 ( .A1(n901), .A2(n900), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(G142), .A2(n902), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(G106), .A2(n590), .ZN(n903) );
  NAND2_X1 U1006 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1007 ( .A(n905), .B(KEYINPUT45), .Z(n906) );
  NOR2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n908), .B(G162), .ZN(n933) );
  XOR2_X1 U1010 ( .A(KEYINPUT118), .B(KEYINPUT120), .Z(n910) );
  XNOR2_X1 U1011 ( .A(KEYINPUT48), .B(KEYINPUT117), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1013 ( .A(n911), .B(KEYINPUT46), .Z(n913) );
  XNOR2_X1 U1014 ( .A(n959), .B(KEYINPUT119), .ZN(n912) );
  XNOR2_X1 U1015 ( .A(n913), .B(n912), .ZN(n923) );
  NAND2_X1 U1016 ( .A1(G139), .A2(n587), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(G103), .A2(n590), .ZN(n914) );
  NAND2_X1 U1018 ( .A1(n915), .A2(n914), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(G115), .A2(n916), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(G127), .A2(n917), .ZN(n918) );
  NAND2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1022 ( .A(KEYINPUT47), .B(n920), .Z(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n969) );
  XOR2_X1 U1024 ( .A(n923), .B(n969), .Z(n926) );
  XNOR2_X1 U1025 ( .A(G164), .B(n924), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n926), .B(n925), .ZN(n928) );
  XOR2_X1 U1027 ( .A(n928), .B(n927), .Z(n931) );
  XOR2_X1 U1028 ( .A(G160), .B(n929), .Z(n930) );
  XNOR2_X1 U1029 ( .A(n931), .B(n930), .ZN(n932) );
  XOR2_X1 U1030 ( .A(n933), .B(n932), .Z(n934) );
  NOR2_X1 U1031 ( .A1(G37), .A2(n934), .ZN(G395) );
  XNOR2_X1 U1032 ( .A(G286), .B(n1015), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(n936), .B(n935), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(n937), .B(G171), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(G37), .A2(n938), .ZN(G397) );
  NOR2_X1 U1036 ( .A1(G227), .A2(G229), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(n940), .B(n939), .ZN(n941) );
  XOR2_X1 U1039 ( .A(KEYINPUT49), .B(n941), .Z(n952) );
  XOR2_X1 U1040 ( .A(G2451), .B(G2430), .Z(n943) );
  XNOR2_X1 U1041 ( .A(G2438), .B(G2443), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(n943), .B(n942), .ZN(n949) );
  XOR2_X1 U1043 ( .A(G2435), .B(G2454), .Z(n945) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G1348), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(n945), .B(n944), .ZN(n947) );
  XOR2_X1 U1046 ( .A(G2446), .B(G2427), .Z(n946) );
  XNOR2_X1 U1047 ( .A(n947), .B(n946), .ZN(n948) );
  XOR2_X1 U1048 ( .A(n949), .B(n948), .Z(n950) );
  NAND2_X1 U1049 ( .A1(G14), .A2(n950), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(G319), .A2(n955), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(G395), .A2(G397), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(G225) );
  INV_X1 U1054 ( .A(G225), .ZN(G308) );
  INV_X1 U1055 ( .A(G69), .ZN(G235) );
  INV_X1 U1056 ( .A(n955), .ZN(G401) );
  NOR2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n965) );
  XOR2_X1 U1058 ( .A(G2084), .B(G160), .Z(n958) );
  NOR2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n977) );
  XOR2_X1 U1063 ( .A(G2090), .B(G162), .Z(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1065 ( .A(KEYINPUT51), .B(n968), .Z(n975) );
  XOR2_X1 U1066 ( .A(G164), .B(G2078), .Z(n972) );
  XNOR2_X1 U1067 ( .A(n970), .B(n969), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(KEYINPUT50), .B(n973), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(KEYINPUT52), .B(n978), .ZN(n979) );
  INV_X1 U1073 ( .A(KEYINPUT55), .ZN(n1003) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n1003), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n980), .A2(G29), .ZN(n1063) );
  XOR2_X1 U1076 ( .A(G2090), .B(G35), .Z(n997) );
  XNOR2_X1 U1077 ( .A(G32), .B(n981), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(G2067), .B(G26), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(G2072), .B(G33), .ZN(n982) );
  NOR2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(G27), .B(n986), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n989), .B(G25), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n990), .A2(G28), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(n991), .B(KEYINPUT123), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1088 ( .A(n994), .B(KEYINPUT124), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n995), .B(KEYINPUT53), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(n998), .B(KEYINPUT125), .ZN(n1001) );
  XOR2_X1 U1092 ( .A(G2084), .B(G34), .Z(n999) );
  XNOR2_X1 U1093 ( .A(KEYINPUT54), .B(n999), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1095 ( .A(n1003), .B(n1002), .ZN(n1005) );
  INV_X1 U1096 ( .A(G29), .ZN(n1004) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(G11), .A2(n1006), .ZN(n1061) );
  XNOR2_X1 U1099 ( .A(G16), .B(KEYINPUT56), .ZN(n1034) );
  INV_X1 U1100 ( .A(n1007), .ZN(n1009) );
  NAND2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(G1971), .A2(G303), .ZN(n1013) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1024) );
  XNOR2_X1 U1106 ( .A(G301), .B(G1961), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(n1015), .B(G1348), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(G1956), .B(n1018), .Z(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1032) );
  XNOR2_X1 U1113 ( .A(n1025), .B(G1341), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(G1966), .B(G168), .Z(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT57), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1059) );
  INV_X1 U1120 ( .A(G16), .ZN(n1057) );
  XOR2_X1 U1121 ( .A(G1966), .B(G21), .Z(n1044) );
  XNOR2_X1 U1122 ( .A(G1348), .B(KEYINPUT59), .ZN(n1035) );
  XNOR2_X1 U1123 ( .A(n1035), .B(G4), .ZN(n1039) );
  XNOR2_X1 U1124 ( .A(G1341), .B(G19), .ZN(n1037) );
  XNOR2_X1 U1125 ( .A(G6), .B(G1981), .ZN(n1036) );
  NOR2_X1 U1126 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1127 ( .A1(n1039), .A2(n1038), .ZN(n1041) );
  XNOR2_X1 U1128 ( .A(G20), .B(G1956), .ZN(n1040) );
  NOR2_X1 U1129 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1130 ( .A(n1042), .B(KEYINPUT60), .ZN(n1043) );
  NAND2_X1 U1131 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1132 ( .A(KEYINPUT127), .B(n1045), .ZN(n1054) );
  XNOR2_X1 U1133 ( .A(G1961), .B(G5), .ZN(n1052) );
  XNOR2_X1 U1134 ( .A(G1971), .B(G22), .ZN(n1047) );
  XNOR2_X1 U1135 ( .A(G23), .B(G1976), .ZN(n1046) );
  NOR2_X1 U1136 ( .A1(n1047), .A2(n1046), .ZN(n1049) );
  XOR2_X1 U1137 ( .A(G1986), .B(G24), .Z(n1048) );
  NAND2_X1 U1138 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XNOR2_X1 U1139 ( .A(KEYINPUT58), .B(n1050), .ZN(n1051) );
  NOR2_X1 U1140 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  NAND2_X1 U1141 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  XOR2_X1 U1142 ( .A(KEYINPUT61), .B(n1055), .Z(n1056) );
  NAND2_X1 U1143 ( .A1(n1057), .A2(n1056), .ZN(n1058) );
  NAND2_X1 U1144 ( .A1(n1059), .A2(n1058), .ZN(n1060) );
  NOR2_X1 U1145 ( .A1(n1061), .A2(n1060), .ZN(n1062) );
  NAND2_X1 U1146 ( .A1(n1063), .A2(n1062), .ZN(n1064) );
  XOR2_X1 U1147 ( .A(KEYINPUT62), .B(n1064), .Z(G311) );
  INV_X1 U1148 ( .A(G311), .ZN(G150) );
endmodule

