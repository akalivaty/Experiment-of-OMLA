//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  INV_X1    g0000(.A(KEYINPUT65), .ZN(new_n201));
  XNOR2_X1  g0001(.A(KEYINPUT64), .B(G50), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  AOI21_X1  g0003(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  AND2_X1   g0004(.A1(KEYINPUT64), .A2(G50), .ZN(new_n205));
  NOR2_X1   g0005(.A1(KEYINPUT64), .A2(G50), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n201), .B(new_n203), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n204), .A2(new_n208), .A3(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G97), .A2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G58), .C2(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G1), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT67), .Z(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n228), .A2(new_n222), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(new_n225), .B2(KEYINPUT1), .ZN(new_n231));
  INV_X1    g0031(.A(new_n223), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT0), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n227), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT2), .ZN(new_n241));
  INV_X1    g0041(.A(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G264), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n213), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT69), .ZN(new_n250));
  INV_X1    g0050(.A(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n212), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT70), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G68), .B(G77), .ZN(new_n255));
  INV_X1    g0055(.A(G50), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n254), .B(new_n259), .ZN(G351));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(KEYINPUT7), .B1(new_n263), .B2(new_n222), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  AND4_X1   g0068(.A1(KEYINPUT7), .A2(new_n267), .A3(new_n222), .A4(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(G68), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G159), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n258), .A2(KEYINPUT73), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT73), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n217), .ZN(new_n277));
  OAI21_X1  g0077(.A(G20), .B1(new_n277), .B2(new_n203), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n270), .A2(new_n272), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT16), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n229), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n270), .A2(new_n278), .A3(KEYINPUT16), .A4(new_n272), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT8), .A2(G58), .ZN(new_n286));
  INV_X1    g0086(.A(new_n276), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(KEYINPUT8), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n221), .A2(G13), .A3(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT75), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT75), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n292), .A2(new_n221), .A3(G13), .A4(G20), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  AOI211_X1 g0095(.A(new_n283), .B(new_n294), .C1(new_n221), .C2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n288), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n285), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT79), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n267), .A2(new_n268), .ZN(new_n300));
  INV_X1    g0100(.A(G1698), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(G223), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G87), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(G1698), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n302), .B(new_n303), .C1(new_n304), .C2(new_n242), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT72), .B1(new_n307), .B2(new_n229), .ZN(new_n308));
  INV_X1    g0108(.A(new_n229), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(new_n310), .A3(new_n306), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n307), .A2(new_n229), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n221), .B1(G41), .B2(G45), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G232), .ZN(new_n318));
  INV_X1    g0118(.A(G274), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n313), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n299), .B1(new_n322), .B2(G179), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n305), .B2(new_n312), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(KEYINPUT79), .A3(new_n325), .A4(new_n318), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n298), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT18), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n298), .A2(new_n327), .A3(KEYINPUT18), .A4(new_n329), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n285), .A2(new_n295), .A3(new_n297), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n322), .A2(G200), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n324), .A2(G190), .A3(new_n318), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n335), .A2(new_n336), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n285), .A2(new_n295), .A3(new_n297), .A4(new_n338), .ZN(new_n340));
  INV_X1    g0140(.A(new_n337), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT17), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n334), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n296), .A2(G68), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n266), .A2(G20), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(G77), .B1(new_n271), .B2(G50), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n222), .B2(G68), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n348), .A2(new_n283), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n349), .A2(KEYINPUT11), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n294), .A2(new_n217), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT12), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(KEYINPUT11), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n345), .A2(new_n350), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  OAI211_X1 g0154(.A(G226), .B(new_n301), .C1(new_n261), .C2(new_n262), .ZN(new_n355));
  OAI211_X1 g0155(.A(G232), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G97), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n312), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n317), .A2(G238), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n312), .A3(KEYINPUT78), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n361), .A2(new_n321), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT13), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n320), .B1(new_n359), .B2(new_n360), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(new_n362), .A4(new_n363), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n354), .B1(new_n369), .B2(G200), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(G190), .A3(new_n368), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT76), .ZN(new_n375));
  OR2_X1    g0175(.A1(KEYINPUT15), .A2(G87), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT76), .ZN(new_n377));
  NAND2_X1  g0177(.A1(KEYINPUT15), .A2(G87), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n346), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT8), .B(G58), .Z(new_n383));
  AOI22_X1  g0183(.A1(new_n382), .A2(KEYINPUT77), .B1(new_n271), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G20), .A2(G77), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(new_n385), .C1(KEYINPUT77), .C2(new_n382), .ZN(new_n386));
  INV_X1    g0186(.A(G77), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n386), .A2(new_n283), .B1(new_n387), .B2(new_n294), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n300), .A2(G232), .A3(new_n301), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n389), .B1(new_n251), .B2(new_n300), .C1(new_n304), .C2(new_n218), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n312), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n317), .A2(G244), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n321), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G200), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n296), .A2(G77), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n388), .A2(new_n394), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n344), .A2(new_n373), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n369), .B2(G169), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n369), .A2(new_n325), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n369), .A2(new_n401), .A3(G169), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n354), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n300), .A2(G223), .A3(G1698), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n300), .A2(G222), .A3(new_n301), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n263), .A2(G77), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT71), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n312), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n317), .A2(G226), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n321), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n418), .A2(G179), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n291), .A2(new_n293), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(G50), .ZN(new_n421));
  OAI21_X1  g0221(.A(G20), .B1(new_n204), .B2(new_n208), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT74), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g0224(.A(KEYINPUT74), .B(G20), .C1(new_n204), .C2(new_n208), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n271), .A2(G150), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n288), .A2(new_n346), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n421), .B1(new_n428), .B2(new_n283), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n296), .A2(G50), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n418), .A2(new_n328), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n419), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT9), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n418), .A2(new_n395), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n429), .A2(KEYINPUT9), .A3(new_n430), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n418), .A2(G200), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n436), .A2(new_n437), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT10), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT10), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n442), .A2(new_n443), .A3(new_n437), .A4(new_n436), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n434), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n388), .A2(new_n397), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n393), .A2(new_n328), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n393), .A2(G179), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AND4_X1   g0249(.A1(new_n400), .A2(new_n408), .A3(new_n445), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT21), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT82), .ZN(new_n453));
  INV_X1    g0253(.A(G41), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n221), .A2(G45), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(KEYINPUT5), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G41), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(KEYINPUT82), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n457), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G270), .A3(new_n315), .ZN(new_n465));
  OAI211_X1 g0265(.A(G257), .B(new_n301), .C1(new_n261), .C2(new_n262), .ZN(new_n466));
  OAI211_X1 g0266(.A(G264), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n267), .A2(G303), .A3(new_n268), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n312), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n457), .A2(new_n463), .A3(G274), .A4(new_n458), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n465), .B(new_n470), .C1(new_n314), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n294), .A2(new_n212), .ZN(new_n473));
  INV_X1    g0273(.A(new_n283), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n266), .A2(G1), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n420), .A2(new_n474), .A3(G116), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n212), .A2(G20), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n283), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n222), .C1(G33), .C2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT20), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n283), .A3(new_n478), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT20), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n473), .B(new_n477), .C1(new_n483), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n472), .A2(G169), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n221), .B(G45), .C1(new_n454), .C2(KEYINPUT5), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n453), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT82), .B1(new_n460), .B2(new_n462), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(G274), .A3(new_n315), .A4(new_n458), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(G179), .A3(new_n470), .A4(new_n465), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n452), .A2(new_n488), .B1(new_n495), .B2(new_n487), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n472), .A2(KEYINPUT21), .A3(G169), .A4(new_n487), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT87), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n484), .A2(new_n485), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n499), .A2(new_n500), .B1(new_n212), .B2(new_n294), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n328), .B1(new_n501), .B2(new_n477), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT87), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT21), .A4(new_n472), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G200), .ZN(new_n506));
  OAI211_X1 g0306(.A(G257), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n507));
  OAI211_X1 g0307(.A(G250), .B(new_n301), .C1(new_n261), .C2(new_n262), .ZN(new_n508));
  INV_X1    g0308(.A(G294), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n507), .B(new_n508), .C1(new_n266), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n312), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n464), .A2(G264), .A3(new_n315), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n471), .A2(new_n314), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n506), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n493), .A2(new_n395), .A3(new_n511), .A4(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI211_X1 g0317(.A(new_n475), .B(new_n283), .C1(new_n291), .C2(new_n293), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G107), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n222), .B(G87), .C1(new_n261), .C2(new_n262), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT22), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n300), .A2(new_n523), .A3(new_n222), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n346), .A2(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n251), .A2(G20), .ZN(new_n527));
  XNOR2_X1  g0327(.A(new_n527), .B(KEYINPUT23), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AND4_X1   g0329(.A1(new_n520), .A2(new_n525), .A3(new_n526), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n522), .B2(new_n524), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n520), .B1(new_n531), .B2(new_n526), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n283), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n420), .A2(G107), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT25), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n517), .A2(new_n519), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n472), .A2(G200), .ZN(new_n537));
  INV_X1    g0337(.A(new_n487), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(new_n395), .C2(new_n472), .ZN(new_n539));
  AND4_X1   g0339(.A1(new_n496), .A2(new_n505), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n533), .A2(new_n519), .A3(new_n535), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n511), .A2(new_n512), .ZN(new_n542));
  AOI21_X1  g0342(.A(G169), .B1(new_n542), .B2(new_n493), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n513), .A2(G179), .A3(new_n514), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G250), .B(new_n456), .C1(new_n307), .C2(new_n229), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G244), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n549));
  OAI211_X1 g0349(.A(G238), .B(new_n301), .C1(new_n261), .C2(new_n262), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G116), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n548), .B1(new_n552), .B2(new_n312), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n460), .A2(G274), .ZN(new_n554));
  AOI21_X1  g0354(.A(G169), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n283), .B1(new_n291), .B2(new_n293), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(new_n379), .A3(new_n375), .A4(new_n476), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n222), .B1(new_n357), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(G97), .A2(G107), .ZN(new_n560));
  INV_X1    g0360(.A(G87), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n222), .B(G68), .C1(new_n261), .C2(new_n262), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n558), .B1(new_n357), .B2(G20), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n283), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n380), .A2(new_n294), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n557), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT86), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT86), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n557), .A2(new_n567), .A3(new_n568), .A4(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n555), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n552), .A2(new_n312), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n554), .A3(new_n547), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n325), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n556), .A2(new_n476), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n567), .B(new_n568), .C1(new_n578), .C2(new_n561), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(G200), .B2(new_n575), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(G190), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n573), .A2(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n546), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT84), .ZN(new_n584));
  OAI211_X1 g0384(.A(G244), .B(new_n301), .C1(new_n261), .C2(new_n262), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT4), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n300), .A2(KEYINPUT4), .A3(G244), .A4(new_n301), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n300), .A2(G250), .A3(G1698), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n480), .A4(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n590), .A2(new_n312), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n464), .A2(G257), .A3(new_n315), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n493), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n584), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(new_n312), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n595), .A2(KEYINPUT84), .A3(new_n493), .A4(new_n592), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n328), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n493), .A3(new_n592), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n325), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT81), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n481), .B1(new_n556), .B2(new_n476), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n420), .A2(new_n481), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n601), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(KEYINPUT81), .B(new_n603), .C1(new_n518), .C2(new_n481), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT6), .ZN(new_n608));
  AND2_X1   g0408(.A1(G97), .A2(G107), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(new_n560), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n251), .A2(KEYINPUT6), .A3(G97), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n222), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n271), .A2(G77), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT80), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT80), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n251), .A2(KEYINPUT6), .A3(G97), .ZN(new_n617));
  XNOR2_X1  g0417(.A(G97), .B(G107), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n608), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n616), .B(new_n613), .C1(new_n619), .C2(new_n222), .ZN(new_n620));
  OAI21_X1  g0420(.A(G107), .B1(new_n264), .B2(new_n269), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n615), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n283), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n607), .A2(new_n623), .A3(KEYINPUT85), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT85), .B1(new_n607), .B2(new_n623), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n597), .B(new_n600), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n598), .A2(G200), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT83), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n598), .A2(KEYINPUT83), .A3(G200), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n607), .A2(new_n623), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n493), .A2(new_n592), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT84), .B1(new_n634), .B2(new_n595), .ZN(new_n635));
  AND4_X1   g0435(.A1(KEYINPUT84), .A2(new_n595), .A3(new_n493), .A4(new_n592), .ZN(new_n636));
  OAI21_X1  g0436(.A(G190), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n631), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n540), .A2(new_n583), .A3(new_n626), .A4(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n451), .A2(new_n639), .ZN(G372));
  INV_X1    g0440(.A(new_n449), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n641), .A2(new_n372), .B1(new_n354), .B2(new_n407), .ZN(new_n642));
  INV_X1    g0442(.A(new_n343), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n334), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n441), .A2(new_n444), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n434), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n597), .A2(new_n600), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT88), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n570), .A2(new_n572), .B1(new_n555), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n575), .A2(new_n328), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n651), .A2(KEYINPUT88), .B1(new_n576), .B2(new_n325), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n650), .A2(new_n652), .B1(new_n581), .B2(new_n580), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n647), .A2(new_n648), .A3(new_n653), .A4(new_n632), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT85), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n632), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n607), .A2(new_n623), .A3(KEYINPUT85), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n658), .A2(new_n582), .A3(new_n597), .A4(new_n600), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n659), .A2(KEYINPUT26), .B1(new_n650), .B2(new_n652), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n505), .A2(KEYINPUT89), .A3(new_n496), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT89), .B1(new_n505), .B2(new_n496), .ZN(new_n662));
  INV_X1    g0462(.A(new_n546), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n638), .A2(new_n536), .A3(new_n626), .A4(new_n653), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n654), .B(new_n660), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n646), .B1(new_n451), .B2(new_n667), .ZN(G369));
  INV_X1    g0468(.A(G13), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(G20), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n221), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(KEYINPUT90), .B(G343), .Z(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n538), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n661), .B2(new_n662), .ZN(new_n680));
  INV_X1    g0480(.A(new_n679), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n505), .A2(new_n496), .A3(new_n539), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT91), .Z(new_n684));
  NOR2_X1   g0484(.A1(new_n546), .A2(new_n677), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n541), .A2(new_n677), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n536), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n546), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n684), .A2(G330), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n677), .B1(new_n505), .B2(new_n496), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n546), .B2(new_n677), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n689), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  INV_X1    g0494(.A(new_n665), .ZN(new_n695));
  INV_X1    g0495(.A(new_n662), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n505), .A2(new_n496), .A3(KEYINPUT89), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n546), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n573), .A2(new_n577), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n580), .A2(new_n581), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT26), .B1(new_n626), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n650), .A2(new_n652), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(new_n704), .A3(new_n654), .ZN(new_n705));
  AOI211_X1 g0505(.A(KEYINPUT96), .B(new_n677), .C1(new_n699), .C2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT96), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n666), .B2(new_n678), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n694), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT97), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n647), .A2(new_n648), .A3(new_n658), .A4(new_n582), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n546), .A2(new_n496), .A3(new_n505), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n711), .B(new_n704), .C1(new_n665), .C2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n647), .A2(new_n632), .A3(new_n653), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(KEYINPUT26), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT29), .B(new_n678), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT97), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n694), .C1(new_n706), .C2(new_n708), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n710), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G330), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT31), .B1(new_n639), .B2(new_n677), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n494), .A2(new_n513), .A3(new_n575), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n722), .B(KEYINPUT30), .C1(new_n635), .C2(new_n636), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT94), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n594), .A2(new_n596), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT94), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT30), .A4(new_n722), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n722), .B1(new_n635), .B2(new_n636), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT95), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n472), .A2(new_n325), .A3(new_n575), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT93), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n493), .B2(new_n542), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n599), .B1(KEYINPUT93), .B2(new_n733), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT30), .B1(new_n725), .B2(new_n722), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT95), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n728), .A2(new_n732), .A3(new_n737), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n677), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n721), .A2(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n724), .A2(new_n727), .B1(new_n735), .B2(new_n736), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n731), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n720), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(KEYINPUT98), .B1(new_n719), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n719), .A2(KEYINPUT98), .A3(new_n748), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(new_n221), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n233), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G41), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n562), .A2(G116), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(G1), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(new_n228), .B2(new_n755), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT92), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n752), .A2(new_n760), .ZN(G364));
  AOI21_X1  g0561(.A(new_n221), .B1(new_n670), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n754), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n684), .B2(G330), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G330), .B2(new_n684), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n229), .B1(G20), .B2(new_n328), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n222), .B1(new_n769), .B2(G190), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n263), .B1(new_n770), .B2(new_n509), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n222), .A2(new_n395), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n325), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n222), .A2(G190), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n769), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G322), .A2(new_n775), .B1(new_n778), .B2(G329), .ZN(new_n779));
  INV_X1    g0579(.A(G283), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n506), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n772), .A2(new_n781), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n779), .B1(new_n780), .B2(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT99), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(KEYINPUT99), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n787), .A2(G190), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n771), .B(new_n785), .C1(G326), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n773), .A2(new_n776), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n787), .A2(new_n395), .A3(new_n788), .ZN(new_n794));
  XOR2_X1   g0594(.A(KEYINPUT33), .B(G317), .Z(new_n795));
  OAI221_X1 g0595(.A(new_n791), .B1(new_n792), .B2(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n790), .A2(G50), .B1(new_n287), .B2(new_n775), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n387), .B2(new_n793), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT100), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n782), .A2(new_n251), .ZN(new_n800));
  INV_X1    g0600(.A(new_n784), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n263), .B(new_n800), .C1(G87), .C2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT101), .Z(new_n803));
  NOR2_X1   g0603(.A1(new_n770), .A2(new_n481), .ZN(new_n804));
  INV_X1    g0604(.A(new_n794), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(new_n805), .B2(G68), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n777), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n799), .A2(new_n803), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n768), .B1(new_n796), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G13), .A2(G33), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n767), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n259), .A2(G45), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n753), .A2(new_n300), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(G45), .C2(new_n228), .ZN(new_n818));
  INV_X1    g0618(.A(G355), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n233), .A2(new_n300), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(G116), .B2(new_n233), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n811), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n814), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n764), .B(new_n822), .C1(new_n684), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n766), .A2(new_n824), .ZN(G396));
  AND4_X1   g0625(.A1(new_n446), .A2(new_n447), .A3(new_n448), .A4(new_n678), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n446), .A2(new_n677), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n398), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n826), .B1(new_n449), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n666), .A2(new_n829), .A3(new_n678), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n706), .A2(new_n708), .ZN(new_n832));
  INV_X1    g0632(.A(new_n829), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n747), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT102), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n834), .A2(new_n747), .ZN(new_n838));
  INV_X1    g0638(.A(new_n764), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n834), .A2(KEYINPUT102), .A3(new_n747), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n793), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n790), .A2(G137), .B1(G159), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G143), .ZN(new_n844));
  INV_X1    g0644(.A(G150), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n843), .B1(new_n844), .B2(new_n774), .C1(new_n845), .C2(new_n794), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT34), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n300), .B1(new_n777), .B2(new_n848), .C1(new_n256), .C2(new_n784), .ZN(new_n849));
  INV_X1    g0649(.A(new_n770), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n287), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n847), .B(new_n851), .C1(new_n217), .C2(new_n782), .ZN(new_n852));
  INV_X1    g0652(.A(new_n782), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G116), .A2(new_n842), .B1(new_n853), .B2(G87), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n854), .B1(new_n251), .B2(new_n784), .C1(new_n509), .C2(new_n774), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n263), .B1(new_n777), .B2(new_n792), .C1(new_n794), .C2(new_n780), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n789), .A2(new_n783), .ZN(new_n857));
  OR4_X1    g0657(.A1(new_n804), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n768), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n767), .A2(new_n812), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n387), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n861), .B(new_n764), .C1(new_n829), .C2(new_n813), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n841), .A2(new_n862), .ZN(G384));
  INV_X1    g0663(.A(new_n674), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n298), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n334), .B2(new_n343), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g0667(.A(KEYINPUT105), .B(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n330), .A2(new_n865), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n340), .A2(new_n341), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n872));
  INV_X1    g0672(.A(new_n868), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n872), .A2(new_n330), .A3(new_n865), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n871), .A4(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n865), .B2(KEYINPUT106), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n877), .A2(new_n872), .A3(new_n330), .A4(new_n865), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT106), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n298), .B2(new_n864), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n869), .A2(new_n870), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n343), .A2(KEYINPUT107), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT107), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n339), .A2(new_n884), .A3(new_n342), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(new_n334), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n865), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n875), .B1(new_n888), .B2(KEYINPUT38), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n738), .B(KEYINPUT95), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n678), .B1(new_n890), .B2(new_n744), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT108), .B1(new_n891), .B2(KEYINPUT31), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n741), .A2(KEYINPUT108), .A3(KEYINPUT31), .A4(new_n677), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n743), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g0695(.A(KEYINPUT14), .B(new_n328), .C1(new_n365), .C2(new_n368), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n402), .A2(new_n896), .A3(new_n404), .ZN(new_n897));
  INV_X1    g0697(.A(new_n354), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT104), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT104), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n407), .A2(new_n900), .A3(new_n354), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n354), .A2(new_n677), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n372), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n408), .A2(new_n678), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n889), .A2(new_n895), .A3(new_n829), .A4(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT108), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n911), .A2(new_n893), .B1(new_n721), .B2(new_n742), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n373), .B1(new_n899), .B2(new_n901), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n905), .B1(new_n913), .B2(new_n903), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n912), .A2(new_n914), .A3(new_n833), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n871), .A2(new_n874), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(new_n866), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT40), .B1(new_n875), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(KEYINPUT40), .A2(new_n908), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n451), .A2(new_n912), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n920), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(G330), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n826), .A2(KEYINPUT103), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n826), .A2(KEYINPUT103), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n830), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n875), .A2(new_n918), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(new_n907), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n334), .B2(new_n864), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n902), .A2(new_n677), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n927), .A2(KEYINPUT39), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n875), .B(new_n933), .C1(new_n888), .C2(KEYINPUT38), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n923), .B(new_n936), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n710), .A2(new_n450), .A3(new_n716), .A4(new_n718), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n646), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n221), .B2(new_n670), .ZN(new_n941));
  INV_X1    g0741(.A(new_n619), .ZN(new_n942));
  OAI211_X1 g0742(.A(G20), .B(new_n309), .C1(new_n942), .C2(KEYINPUT35), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n212), .B(new_n943), .C1(KEYINPUT35), .C2(new_n942), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT36), .Z(new_n945));
  NOR3_X1   g0745(.A1(new_n277), .A2(new_n387), .A3(new_n228), .ZN(new_n946));
  INV_X1    g0746(.A(new_n202), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n217), .ZN(new_n948));
  OAI211_X1 g0748(.A(G1), .B(new_n669), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n941), .A2(new_n945), .A3(new_n949), .ZN(G367));
  OAI21_X1  g0750(.A(new_n300), .B1(new_n782), .B2(new_n387), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT113), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n850), .A2(G68), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n775), .A2(G150), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n801), .A2(new_n287), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n842), .A2(new_n947), .ZN(new_n956));
  AND4_X1   g0756(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n778), .A2(G137), .ZN(new_n958));
  AOI22_X1  g0758(.A1(G143), .A2(new_n790), .B1(new_n805), .B2(G159), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n952), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT114), .Z(new_n961));
  NOR2_X1   g0761(.A1(new_n793), .A2(new_n780), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n263), .B1(new_n770), .B2(new_n251), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n774), .A2(new_n783), .B1(new_n782), .B2(new_n481), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(G317), .C2(new_n778), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G294), .A2(new_n805), .B1(new_n790), .B2(G311), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n801), .A2(G116), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n961), .B1(new_n962), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n839), .B1(new_n971), .B2(new_n767), .ZN(new_n972));
  INV_X1    g0772(.A(new_n817), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n815), .B1(new_n233), .B2(new_n380), .C1(new_n247), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n579), .A2(new_n677), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n653), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n704), .B2(new_n975), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n972), .B(new_n974), .C1(new_n823), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n632), .A2(new_n677), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n647), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n638), .A2(new_n626), .ZN(new_n981));
  INV_X1    g0781(.A(new_n979), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n691), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT42), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n626), .B1(new_n983), .B2(new_n546), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n678), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT109), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT109), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n985), .A2(new_n990), .A3(new_n987), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n977), .B(KEYINPUT43), .Z(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n989), .B2(new_n991), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n689), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(new_n983), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n997), .B(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n692), .A2(new_n983), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n692), .A2(new_n983), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  AND4_X1   g0806(.A1(KEYINPUT110), .A2(new_n1003), .A3(new_n689), .A4(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1003), .A2(new_n1006), .B1(new_n689), .B2(KEYINPUT110), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n684), .A2(G330), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT112), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT112), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n684), .A2(new_n1012), .A3(G330), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT111), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n691), .A2(new_n1014), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n688), .A2(new_n690), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1011), .A2(new_n1013), .A3(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1013), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n751), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1009), .A2(new_n1022), .B1(new_n1023), .B2(new_n749), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n754), .B(KEYINPUT41), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n763), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n978), .B1(new_n1001), .B2(new_n1026), .ZN(G387));
  OAI21_X1  g0827(.A(new_n1021), .B1(new_n1023), .B2(new_n749), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n750), .A2(new_n751), .A3(new_n1022), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n1029), .A3(new_n754), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n817), .B1(new_n243), .B2(new_n459), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n383), .A2(new_n256), .ZN(new_n1032));
  AOI211_X1 g0832(.A(G116), .B(new_n562), .C1(new_n1032), .C2(KEYINPUT50), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n459), .C1(KEYINPUT50), .C2(new_n1032), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G68), .B2(G77), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n820), .A2(new_n756), .B1(G107), .B2(new_n233), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT115), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n815), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n764), .C1(new_n688), .C2(new_n823), .ZN(new_n1040));
  INV_X1    g0840(.A(G322), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n792), .A2(new_n794), .B1(new_n789), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT116), .ZN(new_n1043));
  INV_X1    g0843(.A(G317), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n783), .B2(new_n793), .C1(new_n1044), .C2(new_n774), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT48), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n780), .B2(new_n770), .C1(new_n509), .C2(new_n784), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n778), .A2(G326), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n300), .B1(new_n853), .B2(G116), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n793), .A2(new_n217), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n300), .B1(new_n782), .B2(new_n481), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n256), .A2(new_n774), .B1(new_n784), .B2(new_n387), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G150), .C2(new_n778), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n288), .A2(new_n805), .B1(new_n790), .B2(G159), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n381), .A2(new_n850), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1053), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1040), .B1(new_n1061), .B2(new_n767), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n1021), .B2(new_n763), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1030), .A2(new_n1063), .ZN(G393));
  OAI221_X1 g0864(.A(new_n1021), .B1(new_n1008), .B2(new_n1007), .C1(new_n1023), .C2(new_n749), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1028), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(new_n998), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1065), .B(new_n754), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n983), .A2(new_n814), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n770), .A2(new_n387), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n263), .B1(new_n853), .B2(G87), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n217), .B2(new_n784), .C1(new_n844), .C2(new_n777), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT118), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1071), .B(new_n1074), .C1(new_n947), .C2(new_n805), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n842), .A2(new_n383), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n790), .A2(G150), .B1(G159), .B2(new_n775), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1075), .A2(new_n1076), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n263), .B1(new_n212), .B2(new_n770), .C1(new_n794), .C2(new_n783), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n789), .A2(new_n1044), .B1(new_n792), .B2(new_n774), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n784), .A2(new_n780), .B1(new_n777), .B2(new_n1041), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n800), .B(new_n1085), .C1(G294), .C2(new_n842), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1081), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n767), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1070), .A2(new_n1089), .A3(new_n764), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n253), .A2(new_n817), .B1(G97), .B2(new_n753), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n815), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1068), .B2(new_n763), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1069), .A2(new_n1093), .ZN(G390));
  NAND2_X1  g0894(.A1(new_n828), .A2(new_n449), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n678), .B(new_n1095), .C1(new_n713), .C2(new_n715), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n826), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n889), .B(new_n931), .C1(new_n1098), .C2(new_n914), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n932), .A2(new_n934), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n930), .B1(new_n926), .B2(new_n907), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n895), .A2(new_n907), .A3(G330), .A4(new_n829), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n981), .A2(new_n540), .A3(new_n583), .A4(new_n678), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n891), .B1(KEYINPUT31), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n746), .ZN(new_n1107));
  OAI211_X1 g0907(.A(G330), .B(new_n829), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(new_n914), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1099), .B(new_n1109), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n926), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n914), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n1103), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT119), .B1(new_n912), .B2(new_n720), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT119), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n895), .A2(new_n1115), .A3(G330), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n1116), .A3(new_n829), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n914), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1098), .B1(new_n1108), .B2(new_n914), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1113), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n921), .A2(G330), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n938), .A2(new_n646), .A3(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1104), .B(new_n1110), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n911), .A2(new_n893), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n720), .B1(new_n1126), .B2(new_n743), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n833), .B1(new_n1127), .B2(new_n1115), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n907), .B1(new_n1128), .B2(new_n1114), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1112), .A2(new_n1103), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1129), .A2(new_n1119), .B1(new_n1111), .B2(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n938), .A2(new_n646), .A3(new_n1122), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1125), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1124), .A2(new_n1133), .A3(new_n754), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n782), .A2(new_n217), .B1(new_n777), .B2(new_n509), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT121), .Z(new_n1136));
  NAND2_X1  g0936(.A1(new_n775), .A2(G116), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G107), .A2(new_n805), .B1(new_n790), .B2(G283), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n263), .B1(new_n784), .B2(new_n561), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1071), .B(new_n1139), .C1(G97), .C2(new_n842), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT53), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n801), .A2(new_n1142), .A3(G150), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1143), .B1(new_n807), .B2(new_n770), .C1(new_n1144), .C2(new_n789), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G137), .B2(new_n805), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT54), .B(G143), .Z(new_n1147));
  NAND2_X1  g0947(.A1(new_n842), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n300), .B1(new_n782), .B2(new_n202), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT120), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(G125), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n774), .A2(new_n848), .B1(new_n777), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n1150), .B2(new_n1149), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1146), .A2(new_n1148), .A3(new_n1151), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1142), .B1(new_n801), .B2(G150), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1141), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1157), .A2(new_n767), .B1(new_n289), .B2(new_n860), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n764), .B(new_n1158), .C1(new_n1100), .C2(new_n813), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1125), .B2(new_n763), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1134), .A2(new_n1161), .ZN(G378));
  INV_X1    g0962(.A(KEYINPUT123), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n645), .A2(new_n433), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT122), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT122), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n445), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n431), .A2(new_n864), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1169), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1167), .B1(new_n645), .B2(new_n433), .ZN(new_n1172));
  AOI211_X1 g0972(.A(KEYINPUT122), .B(new_n434), .C1(new_n441), .C2(new_n444), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1164), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1170), .A2(new_n1174), .A3(new_n1164), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1163), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n920), .B2(new_n720), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1170), .A2(new_n1174), .A3(new_n1164), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT123), .B1(new_n1180), .B2(new_n1175), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT40), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n915), .B2(new_n889), .ZN(new_n1183));
  AND4_X1   g0983(.A1(new_n829), .A2(new_n919), .A3(new_n895), .A4(new_n907), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1181), .B(G330), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1179), .A2(new_n936), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n936), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n763), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n801), .A2(new_n1147), .B1(new_n842), .B2(G137), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n1152), .B2(new_n789), .C1(new_n845), .C2(new_n770), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G132), .B2(new_n805), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1144), .B2(new_n774), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT59), .Z(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(new_n266), .C1(new_n807), .C2(new_n782), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G41), .B(new_n1194), .C1(G124), .C2(new_n778), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G50), .B1(new_n268), .B2(new_n454), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n454), .B(new_n263), .C1(new_n784), .C2(new_n387), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n775), .A2(G107), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n853), .A2(new_n287), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n778), .A2(G283), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n953), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1197), .B(new_n1201), .C1(new_n381), .C2(new_n842), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n481), .B2(new_n794), .C1(new_n212), .C2(new_n789), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT58), .Z(new_n1204));
  NOR3_X1   g1004(.A1(new_n1195), .A2(new_n1196), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n764), .B1(new_n1205), .B2(new_n768), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n860), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1180), .A2(new_n1175), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1207), .B1(new_n947), .B2(new_n1208), .C1(new_n1209), .C2(new_n813), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1188), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1123), .A2(KEYINPUT124), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT124), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n938), .A2(new_n1214), .A3(new_n646), .A4(new_n1122), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1179), .A2(new_n1185), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n936), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1179), .A2(new_n936), .A3(new_n1185), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1217), .A2(new_n1133), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n754), .B1(new_n1222), .B2(KEYINPUT57), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1125), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n1224), .A2(new_n1216), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1212), .B1(new_n1223), .B2(new_n1227), .ZN(G375));
  NOR2_X1   g1028(.A1(new_n770), .A2(new_n256), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G137), .A2(new_n775), .B1(new_n842), .B2(G150), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n1144), .B2(new_n777), .C1(new_n807), .C2(new_n784), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1229), .B(new_n1231), .C1(new_n805), .C2(new_n1147), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n790), .A2(G132), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT125), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1232), .A2(new_n300), .A3(new_n1199), .A4(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n784), .A2(new_n481), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n774), .A2(new_n780), .B1(new_n777), .B2(new_n783), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G107), .B2(new_n842), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G116), .A2(new_n805), .B1(new_n790), .B2(G294), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n300), .B1(new_n853), .B2(G77), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1059), .A4(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1235), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n767), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(G68), .B2(new_n1208), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n839), .B(new_n1244), .C1(new_n914), .C2(new_n812), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1131), .B2(new_n763), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1025), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1248), .B2(new_n1249), .ZN(G381));
  AOI21_X1  g1050(.A(new_n755), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1222), .A2(KEYINPUT57), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1211), .A2(G378), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(G387), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1257));
  INV_X1    g1057(.A(G396), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1030), .A2(new_n1258), .A3(new_n1063), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1256), .A2(new_n1257), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT126), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1256), .A2(KEYINPUT126), .A3(new_n1257), .A4(new_n1260), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(G407));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(new_n675), .C2(new_n1255), .ZN(G409));
  AND2_X1   g1066(.A1(new_n676), .A2(G213), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1222), .A2(new_n1025), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1254), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1211), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1270));
  INV_X1    g1070(.A(G378), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n1123), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1276), .A2(new_n754), .A3(new_n1247), .A4(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1278), .A2(G384), .A3(new_n1246), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1278), .B2(new_n1246), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1274), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1246), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1278), .A2(G384), .A3(new_n1246), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(new_n1285), .A3(new_n1273), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1281), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT61), .B1(new_n1272), .B2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1269), .B(new_n1289), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT62), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G375), .A2(G378), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1292), .A2(new_n1293), .A3(new_n1269), .A4(new_n1289), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1288), .A2(new_n1291), .A3(new_n1294), .ZN(new_n1295));
  OR2_X1    g1095(.A1(G387), .A2(G390), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(G390), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1258), .B1(new_n1030), .B2(new_n1063), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1299), .A2(KEYINPUT127), .A3(new_n1259), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT127), .B1(new_n1299), .B2(new_n1259), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1296), .B(new_n1297), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1299), .A2(KEYINPUT127), .A3(new_n1259), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1297), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(G387), .A2(G390), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1295), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1269), .A4(new_n1289), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1290), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(new_n1272), .B2(new_n1287), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1310), .B(new_n1311), .C1(new_n1312), .C2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1309), .A2(new_n1315), .ZN(G405));
  NOR2_X1   g1116(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1289), .B1(new_n1256), .B2(new_n1317), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1292), .B(new_n1255), .C1(new_n1280), .C2(new_n1279), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1307), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1308), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(G402));
endmodule


