//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1202, new_n1203, new_n1204, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G257), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G77), .B2(G244), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n212), .A2(new_n213), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n205), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(new_n202), .A2(G50), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT64), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G250), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n205), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n231), .B(new_n233), .C1(new_n208), .C2(new_n210), .ZN(new_n234));
  AOI22_X1  g0034(.A1(new_n227), .A2(new_n230), .B1(new_n234), .B2(KEYINPUT0), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n225), .B(new_n235), .C1(KEYINPUT0), .C2(new_n234), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n215), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n222), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT66), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G50), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G107), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n221), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT67), .B(G45), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n255), .B(G274), .C1(new_n257), .C2(G41), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G226), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G222), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(new_n265), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(new_n266), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n270), .B1(G223), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n259), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n258), .B(new_n264), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n279), .A2(G179), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G50), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n228), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n255), .A2(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n214), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT68), .A2(G58), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT68), .A2(G58), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT8), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OR3_X1    g0091(.A1(new_n247), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT69), .B1(new_n247), .B2(KEYINPUT8), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n273), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n297));
  INV_X1    g0097(.A(G150), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n229), .A2(new_n273), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AOI211_X1 g0100(.A(new_n282), .B(new_n288), .C1(new_n300), .C2(new_n284), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n279), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n280), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n301), .A2(KEYINPUT9), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n301), .A2(KEYINPUT9), .B1(new_n279), .B2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n279), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n265), .A2(G232), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n314), .B1(new_n267), .B2(new_n215), .C1(new_n266), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n259), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n263), .A2(G238), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n258), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT70), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT13), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n317), .A2(new_n322), .A3(new_n258), .A4(new_n318), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(G169), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT14), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n320), .A2(G179), .A3(new_n323), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n324), .A2(new_n329), .A3(G169), .A4(new_n325), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n287), .A2(new_n216), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G20), .A2(G33), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n295), .A2(G77), .B1(new_n333), .B2(G50), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n229), .B2(G68), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n335), .A2(new_n284), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n336), .B2(KEYINPUT11), .ZN(new_n337));
  INV_X1    g0137(.A(new_n281), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n216), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT12), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n337), .B(new_n340), .C1(KEYINPUT11), .C2(new_n336), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT71), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n331), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n324), .A2(G200), .A3(new_n325), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n320), .A2(G190), .A3(new_n323), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n265), .A2(G1698), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n348), .A2(new_n217), .B1(new_n209), .B2(new_n265), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n315), .A2(G1698), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n259), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n263), .A2(G244), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n258), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT15), .B(G87), .Z(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n295), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT8), .B(G58), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n358), .B1(new_n229), .B2(new_n269), .C1(new_n299), .C2(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n284), .B1(new_n269), .B2(new_n338), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n269), .B2(new_n287), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n353), .A2(new_n303), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n356), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n313), .A2(new_n344), .A3(new_n347), .A4(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT73), .B1(new_n273), .B2(KEYINPUT3), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT73), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(new_n271), .A3(G33), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n369), .A3(new_n274), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(G20), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n371), .B1(new_n265), .B2(G20), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n216), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G159), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT72), .B1(new_n299), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT72), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n333), .A2(new_n378), .A3(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n289), .A2(new_n290), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n201), .B1(new_n381), .B2(G68), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n380), .B1(new_n382), .B2(new_n229), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n366), .B1(new_n375), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT74), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(KEYINPUT74), .B(new_n366), .C1(new_n375), .C2(new_n383), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n275), .A2(new_n372), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n216), .B1(new_n374), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n285), .B1(new_n392), .B2(KEYINPUT16), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n389), .B1(new_n388), .B2(new_n393), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n294), .A2(new_n286), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT76), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n338), .A2(new_n284), .ZN(new_n398));
  INV_X1    g0198(.A(new_n294), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n397), .A2(new_n398), .B1(new_n338), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n394), .A2(new_n395), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n265), .A2(G223), .A3(new_n266), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n348), .C2(new_n215), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT77), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n276), .A2(G226), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT77), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n403), .A3(new_n408), .A4(new_n404), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(new_n409), .A3(new_n259), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n263), .A2(G232), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n258), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G200), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(new_n308), .A3(new_n412), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n402), .A2(KEYINPUT78), .A3(KEYINPUT17), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  OR2_X1    g0219(.A1(KEYINPUT68), .A2(G58), .ZN(new_n420));
  NAND2_X1  g0220(.A1(KEYINPUT68), .A2(G58), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(G68), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n202), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G20), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n275), .A2(new_n229), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n371), .B1(new_n370), .B2(new_n372), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n424), .B(new_n380), .C1(new_n426), .C2(new_n216), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT74), .B1(new_n427), .B2(new_n366), .ZN(new_n428));
  INV_X1    g0228(.A(new_n387), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n393), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(new_n400), .A3(new_n417), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT78), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n419), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(new_n400), .A3(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n413), .A2(G169), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n355), .B2(new_n413), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n436), .A2(KEYINPUT18), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT18), .B1(new_n436), .B2(new_n438), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n418), .B(new_n435), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n362), .B1(G200), .B2(new_n353), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n354), .A2(G190), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n365), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n285), .B(new_n281), .C1(G1), .C2(new_n273), .ZN(new_n448));
  OR3_X1    g0248(.A1(new_n448), .A2(KEYINPUT85), .A3(new_n221), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT85), .B1(new_n448), .B2(new_n221), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n229), .C1(G33), .C2(new_n207), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(new_n284), .C1(new_n229), .C2(G116), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n455), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n456), .A2(new_n457), .B1(new_n221), .B2(new_n338), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n303), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n255), .A2(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n462));
  AND2_X1   g0262(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n260), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT80), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(KEYINPUT80), .B(new_n260), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  AOI211_X1 g0268(.A(new_n461), .B(new_n462), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n469), .A2(new_n222), .A3(new_n259), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n265), .A2(G257), .A3(new_n266), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n275), .A2(G303), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n348), .C2(new_n210), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n259), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n467), .A2(new_n468), .ZN(new_n475));
  INV_X1    g0275(.A(new_n461), .ZN(new_n476));
  INV_X1    g0276(.A(G274), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n259), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n462), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n475), .A2(new_n476), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT84), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n470), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n469), .A2(new_n478), .B1(new_n259), .B2(new_n473), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G270), .A3(new_n278), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT84), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n459), .B(new_n460), .C1(new_n483), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n482), .B1(new_n470), .B2(new_n481), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n484), .A2(KEYINPUT84), .A3(new_n486), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(KEYINPUT86), .A3(KEYINPUT21), .A4(new_n459), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n451), .A2(new_n458), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n484), .A2(G179), .A3(new_n486), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT87), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n470), .A2(new_n481), .A3(new_n355), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT87), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n500), .A3(new_n495), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n490), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(KEYINPUT88), .B(new_n495), .C1(new_n493), .C2(G200), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT88), .ZN(new_n505));
  OAI21_X1  g0305(.A(G200), .B1(new_n483), .B2(new_n487), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(new_n496), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n493), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G190), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n503), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n485), .A2(G257), .A3(new_n278), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT81), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n272), .A2(new_n274), .A3(G244), .A4(new_n266), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n452), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n469), .A2(new_n478), .B1(new_n519), .B2(new_n259), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT81), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n485), .A2(new_n521), .A3(G257), .A4(new_n278), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n513), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G200), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT82), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n513), .A2(G190), .A3(new_n520), .A4(new_n522), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n281), .A2(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n448), .A2(new_n207), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n207), .A2(new_n209), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n530), .B1(new_n533), .B2(KEYINPUT6), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G20), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n299), .A2(new_n269), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n537), .C1(new_n426), .C2(new_n209), .ZN(new_n538));
  AOI211_X1 g0338(.A(new_n528), .B(new_n529), .C1(new_n538), .C2(new_n284), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n527), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n523), .A2(KEYINPUT82), .A3(G200), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n526), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n523), .A2(G169), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n513), .A2(G179), .A3(new_n520), .A4(new_n522), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n539), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  INV_X1    g0348(.A(G244), .ZN(new_n549));
  OAI221_X1 g0349(.A(new_n548), .B1(new_n348), .B2(new_n549), .C1(new_n217), .C2(new_n267), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n259), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n461), .A2(new_n477), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n278), .A2(G250), .A3(new_n461), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(new_n355), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n265), .A2(new_n229), .A3(G68), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n229), .B1(new_n314), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n532), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n557), .B1(new_n314), .B2(G20), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n556), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n284), .ZN(new_n564));
  INV_X1    g0364(.A(new_n357), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n338), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n566), .C1(new_n565), .C2(new_n448), .ZN(new_n567));
  INV_X1    g0367(.A(new_n554), .ZN(new_n568));
  AOI211_X1 g0368(.A(new_n552), .B(new_n568), .C1(new_n550), .C2(new_n259), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n555), .B(new_n567), .C1(new_n569), .C2(G169), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n551), .A2(G190), .A3(new_n553), .A4(new_n554), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n448), .A2(new_n559), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n572), .A2(new_n566), .A3(new_n564), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n573), .C1(new_n569), .C2(new_n414), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT83), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n542), .A2(new_n547), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n542), .A2(new_n575), .A3(new_n547), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT83), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n265), .A2(new_n229), .A3(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT89), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT89), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n265), .A2(new_n582), .A3(new_n229), .A4(G87), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(KEYINPUT22), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n229), .A2(G107), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n585), .B(KEYINPUT23), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT22), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n580), .A2(KEYINPUT89), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n295), .A2(G116), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n584), .A2(new_n586), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT24), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n588), .A2(new_n589), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n586), .A4(new_n584), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n284), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n448), .A2(new_n209), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n338), .A2(new_n209), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n599), .B(KEYINPUT25), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n596), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n485), .A2(G264), .A3(new_n278), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n231), .A2(new_n267), .B1(new_n348), .B2(new_n208), .ZN(new_n604));
  INV_X1    g0404(.A(G294), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n273), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n259), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n607), .A3(new_n480), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n414), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n603), .A2(new_n607), .A3(new_n308), .A4(new_n480), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT90), .B1(new_n602), .B2(new_n612), .ZN(new_n613));
  AOI211_X1 g0413(.A(new_n597), .B(new_n600), .C1(new_n595), .C2(new_n284), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT90), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n611), .ZN(new_n616));
  INV_X1    g0416(.A(new_n608), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(G169), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n355), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n613), .A2(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n511), .A2(new_n577), .A3(new_n579), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n447), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n618), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n602), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n625), .A2(new_n494), .A3(new_n490), .A4(new_n502), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n542), .A2(new_n547), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n613), .A2(new_n616), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n575), .A4(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n575), .A2(new_n545), .A3(new_n546), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT26), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n545), .B(KEYINPUT91), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(new_n575), .A4(new_n546), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n629), .A2(new_n570), .A3(new_n631), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n446), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n440), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n436), .A2(KEYINPUT18), .A3(new_n438), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n418), .A2(new_n435), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n364), .A2(KEYINPUT92), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n364), .A2(KEYINPUT92), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n331), .A2(new_n343), .B1(new_n347), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n639), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n311), .A2(new_n312), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n305), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n636), .A2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(G13), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(G20), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n255), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n496), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n511), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n503), .A2(new_n659), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n628), .B(new_n625), .C1(new_n614), .C2(new_n658), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT93), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n619), .A2(new_n665), .A3(new_n620), .A4(new_n657), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT93), .B1(new_n625), .B2(new_n658), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n663), .A2(G330), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n625), .A2(new_n657), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n503), .A2(new_n658), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT94), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n673), .B2(new_n669), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(G399));
  NOR2_X1   g0475(.A1(new_n233), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n560), .A2(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n227), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n677), .ZN(new_n681));
  XOR2_X1   g0481(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n682));
  XNOR2_X1  g0482(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n569), .A2(new_n603), .A3(new_n607), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n684), .A2(new_n523), .A3(new_n497), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT30), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n523), .A2(new_n355), .ZN(new_n687));
  NOR4_X1   g0487(.A1(new_n509), .A2(new_n687), .A3(new_n569), .A4(new_n617), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n657), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI211_X1 g0489(.A(KEYINPUT31), .B(new_n689), .C1(new_n622), .C2(new_n657), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n689), .A2(KEYINPUT31), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n629), .A2(new_n570), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT97), .ZN(new_n694));
  INV_X1    g0494(.A(new_n630), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(KEYINPUT26), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n630), .A2(KEYINPUT97), .A3(new_n633), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n632), .A2(new_n575), .A3(new_n546), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n633), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n657), .B1(new_n693), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n635), .A2(new_n658), .ZN(new_n702));
  XNOR2_X1  g0502(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI22_X1  g0504(.A1(G330), .A2(new_n692), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n683), .B1(new_n705), .B2(G1), .ZN(G364));
  NAND2_X1  g0506(.A1(new_n663), .A2(G330), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n651), .A2(G45), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n677), .A2(G1), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n661), .A2(new_n710), .A3(new_n662), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n709), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n228), .B1(G20), .B2(new_n303), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n229), .A2(G190), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n355), .A2(G200), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G311), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n275), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n355), .A2(new_n414), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n716), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G317), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT33), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(KEYINPUT33), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n229), .A2(new_n308), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n717), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G322), .ZN(new_n731));
  INV_X1    g0531(.A(G283), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n414), .A2(G179), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n716), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n727), .B(new_n731), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G179), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n716), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT102), .Z(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n720), .B(new_n735), .C1(G329), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n721), .A2(new_n728), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT100), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n741), .A2(new_n742), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n229), .B1(new_n736), .B2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n747), .A2(G326), .B1(G294), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT101), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n740), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G303), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n728), .A2(new_n733), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n752), .B1(KEYINPUT101), .B2(new_n750), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n737), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G159), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n757), .A2(KEYINPUT32), .B1(new_n207), .B2(new_n748), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n275), .B(new_n758), .C1(KEYINPUT32), .C2(new_n757), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n723), .A2(G68), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n729), .B(KEYINPUT99), .ZN(new_n761));
  INV_X1    g0561(.A(new_n734), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n761), .A2(new_n381), .B1(G107), .B2(new_n762), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n754), .A2(new_n559), .B1(new_n718), .B2(new_n269), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n747), .B2(G50), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n759), .A2(new_n760), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n715), .B1(new_n755), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n233), .A2(new_n265), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n768), .B1(new_n680), .B2(new_n257), .C1(new_n250), .C2(new_n261), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n265), .A2(new_n232), .ZN(new_n770));
  XOR2_X1   g0570(.A(G355), .B(KEYINPUT98), .Z(new_n771));
  OAI221_X1 g0571(.A(new_n769), .B1(G116), .B2(new_n232), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n714), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n767), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n775), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n713), .B(new_n777), .C1(new_n663), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n712), .A2(new_n779), .ZN(G396));
  NAND2_X1  g0580(.A1(new_n692), .A2(G330), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n362), .A2(new_n657), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT104), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n364), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n356), .A2(KEYINPUT104), .A3(new_n362), .A4(new_n363), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT105), .ZN(new_n788));
  AND3_X1   g0588(.A1(new_n787), .A2(new_n788), .A3(new_n444), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(new_n787), .B2(new_n444), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n782), .B1(new_n642), .B2(new_n643), .ZN(new_n791));
  OR3_X1    g0591(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n702), .B(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n781), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n709), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT103), .B(G283), .ZN(new_n796));
  INV_X1    g0596(.A(new_n754), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n723), .A2(new_n796), .B1(new_n797), .B2(G107), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n798), .B1(new_n221), .B2(new_n718), .C1(new_n605), .C2(new_n729), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n734), .A2(new_n559), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n799), .A2(new_n265), .A3(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G303), .A2(new_n747), .B1(new_n739), .B2(G311), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(new_n207), .C2(new_n748), .ZN(new_n803));
  INV_X1    g0603(.A(new_n718), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n747), .A2(G137), .B1(G159), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G143), .ZN(new_n806));
  INV_X1    g0606(.A(new_n761), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(new_n806), .B2(new_n807), .C1(new_n298), .C2(new_n722), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT34), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G68), .A2(new_n762), .B1(new_n749), .B2(new_n381), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n265), .B1(new_n214), .B2(new_n754), .C1(new_n738), .C2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n803), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n714), .A2(new_n773), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n814), .A2(new_n714), .B1(new_n269), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n816), .B(new_n713), .C1(new_n792), .C2(new_n774), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n795), .A2(new_n817), .ZN(G384));
  AOI21_X1  g0618(.A(new_n221), .B1(new_n534), .B2(KEYINPUT35), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(new_n230), .C1(KEYINPUT35), .C2(new_n534), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT36), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n227), .A2(G77), .A3(new_n422), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(G50), .B2(new_n216), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n823), .A2(G1), .A3(new_n650), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n651), .A2(new_n255), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT108), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n344), .A2(new_n657), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n402), .A2(new_n655), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n441), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n655), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n436), .B1(new_n438), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n433), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT37), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(new_n838), .A3(new_n433), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n830), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n393), .B1(KEYINPUT16), .B2(new_n392), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n400), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n438), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n833), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT37), .B1(new_n836), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n846), .ZN(new_n849));
  AOI221_X4 g0649(.A(new_n842), .B1(new_n848), .B2(new_n839), .C1(new_n441), .C2(new_n849), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n841), .A2(new_n850), .A3(KEYINPUT39), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n846), .B1(new_n640), .B2(new_n639), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n839), .A2(new_n848), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n842), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n441), .A2(new_n849), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(KEYINPUT38), .A3(new_n854), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n852), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT106), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n857), .B2(new_n854), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT39), .B1(new_n850), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT106), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n828), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n639), .A2(new_n833), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n344), .B(new_n347), .C1(new_n342), .C2(new_n658), .ZN(new_n867));
  INV_X1    g0667(.A(new_n347), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n343), .B(new_n657), .C1(new_n331), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n635), .A2(new_n658), .A3(new_n792), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n785), .A2(new_n786), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n873), .A2(new_n657), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n871), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n856), .A2(new_n858), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n866), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n826), .B1(new_n865), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n441), .A2(new_n831), .B1(new_n837), .B2(new_n839), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n858), .B(new_n852), .C1(new_n881), .C2(new_n830), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n863), .B1(new_n862), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT106), .B1(new_n877), .B2(KEYINPUT39), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n827), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(KEYINPUT108), .A3(new_n878), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n701), .A2(new_n446), .A3(new_n704), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n648), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT109), .Z(new_n890));
  XNOR2_X1  g0690(.A(new_n887), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n858), .B1(new_n881), .B2(new_n830), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n867), .B2(new_n869), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n892), .A2(new_n690), .A3(new_n691), .A4(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n690), .A2(new_n894), .A3(new_n691), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT40), .B1(new_n856), .B2(new_n858), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n895), .A2(KEYINPUT40), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n692), .A2(new_n446), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n898), .B(new_n899), .Z(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n710), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n825), .B1(new_n891), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT110), .Z(new_n903));
  NOR2_X1   g0703(.A1(new_n891), .A2(new_n901), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n821), .B(new_n824), .C1(new_n903), .C2(new_n904), .ZN(G367));
  INV_X1    g0705(.A(new_n768), .ZN(new_n906));
  OAI221_X1 g0706(.A(new_n776), .B1(new_n232), .B2(new_n565), .C1(new_n244), .C2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n575), .B1(new_n573), .B2(new_n658), .ZN(new_n908));
  OR3_X1    g0708(.A1(new_n570), .A2(new_n573), .A3(new_n658), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n713), .B(new_n907), .C1(new_n910), .C2(new_n778), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n797), .A2(KEYINPUT46), .A3(G116), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(KEYINPUT113), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(KEYINPUT113), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT114), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT46), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n754), .B2(new_n221), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n913), .B(new_n918), .C1(G311), .C2(new_n747), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n804), .A2(new_n796), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n761), .A2(G303), .B1(new_n915), .B2(new_n917), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n722), .A2(new_n605), .B1(new_n737), .B2(new_n724), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n275), .B1(new_n748), .B2(new_n209), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n734), .A2(new_n207), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n749), .A2(G68), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n298), .B2(new_n729), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT115), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT115), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n929), .B(new_n930), .C1(new_n806), .C2(new_n746), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT116), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n762), .A2(G77), .ZN(new_n935));
  INV_X1    g0735(.A(G137), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n935), .B1(new_n214), .B2(new_n718), .C1(new_n936), .C2(new_n737), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n275), .B(new_n937), .C1(new_n381), .C2(new_n797), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n933), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n722), .A2(new_n376), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n926), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT47), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n911), .B1(new_n714), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT117), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n627), .B1(new_n539), .B2(new_n658), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n632), .A2(new_n546), .A3(new_n657), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n673), .A2(new_n669), .A3(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT42), .Z(new_n951));
  INV_X1    g0751(.A(new_n949), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n547), .B1(new_n952), .B2(new_n625), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n658), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n946), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n670), .A2(new_n952), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n955), .A2(new_n946), .A3(new_n956), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n708), .A2(G1), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT111), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n674), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n673), .A2(new_n669), .ZN(new_n968));
  INV_X1    g0768(.A(new_n671), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n967), .B1(new_n970), .B2(new_n952), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(KEYINPUT44), .A3(new_n952), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT44), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n674), .B2(new_n949), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n966), .A2(new_n971), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n965), .B1(new_n975), .B2(new_n670), .ZN(new_n976));
  INV_X1    g0776(.A(new_n673), .ZN(new_n977));
  INV_X1    g0777(.A(new_n670), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n669), .B1(new_n663), .B2(G330), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n979), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n670), .A3(new_n673), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(KEYINPUT112), .A3(new_n705), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT112), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n701), .A2(new_n704), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n781), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n980), .A2(new_n982), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n976), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n971), .A2(new_n966), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n972), .A2(new_n974), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n978), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n975), .A2(new_n670), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n965), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n705), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n676), .B(KEYINPUT41), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n964), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n944), .B1(new_n963), .B2(new_n999), .ZN(G387));
  NAND2_X1  g0800(.A1(new_n984), .A2(new_n989), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n676), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT119), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n987), .A2(new_n988), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1001), .A2(KEYINPUT119), .A3(new_n676), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n983), .A2(new_n964), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n747), .A2(G322), .B1(G303), .B2(new_n804), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n719), .B2(new_n722), .C1(new_n724), .C2(new_n807), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT48), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n605), .B2(new_n754), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n749), .B2(new_n796), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT49), .Z(new_n1014));
  AOI21_X1  g0814(.A(new_n265), .B1(new_n756), .B2(G326), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n221), .C2(new_n734), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G77), .A2(new_n797), .B1(new_n804), .B2(G68), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n214), .B2(new_n729), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n924), .B(new_n1018), .C1(G150), .C2(new_n756), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n747), .A2(G159), .B1(new_n294), .B2(new_n723), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n565), .C2(new_n748), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1016), .B1(new_n275), .B2(new_n1021), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n359), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT50), .B1(new_n359), .B2(G50), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1023), .A2(new_n261), .A3(new_n678), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n216), .A2(new_n269), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n768), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT118), .Z(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n241), .B2(new_n256), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(G107), .B2(new_n232), .C1(new_n678), .C2(new_n770), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1022), .A2(new_n714), .B1(new_n776), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(new_n713), .C1(new_n669), .C2(new_n778), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1007), .A2(new_n1008), .A3(new_n1032), .ZN(G393));
  NAND3_X1  g0833(.A1(new_n994), .A2(new_n995), .A3(new_n964), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n776), .B1(new_n207), .B2(new_n232), .C1(new_n253), .C2(new_n906), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n747), .A2(G150), .B1(G159), .B2(new_n730), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT51), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n748), .A2(new_n269), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1036), .A2(KEYINPUT51), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n756), .A2(G143), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n216), .B2(new_n754), .C1(new_n359), .C2(new_n718), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n800), .B(new_n1042), .C1(G50), .C2(new_n723), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n746), .A2(new_n724), .B1(new_n719), .B2(new_n729), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT52), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n797), .A2(new_n796), .B1(new_n756), .B2(G322), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT120), .Z(new_n1048));
  NOR2_X1   g0848(.A1(new_n718), .A2(new_n605), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n275), .B1(new_n734), .B2(new_n209), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G116), .C2(new_n749), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1046), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n722), .A2(new_n753), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1044), .A2(new_n275), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n709), .B1(new_n1054), .B2(new_n714), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1035), .B(new_n1055), .C1(new_n949), .C2(new_n778), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n676), .B1(new_n990), .B2(new_n996), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n989), .A2(new_n984), .B1(new_n994), .B2(new_n995), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1034), .B(new_n1056), .C1(new_n1057), .C2(new_n1058), .ZN(G390));
  NAND2_X1  g0859(.A1(new_n872), .A2(new_n875), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n690), .A2(G330), .A3(new_n691), .A4(new_n792), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1061), .A2(new_n871), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n871), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n692), .A2(G330), .A3(new_n792), .A4(new_n870), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n874), .B1(new_n700), .B2(new_n792), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1061), .A2(new_n871), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n692), .A2(G330), .A3(new_n446), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n888), .A3(new_n648), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1060), .A2(new_n870), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n828), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n860), .A2(new_n1075), .A3(new_n864), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n892), .B(new_n828), .C1(new_n1066), .C2(new_n871), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n1065), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1065), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1073), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n827), .B1(new_n1060), .B2(new_n870), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n883), .A2(new_n1081), .A3(new_n884), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1077), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1063), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1076), .A2(new_n1077), .A3(new_n1065), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1071), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1080), .A2(new_n676), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n964), .A3(new_n1085), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n860), .A2(new_n773), .A3(new_n864), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT54), .B(G143), .Z(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1092), .A2(new_n718), .B1(new_n936), .B2(new_n722), .ZN(new_n1093));
  INV_X1    g0893(.A(G125), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n738), .A2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(G128), .C2(new_n747), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n265), .B1(new_n748), .B2(new_n376), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n754), .A2(new_n298), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1097), .B(new_n1100), .C1(G132), .C2(new_n730), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1096), .B(new_n1101), .C1(new_n214), .C2(new_n734), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n747), .A2(G283), .B1(G107), .B2(new_n723), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n207), .B2(new_n718), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT122), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n275), .B1(new_n729), .B2(new_n221), .C1(new_n559), .C2(new_n754), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n739), .B2(G294), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1105), .B(new_n1107), .C1(new_n216), .C2(new_n734), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1102), .B1(new_n1108), .B2(new_n1038), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1109), .A2(new_n714), .B1(new_n399), .B2(new_n815), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1090), .A2(new_n713), .A3(new_n1110), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1088), .A2(new_n1089), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G378));
  INV_X1    g0913(.A(KEYINPUT57), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1087), .A2(new_n1072), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n313), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n301), .A2(new_n655), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n313), .B1(new_n301), .B2(new_n655), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT55), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT55), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1118), .A2(new_n1122), .A3(new_n1119), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT56), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1121), .A2(KEYINPUT56), .A3(new_n1123), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT40), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n896), .B2(new_n892), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n690), .A2(new_n894), .A3(new_n691), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n850), .A2(new_n861), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT40), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n1128), .C1(new_n1130), .C2(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n898), .B2(new_n710), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n880), .A2(new_n886), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1134), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n885), .A2(KEYINPUT108), .A3(new_n878), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT108), .B1(new_n885), .B2(new_n878), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1114), .B1(new_n1115), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1087), .A2(new_n1072), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(KEYINPUT57), .A3(new_n1137), .A4(new_n1141), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n676), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n964), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n815), .A2(new_n214), .ZN(new_n1149));
  INV_X1    g0949(.A(G124), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n273), .B(new_n260), .C1(new_n737), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n748), .A2(new_n298), .ZN(new_n1152));
  INV_X1    g0952(.A(G128), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1153), .A2(new_n729), .B1(new_n722), .B2(new_n812), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(new_n797), .C2(new_n1091), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n1094), .B2(new_n746), .C1(new_n936), .C2(new_n718), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1151), .B1(new_n1156), .B2(KEYINPUT59), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(KEYINPUT59), .B2(new_n1156), .C1(new_n376), .C2(new_n734), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G50), .B1(new_n273), .B2(new_n260), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n265), .B2(G41), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n746), .A2(new_n221), .B1(new_n738), .B2(new_n732), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n730), .A2(G107), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n723), .A2(G97), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n762), .A2(new_n381), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n927), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n260), .B(new_n275), .C1(new_n754), .C2(new_n269), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT123), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(new_n565), .C2(new_n718), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT58), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1158), .A2(new_n1160), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n709), .B1(new_n1171), .B2(new_n714), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1149), .B(new_n1172), .C1(new_n1128), .C2(new_n774), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT124), .Z(new_n1174));
  NOR2_X1   g0974(.A1(new_n1148), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1146), .A2(new_n1175), .ZN(G375));
  NOR2_X1   g0976(.A1(new_n870), .A2(new_n774), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n738), .A2(new_n753), .B1(new_n207), .B2(new_n754), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT125), .Z(new_n1179));
  NOR2_X1   g0979(.A1(new_n565), .A2(new_n748), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G116), .A2(new_n723), .B1(new_n804), .B2(G107), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n732), .B2(new_n729), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(G294), .C2(new_n747), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1179), .A2(new_n1183), .A3(new_n275), .A4(new_n935), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G159), .A2(new_n797), .B1(new_n723), .B2(new_n1091), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n1164), .C1(new_n298), .C2(new_n718), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n275), .B(new_n1186), .C1(G50), .C2(new_n749), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n747), .A2(G132), .B1(G137), .B2(new_n761), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n1153), .C2(new_n738), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n715), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n714), .A2(G68), .A3(new_n773), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1177), .A2(new_n709), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1069), .B2(new_n964), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1064), .A2(new_n1071), .A3(new_n1068), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n998), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1195), .B2(new_n1086), .ZN(G381));
  OR3_X1    g0996(.A1(G387), .A2(G384), .A3(G381), .ZN(new_n1197));
  INV_X1    g0997(.A(G396), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1007), .A2(new_n1198), .A3(new_n1008), .A4(new_n1032), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1146), .A2(new_n1112), .A3(new_n1175), .ZN(new_n1200));
  OR4_X1    g1000(.A1(G390), .A2(new_n1197), .A3(new_n1199), .A4(new_n1200), .ZN(G407));
  NAND2_X1  g1001(.A1(new_n656), .A2(G213), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT126), .Z(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(G407), .B(G213), .C1(new_n1200), .C2(new_n1204), .ZN(G409));
  NAND2_X1  g1005(.A1(new_n1142), .A2(KEYINPUT127), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT127), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1137), .A2(new_n1141), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1147), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1144), .A2(new_n998), .A3(new_n1137), .A4(new_n1141), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1173), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1203), .B1(new_n1212), .B2(new_n1112), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(G375), .A2(G378), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT60), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1194), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1064), .A2(new_n1068), .A3(KEYINPUT60), .A4(new_n1071), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1216), .A2(new_n1073), .A3(new_n676), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1193), .ZN(new_n1219));
  INV_X1    g1019(.A(G384), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(G384), .A3(new_n1193), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1213), .A2(new_n1214), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1203), .A2(G2897), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1223), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1221), .A2(new_n1222), .A3(new_n1226), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT63), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1225), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1199), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n961), .A2(new_n962), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n998), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n993), .A2(new_n978), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n975), .A2(new_n670), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT111), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1240), .A2(new_n989), .A3(new_n984), .A4(new_n976), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1237), .B1(new_n1241), .B2(new_n705), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1236), .B1(new_n1242), .B2(new_n964), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G390), .B1(new_n1243), .B2(new_n944), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n944), .B(G390), .C1(new_n963), .C2(new_n999), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1235), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G390), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G387), .A2(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1249), .A2(new_n1199), .A3(new_n1234), .A4(new_n1245), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1137), .A2(new_n1141), .A3(new_n1207), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1207), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n964), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1254), .A2(new_n1112), .A3(new_n1173), .A4(new_n1210), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1204), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1112), .B1(new_n1146), .B2(new_n1175), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1256), .A2(new_n1257), .A3(new_n1223), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1251), .B1(new_n1258), .B2(KEYINPUT63), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1233), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT62), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1224), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1260), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(new_n1256), .A2(new_n1257), .A3(KEYINPUT62), .A4(new_n1223), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1264), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1251), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1261), .B1(new_n1269), .B2(new_n1270), .ZN(G405));
  NAND2_X1  g1071(.A1(new_n1214), .A2(new_n1200), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1224), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1214), .A2(new_n1200), .A3(new_n1223), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(new_n1270), .ZN(G402));
endmodule


