//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n191), .A2(KEYINPUT73), .A3(G125), .ZN(new_n192));
  AOI21_X1  g006(.A(KEYINPUT73), .B1(new_n191), .B2(G125), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT74), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n191), .B2(G125), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT74), .A3(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n190), .B1(new_n194), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n190), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(G146), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n193), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n191), .A2(KEYINPUT73), .A3(G125), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n199), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(new_n202), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT71), .B1(new_n212), .B2(G128), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n213), .A2(KEYINPUT23), .B1(new_n212), .B2(G128), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G119), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(KEYINPUT71), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G110), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT72), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT72), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n222), .A3(G110), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n212), .A2(G128), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT24), .B(G110), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n211), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT75), .B1(new_n219), .B2(G110), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n227), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n232));
  INV_X1    g046(.A(G110), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n214), .A2(new_n232), .A3(new_n233), .A4(new_n218), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n197), .A2(G140), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n201), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G146), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n204), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G137), .ZN(new_n241));
  INV_X1    g055(.A(G953), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n242), .A2(G221), .A3(G234), .ZN(new_n243));
  XOR2_X1   g057(.A(new_n241), .B(new_n243), .Z(new_n244));
  AND3_X1   g058(.A1(new_n229), .A2(new_n240), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n229), .B2(new_n240), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT25), .B1(new_n247), .B2(new_n188), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT25), .ZN(new_n249));
  NOR4_X1   g063(.A1(new_n245), .A2(new_n246), .A3(new_n249), .A4(G902), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n189), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n247), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n189), .A2(G902), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(G472), .A2(G902), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n209), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G143), .B(G146), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT65), .A3(new_n260), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT0), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n215), .A3(KEYINPUT64), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n268), .B1(KEYINPUT0), .B2(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n260), .B1(new_n257), .B2(new_n259), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n263), .A2(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT11), .B1(new_n273), .B2(G137), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(G134), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G131), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n276), .B2(G134), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n273), .A2(KEYINPUT67), .A3(G137), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n278), .A2(new_n279), .A3(new_n281), .A4(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n281), .A2(new_n282), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n279), .B1(new_n285), .B2(new_n278), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n272), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT2), .B(G113), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n212), .A2(G116), .ZN(new_n290));
  INV_X1    g104(.A(G116), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G119), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n292), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n288), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT68), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n273), .B2(G137), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n273), .A2(G137), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n276), .A2(KEYINPUT68), .A3(G134), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G131), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n257), .B(new_n259), .C1(KEYINPUT1), .C2(new_n215), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n257), .A2(new_n259), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(G128), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n283), .A2(new_n304), .A3(new_n305), .A4(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n287), .A2(new_n298), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT28), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n287), .A2(new_n312), .A3(new_n298), .A4(new_n309), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n271), .A2(new_n270), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT65), .B1(new_n264), .B2(new_n260), .ZN(new_n316));
  AND4_X1   g130(.A1(KEYINPUT65), .A2(new_n257), .A3(new_n259), .A4(new_n260), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT66), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n263), .A2(new_n265), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT66), .A3(new_n315), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n274), .A2(new_n277), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n281), .A2(new_n282), .ZN(new_n324));
  OAI21_X1  g138(.A(G131), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n283), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n309), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n297), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n314), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(G237), .A2(G953), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G210), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT27), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G101), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n287), .A2(KEYINPUT30), .A3(new_n309), .ZN(new_n338));
  INV_X1    g152(.A(new_n309), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n318), .A2(new_n319), .B1(new_n325), .B2(new_n283), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n322), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n297), .B(new_n338), .C1(new_n341), .C2(KEYINPUT30), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT31), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT69), .B1(new_n310), .B2(new_n335), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n310), .A2(KEYINPUT69), .A3(new_n335), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n310), .A2(KEYINPUT69), .A3(new_n335), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n343), .B1(new_n350), .B2(new_n342), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n256), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT32), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT32), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n354), .B(new_n256), .C1(new_n347), .C2(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n314), .A2(new_n335), .A3(new_n329), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n335), .B1(new_n342), .B2(new_n310), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT70), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n342), .A2(new_n310), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n336), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n311), .A2(new_n313), .B1(new_n328), .B2(new_n297), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n364), .B2(new_n335), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT70), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n287), .A2(new_n309), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n297), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n314), .A2(KEYINPUT29), .A3(new_n335), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n188), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n361), .A2(new_n367), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G472), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n255), .B1(new_n356), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G107), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n379), .A2(KEYINPUT3), .A3(G104), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT3), .B1(new_n379), .B2(G104), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(G101), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n384), .A2(new_n321), .A3(new_n315), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT76), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n377), .B2(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n379), .A2(KEYINPUT3), .A3(G104), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n388), .A2(new_n389), .B1(new_n377), .B2(G107), .ZN(new_n390));
  INV_X1    g204(.A(G101), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n386), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n382), .A2(KEYINPUT76), .A3(G101), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n391), .B(new_n378), .C1(new_n380), .C2(new_n381), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT4), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n385), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n308), .A2(new_n305), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT77), .B1(new_n379), .B2(G104), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT77), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n377), .A3(G107), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n379), .A2(G104), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G101), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT78), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n405), .A2(new_n406), .A3(new_n394), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n406), .B1(new_n405), .B2(new_n394), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n399), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n326), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n405), .A2(new_n394), .A3(new_n308), .A4(new_n305), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n398), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n396), .A2(new_n409), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n396), .A2(new_n409), .A3(new_n412), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n414), .A2(new_n415), .A3(new_n326), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n414), .B2(new_n326), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G140), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n242), .A2(G227), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n421), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n397), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n407), .A2(new_n408), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n411), .ZN(new_n427));
  OAI221_X1 g241(.A(new_n326), .B1(KEYINPUT79), .B2(KEYINPUT12), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n326), .B1(new_n426), .B2(new_n427), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT12), .B1(new_n326), .B2(KEYINPUT79), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n424), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n422), .B2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT81), .B(G469), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n428), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n423), .B1(new_n437), .B2(new_n413), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n414), .A2(new_n326), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT80), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n414), .A2(new_n415), .A3(new_n326), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n424), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n188), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n434), .A2(new_n436), .B1(new_n443), .B2(G469), .ZN(new_n444));
  INV_X1    g258(.A(G221), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT9), .B(G234), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n447), .B2(new_n188), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n376), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n440), .A2(new_n441), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n423), .B1(new_n450), .B2(new_n413), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n188), .B(new_n436), .C1(new_n451), .C2(new_n432), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n443), .A2(G469), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT82), .ZN(new_n455));
  OAI21_X1  g269(.A(G210), .B1(G237), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G122), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n297), .A2(new_n384), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT76), .B1(new_n382), .B2(G101), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n460), .B1(new_n463), .B2(new_n393), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g280(.A(G113), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n294), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n405), .A2(new_n394), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT78), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n405), .A2(new_n406), .A3(new_n394), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n459), .B1(new_n464), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n395), .A2(new_n297), .A3(new_n384), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n294), .B(new_n469), .C1(new_n407), .C2(new_n408), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n458), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n480), .B(new_n459), .C1(new_n464), .C2(new_n474), .ZN(new_n481));
  AOI21_X1  g295(.A(G125), .B1(new_n308), .B2(new_n305), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n272), .B2(new_n197), .ZN(new_n484));
  INV_X1    g298(.A(G224), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(G953), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n484), .B(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n479), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n465), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n293), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n468), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n492), .B(new_n294), .C1(new_n407), .C2(new_n408), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n470), .A2(new_n471), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n458), .B(KEYINPUT8), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n197), .B1(new_n321), .B2(new_n315), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n499));
  OAI22_X1  g313(.A1(new_n498), .A2(new_n482), .B1(new_n499), .B2(new_n486), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n486), .A2(new_n499), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n483), .B(new_n501), .C1(new_n197), .C2(new_n272), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n478), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n188), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n457), .B1(new_n488), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n502), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n464), .A2(new_n474), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n507), .B2(new_n458), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n495), .A2(new_n496), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n479), .A2(new_n481), .A3(new_n487), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n456), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(KEYINPUT85), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G214), .B1(G237), .B2(G902), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(KEYINPUT83), .Z(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n510), .A2(new_n511), .A3(new_n456), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT85), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G478), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n446), .A2(new_n187), .A3(G953), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(KEYINPUT91), .A2(G122), .ZN(new_n525));
  NAND2_X1  g339(.A1(KEYINPUT91), .A2(G122), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n291), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G122), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT14), .B1(new_n528), .B2(G116), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n291), .A3(G122), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G107), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n258), .A2(G128), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n215), .A2(G143), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n534), .A2(new_n535), .A3(G134), .ZN(new_n536));
  AOI21_X1  g350(.A(G134), .B1(new_n534), .B2(new_n535), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n526), .ZN(new_n539));
  NOR2_X1   g353(.A1(KEYINPUT91), .A2(G122), .ZN(new_n540));
  OAI21_X1  g354(.A(G116), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n528), .A2(G116), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n379), .A3(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n533), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G107), .B1(new_n527), .B2(new_n542), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n258), .A2(G128), .ZN(new_n547));
  OAI21_X1  g361(.A(G134), .B1(new_n547), .B2(KEYINPUT13), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n534), .A2(new_n535), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT13), .A4(G134), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n546), .A2(new_n544), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n545), .A2(new_n552), .A3(KEYINPUT92), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n546), .A2(new_n544), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n551), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n533), .A2(new_n538), .A3(new_n544), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n524), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT92), .B1(new_n545), .B2(new_n552), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n554), .A3(new_n558), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n523), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT93), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n522), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n563), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n523), .B1(new_n561), .B2(new_n562), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n188), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT93), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n564), .A2(new_n565), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n566), .B1(new_n572), .B2(new_n522), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n331), .A2(G143), .A3(G214), .ZN(new_n574));
  AOI21_X1  g388(.A(G143), .B1(new_n331), .B2(G214), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT17), .B(G131), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT89), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n331), .A2(G214), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n258), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n331), .A2(G143), .A3(G214), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n582), .A2(KEYINPUT89), .A3(KEYINPUT17), .A4(G131), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(G131), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(new_n279), .A3(new_n581), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n584), .A2(new_n204), .A3(new_n210), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n582), .A2(KEYINPUT18), .A3(G131), .ZN(new_n590));
  NAND2_X1  g404(.A1(KEYINPUT18), .A2(G131), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n580), .A2(new_n581), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n209), .B1(new_n194), .B2(new_n199), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n590), .B(new_n592), .C1(new_n238), .C2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(G113), .B(G122), .Z(new_n595));
  XOR2_X1   g409(.A(KEYINPUT88), .B(G104), .Z(new_n596));
  XOR2_X1   g410(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND3_X1  g411(.A1(new_n589), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT90), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT90), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n589), .A2(new_n600), .A3(new_n594), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT19), .ZN(new_n603));
  AOI211_X1 g417(.A(KEYINPUT87), .B(new_n603), .C1(new_n194), .C2(new_n199), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n236), .A2(new_n201), .A3(new_n603), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT87), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n207), .B2(KEYINPUT19), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n209), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n585), .A2(new_n587), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n204), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n597), .B1(new_n610), .B2(new_n594), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT20), .ZN(new_n614));
  NOR2_X1   g428(.A1(G475), .A2(G902), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n611), .B1(new_n599), .B2(new_n601), .ZN(new_n619));
  INV_X1    g433(.A(new_n615), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n597), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n589), .A2(new_n594), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n599), .A2(new_n601), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(G475), .B1(new_n625), .B2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(G234), .A2(G237), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n627), .A2(G952), .A3(new_n242), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(G902), .A3(G953), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT94), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT21), .B(G898), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n573), .A2(new_n622), .A3(new_n626), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n520), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n375), .A2(new_n449), .A3(new_n455), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  NOR2_X1   g451(.A1(new_n564), .A2(G478), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n560), .A2(KEYINPUT33), .A3(new_n563), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT33), .B1(new_n560), .B2(new_n563), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n188), .A2(G478), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n622), .B2(new_n626), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n515), .B1(new_n505), .B2(new_n512), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n633), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n644), .A2(KEYINPUT96), .A3(new_n633), .A4(new_n645), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n454), .A2(KEYINPUT82), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n376), .B(new_n448), .C1(new_n452), .C2(new_n453), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n188), .B1(new_n347), .B2(new_n351), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT95), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(G472), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n252), .A2(new_n254), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n229), .A2(new_n240), .ZN(new_n659));
  INV_X1    g473(.A(new_n244), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n229), .A2(new_n240), .A3(new_n244), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n188), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n249), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n657), .B1(new_n665), .B2(new_n189), .ZN(new_n666));
  INV_X1    g480(.A(G472), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n345), .A2(new_n344), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT30), .B1(new_n327), .B2(new_n309), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n287), .A2(KEYINPUT30), .A3(new_n309), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n669), .A2(new_n298), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT31), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n346), .A3(new_n337), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n667), .B1(new_n673), .B2(new_n188), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT95), .B1(new_n673), .B2(new_n256), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n656), .B(new_n666), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n650), .A2(new_n653), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n377), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G6));
  NOR2_X1   g495(.A1(new_n564), .A2(new_n565), .ZN(new_n682));
  AOI211_X1 g496(.A(KEYINPUT93), .B(G902), .C1(new_n560), .C2(new_n563), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n522), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n566), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n632), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n613), .A2(new_n617), .A3(new_n615), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n624), .A2(new_n623), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n602), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n188), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n687), .A2(new_n621), .B1(new_n690), .B2(G475), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n645), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n653), .A2(new_n677), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G107), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  NOR2_X1   g510(.A1(new_n660), .A2(KEYINPUT36), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n659), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n253), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n251), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n700), .B(new_n656), .C1(new_n674), .C2(new_n675), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT99), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n654), .A2(G472), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n352), .A2(new_n655), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(KEYINPUT99), .A3(new_n656), .A4(new_n700), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n653), .A2(new_n635), .A3(new_n703), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT37), .B(G110), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G12));
  NAND2_X1  g524(.A1(new_n687), .A2(new_n621), .ZN(new_n711));
  INV_X1    g525(.A(new_n628), .ZN(new_n712));
  INV_X1    g526(.A(G900), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n630), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n712), .B1(new_n714), .B2(KEYINPUT100), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(KEYINPUT100), .B2(new_n714), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n711), .A2(new_n626), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(KEYINPUT101), .B1(new_n718), .B2(new_n573), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT101), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n684), .A2(new_n685), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n691), .A2(new_n720), .A3(new_n721), .A4(new_n717), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n353), .A2(new_n355), .B1(new_n373), .B2(G472), .ZN(new_n725));
  INV_X1    g539(.A(new_n645), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n665), .A2(new_n189), .B1(new_n253), .B2(new_n698), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n653), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G128), .ZN(G30));
  NAND2_X1  g544(.A1(new_n449), .A2(new_n455), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n716), .B(KEYINPUT39), .Z(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  OR3_X1    g547(.A1(new_n731), .A2(KEYINPUT40), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT40), .B1(new_n731), .B2(new_n733), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n512), .A2(KEYINPUT85), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n456), .B1(new_n510), .B2(new_n511), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n517), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n736), .B1(new_n738), .B2(KEYINPUT85), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT38), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n617), .B1(new_n613), .B2(new_n615), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n619), .A2(KEYINPUT20), .A3(new_n620), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n626), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n668), .A2(new_n671), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n335), .B1(new_n369), .B2(new_n310), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n188), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(G472), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n356), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n700), .A2(new_n515), .ZN(new_n749));
  AND4_X1   g563(.A1(new_n743), .A2(new_n748), .A3(new_n721), .A4(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n734), .A2(new_n735), .A3(new_n740), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G143), .ZN(G45));
  INV_X1    g566(.A(new_n643), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n743), .A2(new_n753), .A3(new_n717), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n653), .A2(new_n728), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G146), .ZN(G48));
  AOI21_X1  g571(.A(new_n432), .B1(new_n418), .B2(new_n421), .ZN(new_n758));
  OAI21_X1  g572(.A(G469), .B1(new_n758), .B2(G902), .ZN(new_n759));
  INV_X1    g573(.A(new_n448), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n452), .A3(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n725), .A2(new_n255), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n650), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT41), .B(G113), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G15));
  AOI21_X1  g579(.A(new_n354), .B1(new_n673), .B2(new_n256), .ZN(new_n766));
  INV_X1    g580(.A(new_n355), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n374), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n759), .A2(new_n452), .A3(new_n760), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n692), .A2(new_n768), .A3(new_n769), .A4(new_n666), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G116), .ZN(G18));
  OAI211_X1 g585(.A(new_n626), .B(new_n633), .C1(new_n741), .C2(new_n742), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n721), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n767), .A2(new_n766), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n363), .A2(new_n365), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n371), .B1(new_n775), .B2(KEYINPUT70), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n667), .B1(new_n776), .B2(new_n367), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n773), .B(new_n700), .C1(new_n774), .C2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n645), .A2(new_n759), .A3(new_n452), .A4(new_n760), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT102), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n727), .B1(new_n356), .B2(new_n374), .ZN(new_n781));
  INV_X1    g595(.A(new_n779), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT102), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .A4(new_n773), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G119), .ZN(G21));
  AND4_X1   g600(.A1(new_n760), .A2(new_n759), .A3(new_n452), .A4(new_n633), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n645), .A2(new_n743), .A3(new_n721), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n335), .B1(new_n314), .B2(new_n369), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT103), .B1(new_n351), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT103), .ZN(new_n791));
  INV_X1    g605(.A(new_n789), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n672), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n793), .A3(new_n346), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n674), .B1(new_n794), .B2(new_n256), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n787), .A2(new_n788), .A3(new_n666), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G122), .ZN(G24));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n256), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n798), .A2(new_n704), .A3(new_n700), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n754), .A2(KEYINPUT104), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT104), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n644), .A2(new_n801), .A3(new_n717), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n799), .A2(new_n782), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT105), .B(G125), .Z(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G27));
  INV_X1    g619(.A(KEYINPUT42), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT106), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n739), .B2(new_n515), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n513), .A2(new_n519), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(KEYINPUT106), .A3(new_n516), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n808), .A2(new_n375), .A3(new_n454), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n800), .A2(new_n802), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n806), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT106), .B1(new_n809), .B2(new_n516), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n807), .B(new_n515), .C1(new_n513), .C2(new_n519), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n452), .A2(new_n453), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n760), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n812), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(KEYINPUT42), .A3(new_n819), .A4(new_n375), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n813), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G131), .ZN(G33));
  INV_X1    g636(.A(KEYINPUT107), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n811), .B2(new_n723), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n818), .A2(KEYINPUT107), .A3(new_n375), .A4(new_n724), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G134), .ZN(G36));
  INV_X1    g641(.A(KEYINPUT109), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n438), .A2(new_n442), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT45), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(G469), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT108), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n829), .A2(new_n830), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(KEYINPUT108), .A3(G469), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(G469), .A2(G902), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT46), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n837), .A2(KEYINPUT46), .A3(new_n838), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n452), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n760), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n828), .B1(new_n844), .B2(new_n733), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(KEYINPUT109), .A3(new_n760), .A4(new_n732), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n727), .B1(new_n706), .B2(new_n656), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n753), .A2(new_n622), .A3(new_n626), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n848), .A2(KEYINPUT43), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(KEYINPUT43), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT44), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n814), .A2(new_n815), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n851), .B2(new_n853), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n845), .A2(new_n846), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(KEYINPUT111), .B(G137), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n859), .B(new_n860), .ZN(G39));
  XNOR2_X1  g675(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n844), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n843), .A2(new_n760), .A3(new_n862), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n808), .A2(new_n810), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n866), .A2(new_n768), .A3(new_n666), .A4(new_n754), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(G140), .ZN(G42));
  NOR2_X1   g683(.A1(new_n866), .A2(new_n761), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n748), .A2(new_n255), .A3(new_n712), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT119), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(KEYINPUT119), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n622), .A2(new_n626), .A3(new_n643), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n849), .A2(new_n628), .A3(new_n850), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n870), .A2(new_n799), .A3(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n798), .A2(new_n666), .A3(new_n704), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n740), .A2(new_n516), .A3(new_n761), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n881), .A2(KEYINPUT50), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT50), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n864), .A2(new_n865), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n759), .A2(new_n452), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n448), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n881), .A2(new_n855), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n873), .A2(new_n644), .A3(new_n874), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n870), .A2(new_n375), .A3(new_n878), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT48), .ZN(new_n898));
  INV_X1    g712(.A(G952), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n899), .B(G953), .C1(new_n881), .C2(new_n782), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n896), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT120), .Z(new_n902));
  OAI211_X1 g716(.A(new_n886), .B(KEYINPUT51), .C1(new_n891), .C2(new_n892), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n895), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT116), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n721), .A2(new_n622), .A3(new_n626), .A4(new_n633), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n520), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n677), .A2(new_n449), .A3(new_n455), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n703), .A2(new_n707), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n449), .A2(new_n455), .A3(new_n635), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT115), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n908), .B(KEYINPUT115), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n743), .A2(new_n633), .A3(new_n753), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(KEYINPUT114), .A3(new_n516), .A4(new_n739), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT114), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n644), .A2(new_n633), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n520), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n677), .A2(new_n449), .A3(new_n455), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n636), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n905), .B1(new_n915), .B2(new_n924), .ZN(new_n925));
  AOI211_X1 g739(.A(KEYINPUT116), .B(new_n923), .C1(new_n913), .C2(new_n914), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n718), .A2(new_n721), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n781), .A2(new_n449), .A3(new_n455), .A4(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n930), .B2(new_n866), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n781), .A2(new_n929), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n932), .A2(new_n653), .A3(new_n855), .A4(KEYINPUT117), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n808), .A2(new_n454), .A3(new_n810), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n826), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n759), .A2(new_n452), .A3(new_n760), .A4(new_n633), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n645), .A2(new_n743), .A3(new_n721), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI22_X1  g756(.A1(new_n762), .A2(new_n692), .B1(new_n880), .B2(new_n942), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n725), .A2(new_n634), .A3(new_n727), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n783), .B1(new_n944), .B2(new_n782), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n778), .A2(KEYINPUT102), .A3(new_n779), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n763), .B(new_n943), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n813), .B2(new_n820), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n781), .A2(new_n449), .A3(new_n455), .A4(new_n645), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n803), .B1(new_n949), .B2(new_n723), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT52), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n700), .A2(new_n716), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n748), .A2(new_n788), .A3(new_n454), .A4(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n951), .A2(new_n952), .A3(new_n756), .A4(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n729), .A2(new_n756), .A3(new_n803), .A4(new_n954), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT52), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n939), .A2(new_n948), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT53), .B1(new_n950), .B2(KEYINPUT52), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n927), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT115), .B1(new_n708), .B2(new_n908), .ZN(new_n961));
  INV_X1    g775(.A(new_n914), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n924), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT116), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n915), .A2(new_n905), .A3(new_n924), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n947), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n937), .B1(new_n931), .B2(new_n933), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n968), .A3(new_n821), .A4(new_n826), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n955), .A2(new_n957), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT53), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT54), .B1(new_n960), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT53), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n927), .B2(new_n958), .ZN(new_n975));
  AND4_X1   g789(.A1(KEYINPUT118), .A2(new_n785), .A3(new_n763), .A4(new_n943), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n768), .A2(new_n769), .A3(new_n666), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n648), .B2(new_n649), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n770), .A2(new_n796), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT118), .B1(new_n980), .B2(new_n785), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n974), .B1(new_n950), .B2(KEYINPUT52), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n968), .A2(new_n983), .A3(new_n821), .A4(new_n826), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n970), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n966), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT54), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n975), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n973), .A2(new_n989), .ZN(new_n990));
  OAI22_X1  g804(.A1(new_n904), .A2(new_n990), .B1(G952), .B2(G953), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT113), .ZN(new_n992));
  NOR4_X1   g806(.A1(new_n848), .A2(new_n255), .A3(new_n448), .A4(new_n515), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n740), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n888), .A2(KEYINPUT49), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n888), .A2(KEYINPUT49), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n995), .A2(new_n996), .A3(new_n748), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n994), .B(new_n997), .C1(new_n992), .C2(new_n993), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n991), .A2(new_n998), .ZN(G75));
  NAND2_X1  g813(.A1(new_n479), .A2(new_n481), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(new_n487), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT55), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n188), .B1(new_n975), .B2(new_n987), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(G210), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT56), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g820(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1007));
  NAND2_X1  g821(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1008), .B1(new_n1003), .B2(G210), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n242), .A2(G952), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT122), .Z(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1006), .A2(new_n1009), .A3(new_n1012), .ZN(G51));
  XOR2_X1   g827(.A(new_n838), .B(KEYINPUT57), .Z(new_n1014));
  AND3_X1   g828(.A1(new_n975), .A2(new_n988), .A3(new_n987), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n988), .B1(new_n975), .B2(new_n987), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n758), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1003), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1010), .B1(new_n1019), .B2(new_n1020), .ZN(G54));
  AND2_X1   g835(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1003), .A2(new_n613), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n613), .B1(new_n1003), .B2(new_n1022), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1023), .A2(new_n1024), .A3(new_n1010), .ZN(G60));
  XOR2_X1   g839(.A(new_n641), .B(KEYINPUT123), .Z(new_n1026));
  NAND2_X1  g840(.A1(G478), .A2(G902), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT59), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1026), .B(new_n1028), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(new_n1011), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1026), .B1(new_n990), .B2(new_n1028), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1030), .A2(new_n1031), .ZN(G63));
  INV_X1    g846(.A(KEYINPUT61), .ZN(new_n1033));
  NAND2_X1  g847(.A1(G217), .A2(G902), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT124), .Z(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT60), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1036), .B1(new_n975), .B2(new_n987), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n698), .B(KEYINPUT125), .Z(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1011), .B1(new_n1037), .B2(new_n247), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1033), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AND2_X1   g856(.A1(new_n975), .A2(new_n987), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n252), .B1(new_n1043), .B2(new_n1036), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1044), .A2(KEYINPUT61), .A3(new_n1011), .A4(new_n1039), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1042), .A2(new_n1045), .ZN(G66));
  NAND2_X1  g860(.A1(new_n966), .A2(new_n967), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1047), .A2(new_n242), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n631), .A2(new_n485), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(G953), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1048), .A2(KEYINPUT126), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1052), .B1(KEYINPUT126), .B2(new_n1048), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1000), .B1(G898), .B2(new_n242), .ZN(new_n1054));
  INV_X1    g868(.A(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g869(.A(new_n1053), .B(new_n1055), .ZN(G69));
  NOR2_X1   g870(.A1(new_n669), .A2(new_n670), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n604), .A2(new_n607), .ZN(new_n1058));
  XNOR2_X1  g872(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1059), .B1(G900), .B2(G953), .ZN(new_n1060));
  NOR3_X1   g874(.A1(new_n725), .A2(new_n941), .A3(new_n255), .ZN(new_n1061));
  OAI211_X1 g875(.A(new_n845), .B(new_n846), .C1(new_n858), .C2(new_n1061), .ZN(new_n1062));
  AND3_X1   g876(.A1(new_n729), .A2(new_n756), .A3(new_n803), .ZN(new_n1063));
  AND3_X1   g877(.A1(new_n1063), .A2(new_n821), .A3(new_n826), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1062), .A2(new_n868), .A3(new_n1064), .ZN(new_n1065));
  OAI21_X1  g879(.A(new_n1060), .B1(new_n1065), .B2(G953), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n751), .A2(new_n1063), .ZN(new_n1067));
  INV_X1    g881(.A(KEYINPUT62), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n751), .A2(new_n1063), .A3(KEYINPUT62), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g885(.A1(new_n731), .A2(new_n733), .ZN(new_n1072));
  INV_X1    g886(.A(new_n644), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n1073), .B1(new_n743), .B2(new_n573), .ZN(new_n1074));
  NAND4_X1  g888(.A1(new_n1072), .A2(new_n375), .A3(new_n855), .A4(new_n1074), .ZN(new_n1075));
  NAND4_X1  g889(.A1(new_n859), .A2(new_n1071), .A3(new_n868), .A4(new_n1075), .ZN(new_n1076));
  AND2_X1   g890(.A1(new_n1076), .A2(new_n242), .ZN(new_n1077));
  INV_X1    g891(.A(new_n1059), .ZN(new_n1078));
  OAI21_X1  g892(.A(new_n1066), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g893(.A1(new_n1059), .A2(KEYINPUT127), .ZN(new_n1080));
  AOI211_X1 g894(.A(new_n242), .B(new_n1080), .C1(G227), .C2(G900), .ZN(new_n1081));
  XNOR2_X1  g895(.A(new_n1079), .B(new_n1081), .ZN(G72));
  NAND2_X1  g896(.A1(G472), .A2(G902), .ZN(new_n1083));
  XOR2_X1   g897(.A(new_n1083), .B(KEYINPUT63), .Z(new_n1084));
  OAI21_X1  g898(.A(new_n1084), .B1(new_n1065), .B2(new_n1047), .ZN(new_n1085));
  NAND2_X1  g899(.A1(new_n1085), .A2(new_n336), .ZN(new_n1086));
  OAI21_X1  g900(.A(new_n1084), .B1(new_n1076), .B2(new_n1047), .ZN(new_n1087));
  NAND2_X1  g901(.A1(new_n1087), .A2(new_n362), .ZN(new_n1088));
  AOI21_X1  g902(.A(new_n360), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OAI221_X1 g903(.A(new_n1084), .B1(new_n744), .B2(new_n360), .C1(new_n960), .C2(new_n972), .ZN(new_n1090));
  OAI21_X1  g904(.A(new_n1090), .B1(G952), .B2(new_n242), .ZN(new_n1091));
  NOR2_X1   g905(.A1(new_n1089), .A2(new_n1091), .ZN(G57));
endmodule


