//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT35), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G78gat), .B(G106gat), .ZN(new_n206));
  INV_X1    g005(.A(G50gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G228gat), .ZN(new_n210));
  INV_X1    g009(.A(G233gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n218), .B1(G155gat), .B2(G162gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G141gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G155gat), .B(G162gat), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT2), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n220), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(KEYINPUT29), .ZN(new_n233));
  OR2_X1    g032(.A1(G211gat), .A2(G218gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(G211gat), .A2(G218gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(KEYINPUT77), .A3(new_n235), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(KEYINPUT76), .A3(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(G197gat), .A2(G204gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(G197gat), .A2(G204gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n241), .A2(new_n242), .B1(new_n243), .B2(new_n235), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n244), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n246), .A2(KEYINPUT76), .A3(new_n238), .A4(new_n239), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n213), .B1(new_n233), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n239), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n246), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT29), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n238), .A2(new_n239), .A3(new_n244), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT87), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT87), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n251), .A2(new_n256), .A3(new_n252), .A4(new_n253), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n231), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n220), .A2(new_n230), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT80), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n220), .A2(new_n230), .A3(KEYINPUT80), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n249), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT29), .B1(new_n245), .B2(new_n247), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n259), .B1(new_n266), .B2(KEYINPUT3), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n245), .A2(new_n247), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(KEYINPUT29), .B2(new_n232), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n213), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G22gat), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT86), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(G22gat), .B1(new_n265), .B2(new_n270), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n209), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT86), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n258), .A2(new_n264), .ZN(new_n277));
  INV_X1    g076(.A(new_n249), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n267), .A2(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n212), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n281), .A3(new_n272), .ZN(new_n282));
  AND4_X1   g081(.A1(new_n276), .A2(new_n282), .A3(new_n209), .A4(new_n274), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n205), .B1(new_n275), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n274), .A3(new_n276), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n208), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n273), .A2(new_n209), .A3(new_n274), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n204), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n290));
  INV_X1    g089(.A(G183gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT27), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT27), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G183gat), .ZN(new_n294));
  INV_X1    g093(.A(G190gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT28), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT27), .B1(new_n298), .B2(new_n291), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n293), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n307), .A2(KEYINPUT26), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(KEYINPUT26), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(new_n291), .B2(new_n295), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n303), .B1(new_n297), .B2(new_n302), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT23), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  OAI211_X1 g116(.A(KEYINPUT25), .B(new_n315), .C1(new_n317), .C2(new_n308), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n291), .A2(new_n295), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT65), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n318), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n316), .A2(G169gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT23), .B1(new_n305), .B2(new_n306), .ZN(new_n330));
  INV_X1    g129(.A(new_n308), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n328), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n322), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(new_n319), .A3(new_n320), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT25), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI22_X1  g134(.A1(new_n313), .A2(new_n314), .B1(new_n325), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G120gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G113gat), .ZN(new_n338));
  INV_X1    g137(.A(G113gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G120gat), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT1), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G127gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G134gat), .ZN(new_n346));
  INV_X1    g145(.A(G134gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G127gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n348), .A3(KEYINPUT68), .ZN(new_n349));
  OR3_X1    g148(.A1(new_n347), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT69), .B1(new_n351), .B2(new_n341), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n338), .A2(new_n340), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n349), .A4(new_n350), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n344), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n324), .A2(new_n321), .ZN(new_n360));
  INV_X1    g159(.A(new_n318), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n332), .A2(new_n334), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(KEYINPUT25), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n351), .A2(KEYINPUT69), .A3(new_n341), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n347), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(new_n342), .B2(KEYINPUT68), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n356), .B1(new_n367), .B2(new_n355), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n343), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n297), .A2(new_n302), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT67), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n304), .A3(new_n312), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n364), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n359), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n290), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n375), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT72), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT34), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI211_X1 g179(.A(new_n377), .B(new_n380), .C1(new_n359), .C2(new_n373), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n359), .A2(new_n377), .A3(new_n373), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT32), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT71), .B(G71gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G99gat), .ZN(new_n388));
  XOR2_X1   g187(.A(G15gat), .B(G43gat), .Z(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n384), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n383), .B(KEYINPUT32), .C1(new_n385), .C2(new_n390), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n382), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT74), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n382), .A2(new_n392), .A3(new_n396), .A4(new_n393), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT73), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n374), .A2(new_n375), .ZN(new_n400));
  INV_X1    g199(.A(new_n290), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n374), .B(new_n375), .C1(new_n378), .C2(new_n379), .ZN(new_n403));
  AOI221_X4 g202(.A(new_n399), .B1(new_n402), .B2(new_n403), .C1(new_n392), .C2(new_n393), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n392), .A2(new_n393), .ZN(new_n405));
  INV_X1    g204(.A(new_n382), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT73), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n395), .A2(new_n398), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n289), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n410), .B(KEYINPUT78), .Z(new_n411));
  AOI21_X1  g210(.A(new_n411), .B1(new_n336), .B2(new_n252), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n364), .B2(new_n372), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n268), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n336), .A2(new_n411), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n364), .B2(new_n372), .ZN(new_n416));
  INV_X1    g215(.A(new_n410), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n415), .B(new_n248), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  NAND3_X1  g220(.A1(new_n414), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n414), .B2(new_n418), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(KEYINPUT79), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT79), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n414), .A2(new_n418), .A3(new_n428), .A4(new_n421), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n423), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n259), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(new_n343), .C1(new_n365), .C2(new_n368), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT4), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT83), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n263), .A2(new_n358), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(new_n438), .A3(KEYINPUT4), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n231), .B1(new_n220), .B2(new_n230), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n232), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n369), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n436), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n263), .A2(new_n358), .A3(KEYINPUT4), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n453), .A2(KEYINPUT5), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT81), .B1(new_n358), .B2(new_n432), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n369), .A2(new_n259), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n369), .A2(KEYINPUT81), .A3(new_n259), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n442), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT82), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  AND4_X1   g259(.A1(KEYINPUT82), .A2(new_n459), .A3(KEYINPUT5), .A4(new_n453), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n450), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G1gat), .B(G29gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT0), .ZN(new_n464));
  XNOR2_X1  g263(.A(G57gat), .B(G85gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n464), .B(new_n465), .Z(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT84), .B(KEYINPUT6), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n457), .A2(new_n442), .A3(new_n458), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n453), .A2(KEYINPUT5), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n459), .A2(KEYINPUT82), .A3(KEYINPUT5), .A4(new_n453), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n449), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n468), .A2(new_n469), .A3(new_n476), .ZN(new_n477));
  OR3_X1    g276(.A1(new_n475), .A2(new_n466), .A3(new_n469), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n431), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n203), .B1(new_n409), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n284), .A2(new_n288), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n482), .A2(new_n397), .B1(new_n405), .B2(new_n406), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n203), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n469), .B1(new_n475), .B2(new_n466), .ZN(new_n486));
  AOI211_X1 g285(.A(new_n467), .B(new_n449), .C1(new_n473), .C2(new_n474), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n468), .A2(KEYINPUT89), .A3(new_n476), .A4(new_n469), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n478), .ZN(new_n490));
  INV_X1    g289(.A(new_n431), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n484), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(KEYINPUT91), .A3(new_n491), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n480), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT38), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n421), .A2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n425), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n414), .A2(new_n418), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT37), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n497), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n425), .A2(new_n499), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n248), .B1(new_n412), .B2(new_n413), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n415), .B(new_n268), .C1(new_n416), .C2(new_n417), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT37), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n497), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n427), .B(new_n429), .C1(new_n504), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n488), .A2(new_n489), .A3(new_n478), .A4(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n457), .A2(new_n458), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n512), .B(KEYINPUT39), .C1(new_n513), .C2(new_n442), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n369), .A2(new_n444), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n439), .A2(new_n437), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n438), .B1(new_n433), .B2(KEYINPUT4), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n442), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n442), .B1(new_n457), .B2(new_n458), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT39), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT88), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n441), .B1(new_n440), .B2(new_n515), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n467), .B1(new_n524), .B2(new_n521), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n523), .A2(KEYINPUT40), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT40), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n430), .A2(new_n426), .B1(new_n462), .B2(new_n467), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n528), .A2(new_n529), .B1(new_n288), .B2(new_n284), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n511), .A2(new_n530), .A3(KEYINPUT90), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT90), .B1(new_n511), .B2(new_n530), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI22_X1  g334(.A1(new_n408), .A2(new_n533), .B1(new_n483), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n479), .B2(new_n481), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n531), .A2(new_n532), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n496), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(G29gat), .A2(G36gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT14), .Z(new_n541));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n544));
  INV_X1    g343(.A(G29gat), .ZN(new_n545));
  INV_X1    g344(.A(G36gat), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT92), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n541), .A2(new_n543), .A3(new_n544), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n540), .B(KEYINPUT14), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT15), .B(new_n542), .C1(new_n550), .C2(new_n547), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G15gat), .B(G22gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT16), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(G1gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(G1gat), .B2(new_n555), .ZN(new_n558));
  INV_X1    g357(.A(G8gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n549), .A2(KEYINPUT17), .A3(new_n551), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n558), .B(G8gat), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n552), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n554), .A2(new_n560), .A3(new_n563), .A4(new_n561), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n566), .A2(new_n567), .B1(G229gat), .B2(G233gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT94), .B1(new_n568), .B2(KEYINPUT18), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G197gat), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT11), .B(G169gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT12), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n568), .A2(KEYINPUT18), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n560), .B(new_n552), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT13), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n579), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT18), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n576), .A2(new_n577), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n577), .ZN(new_n588));
  OAI22_X1  g387(.A1(new_n568), .A2(KEYINPUT18), .B1(new_n578), .B2(new_n581), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n569), .B(new_n575), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n202), .B1(new_n539), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(KEYINPUT95), .B(new_n591), .C1(new_n496), .C2(new_n538), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(G64gat), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT9), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(G64gat), .B1(new_n600), .B2(new_n601), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n596), .B(new_n599), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n597), .B1(new_n596), .B2(new_n603), .ZN(new_n608));
  INV_X1    g407(.A(G57gat), .ZN(new_n609));
  INV_X1    g408(.A(G64gat), .ZN(new_n610));
  OR3_X1    g409(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT98), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n609), .B2(KEYINPUT98), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n608), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G127gat), .B(G155gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  OAI21_X1  g417(.A(new_n560), .B1(new_n615), .B2(new_n614), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT99), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n620), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  INV_X1    g428(.A(G85gat), .ZN(new_n630));
  INV_X1    g429(.A(G92gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(KEYINPUT8), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT7), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n630), .B2(new_n631), .ZN(new_n634));
  NAND3_X1  g433(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G99gat), .B(G106gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n554), .A2(new_n561), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n552), .A2(new_n638), .B1(KEYINPUT41), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G190gat), .B(G218gat), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n644), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n640), .A2(new_n649), .A3(new_n642), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n648), .B1(new_n645), .B2(new_n650), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n628), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n638), .A2(KEYINPUT10), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n657), .B2(new_n614), .ZN(new_n658));
  INV_X1    g457(.A(new_n614), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n659), .A2(KEYINPUT102), .A3(KEYINPUT10), .A4(new_n638), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n614), .A2(new_n638), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n636), .A2(KEYINPUT100), .ZN(new_n664));
  INV_X1    g463(.A(new_n637), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n636), .A2(KEYINPUT100), .A3(new_n637), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n666), .A2(new_n607), .A3(new_n613), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT10), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n662), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI211_X1 g470(.A(KEYINPUT101), .B(KEYINPUT10), .C1(new_n663), .C2(new_n668), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n661), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT103), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n663), .A2(new_n668), .A3(new_n675), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(KEYINPUT104), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n677), .B2(new_n678), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(KEYINPUT105), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n687), .B(new_n681), .C1(new_n677), .C2(new_n678), .ZN(new_n688));
  OAI22_X1  g487(.A1(new_n683), .A2(new_n684), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n655), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT106), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(KEYINPUT106), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n595), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n477), .A2(new_n478), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT107), .B(G1gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1324gat));
  NOR2_X1   g497(.A1(new_n556), .A2(new_n559), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n700));
  NOR4_X1   g499(.A1(new_n694), .A2(new_n491), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(KEYINPUT42), .ZN(new_n702));
  INV_X1    g501(.A(new_n694), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n559), .B1(new_n703), .B2(new_n431), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT42), .B1(new_n704), .B2(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(G1325gat));
  INV_X1    g505(.A(new_n483), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n694), .A2(G15gat), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G15gat), .B1(new_n694), .B2(new_n536), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1326gat));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n481), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  INV_X1    g512(.A(new_n689), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n628), .A3(new_n653), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n715), .B1(new_n593), .B2(new_n594), .ZN(new_n716));
  INV_X1    g515(.A(new_n695), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(new_n545), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n653), .B1(new_n496), .B2(new_n538), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n511), .A2(new_n530), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT90), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n479), .ZN(new_n727));
  OAI221_X1 g526(.A(KEYINPUT36), .B1(new_n404), .B2(new_n407), .C1(new_n395), .C2(new_n398), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n707), .A2(new_n534), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n727), .A2(new_n289), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n511), .A2(new_n530), .A3(KEYINPUT90), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n726), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n490), .A2(KEYINPUT91), .A3(new_n491), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT91), .B1(new_n490), .B2(new_n491), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n733), .A2(new_n734), .A3(new_n484), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n735), .B2(new_n480), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(KEYINPUT44), .A3(new_n653), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n723), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n592), .A2(new_n689), .A3(new_n627), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G29gat), .B1(new_n740), .B2(new_n695), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n718), .A2(new_n719), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n720), .A2(new_n741), .A3(new_n742), .ZN(G1328gat));
  AND3_X1   g542(.A1(new_n716), .A2(new_n546), .A3(new_n431), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n745));
  OR2_X1    g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  OAI21_X1  g546(.A(G36gat), .B1(new_n740), .B2(new_n491), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(G1329gat));
  INV_X1    g548(.A(new_n536), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n723), .A2(new_n750), .A3(new_n737), .A4(new_n739), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G43gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n715), .A2(G43gat), .A3(new_n707), .ZN(new_n753));
  INV_X1    g552(.A(new_n594), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT95), .B1(new_n736), .B2(new_n591), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n752), .A2(KEYINPUT47), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT111), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n752), .A2(new_n759), .A3(KEYINPUT47), .A4(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n756), .A2(KEYINPUT109), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n763), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n752), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n761), .B1(new_n768), .B2(new_n769), .ZN(G1330gat));
  NAND4_X1  g569(.A1(new_n723), .A2(new_n289), .A3(new_n737), .A4(new_n739), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G50gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n481), .A2(G50gat), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n716), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT112), .B1(new_n771), .B2(G50gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n716), .B2(new_n775), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n780), .A2(KEYINPUT113), .A3(new_n772), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT113), .B1(new_n780), .B2(new_n772), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n778), .A2(KEYINPUT48), .B1(new_n781), .B2(new_n782), .ZN(G1331gat));
  NOR4_X1   g582(.A1(new_n539), .A2(new_n591), .A3(new_n655), .A4(new_n714), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n717), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G57gat), .ZN(G1332gat));
  INV_X1    g585(.A(KEYINPUT49), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n784), .B(new_n431), .C1(new_n787), .C2(new_n610), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n610), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1333gat));
  NAND2_X1  g589(.A1(new_n784), .A2(new_n483), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT115), .ZN(new_n792));
  INV_X1    g591(.A(G71gat), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n784), .A2(new_n794), .A3(new_n483), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n784), .A2(G71gat), .A3(new_n750), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT114), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n799), .A3(G71gat), .A4(new_n750), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT50), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n796), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1334gat));
  NAND2_X1  g605(.A1(new_n784), .A2(new_n289), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g607(.A1(new_n714), .A2(new_n591), .A3(new_n627), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n738), .A2(new_n717), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G85gat), .ZN(new_n811));
  INV_X1    g610(.A(new_n721), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n591), .A2(new_n627), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n812), .A2(KEYINPUT51), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT51), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n717), .A2(new_n630), .A3(new_n689), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n811), .B1(new_n816), .B2(new_n817), .ZN(G1336gat));
  NAND4_X1  g617(.A1(new_n723), .A2(new_n431), .A3(new_n737), .A4(new_n809), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(G92gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n689), .A2(new_n631), .A3(new_n431), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT116), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n823), .B(new_n826), .ZN(G1337gat));
  NAND3_X1  g626(.A1(new_n738), .A2(new_n750), .A3(new_n809), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT118), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G99gat), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n828), .A2(KEYINPUT118), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n714), .A2(G99gat), .A3(new_n707), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n830), .A2(new_n831), .B1(new_n816), .B2(new_n832), .ZN(G1338gat));
  NAND4_X1  g632(.A1(new_n723), .A2(new_n289), .A3(new_n737), .A4(new_n809), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G106gat), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n714), .A2(G106gat), .A3(new_n481), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n816), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g637(.A1(new_n690), .A2(new_n592), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n677), .A2(KEYINPUT54), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n681), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT10), .B1(new_n663), .B2(new_n668), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(new_n662), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n676), .B1(new_n658), .B2(new_n660), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n846), .A2(new_n847), .A3(new_n677), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n846), .B2(new_n677), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n841), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n586), .A2(new_n574), .A3(new_n577), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n578), .A2(new_n581), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n583), .B2(new_n579), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n573), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n853), .A2(new_n653), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n841), .B(KEYINPUT55), .C1(new_n848), .C2(new_n849), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n682), .B(KEYINPUT104), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n689), .A2(new_n856), .A3(new_n853), .ZN(new_n863));
  INV_X1    g662(.A(new_n852), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n591), .A3(new_n860), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n653), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n839), .B1(new_n868), .B2(new_n627), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(new_n717), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n491), .A3(new_n409), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(G113gat), .B1(new_n872), .B2(new_n591), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n869), .A2(new_n481), .A3(new_n483), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n717), .A3(new_n491), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n339), .A3(new_n592), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n873), .A2(new_n876), .ZN(G1340gat));
  AOI21_X1  g676(.A(G120gat), .B1(new_n872), .B2(new_n689), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n875), .A2(new_n337), .A3(new_n714), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(G1341gat));
  NAND3_X1  g679(.A1(new_n872), .A2(new_n345), .A3(new_n627), .ZN(new_n881));
  OAI21_X1  g680(.A(G127gat), .B1(new_n875), .B2(new_n628), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1342gat));
  NAND3_X1  g682(.A1(new_n872), .A2(new_n347), .A3(new_n653), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(KEYINPUT56), .ZN(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n875), .B2(new_n867), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(KEYINPUT56), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(G1343gat));
  NAND3_X1  g687(.A1(new_n536), .A2(new_n717), .A3(new_n491), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT120), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n869), .A2(new_n289), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT55), .B1(new_n850), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n841), .B(KEYINPUT121), .C1(new_n848), .C2(new_n849), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n859), .A2(new_n591), .A3(new_n860), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n850), .A2(new_n894), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n901), .A2(KEYINPUT122), .A3(new_n851), .A4(new_n896), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n653), .B1(new_n903), .B2(new_n863), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n628), .B1(new_n904), .B2(new_n862), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n481), .B1(new_n905), .B2(new_n839), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n893), .B1(new_n906), .B2(new_n892), .ZN(new_n907));
  OAI21_X1  g706(.A(G141gat), .B1(new_n907), .B2(new_n592), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n750), .A2(new_n431), .A3(new_n481), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n870), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n221), .A3(new_n591), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT58), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n908), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1344gat));
  NAND3_X1  g716(.A1(new_n911), .A2(new_n223), .A3(new_n689), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n907), .A2(new_n714), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n223), .A2(KEYINPUT59), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n481), .A2(KEYINPUT57), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n900), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT122), .B1(new_n895), .B2(new_n896), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n863), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n867), .ZN(new_n927));
  INV_X1    g726(.A(new_n862), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n627), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n691), .A2(new_n592), .A3(new_n692), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n923), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n869), .A2(new_n289), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT57), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n890), .A2(new_n714), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n922), .B1(new_n936), .B2(G148gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n918), .B1(new_n921), .B2(new_n937), .ZN(G1345gat));
  OAI21_X1  g737(.A(G155gat), .B1(new_n907), .B2(new_n628), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n911), .A2(new_n227), .A3(new_n627), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1346gat));
  OR3_X1    g740(.A1(new_n907), .A2(new_n228), .A3(new_n867), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n228), .B1(new_n910), .B2(new_n867), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(G1347gat));
  NOR2_X1   g743(.A1(new_n717), .A2(new_n491), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT124), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n874), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n948), .A2(new_n305), .A3(new_n592), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n869), .A2(new_n945), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n409), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT123), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n952), .A2(new_n592), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n949), .B1(new_n953), .B2(new_n305), .ZN(G1348gat));
  NOR3_X1   g753(.A1(new_n948), .A2(new_n328), .A3(new_n714), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n952), .A2(new_n714), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n306), .ZN(G1349gat));
  OAI21_X1  g756(.A(G183gat), .B1(new_n948), .B2(new_n628), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n627), .A2(new_n292), .A3(new_n294), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n951), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n948), .B2(new_n867), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT61), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n653), .A2(new_n295), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n952), .B2(new_n964), .ZN(G1351gat));
  NOR2_X1   g764(.A1(new_n750), .A2(new_n481), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(G197gat), .B1(new_n968), .B2(new_n591), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n946), .A2(new_n750), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n934), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n591), .A2(G197gat), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1352gat));
  NOR3_X1   g772(.A1(new_n967), .A2(G204gat), .A3(new_n714), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT62), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n934), .A2(new_n689), .A3(new_n970), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n977));
  OAI21_X1  g776(.A(G204gat), .B1(new_n976), .B2(KEYINPUT125), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1353gat));
  OR3_X1    g778(.A1(new_n967), .A2(G211gat), .A3(new_n628), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n931), .A2(new_n627), .A3(new_n933), .A4(new_n970), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g785(.A(KEYINPUT126), .B(new_n980), .C1(new_n982), .C2(new_n983), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1354gat));
  AOI21_X1  g787(.A(G218gat), .B1(new_n968), .B2(new_n653), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n653), .A2(G218gat), .ZN(new_n990));
  XOR2_X1   g789(.A(new_n990), .B(KEYINPUT127), .Z(new_n991));
  AOI21_X1  g790(.A(new_n989), .B1(new_n971), .B2(new_n991), .ZN(G1355gat));
endmodule


