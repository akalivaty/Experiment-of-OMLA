//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g0008(.A(G250), .B1(G257), .B2(G264), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n202), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n210), .A2(KEYINPUT0), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(KEYINPUT0), .B2(new_n210), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n219), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  INV_X1    g0042(.A(G50), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n245), .B(KEYINPUT67), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G50), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n211), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G1), .B2(new_n212), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n254), .B1(new_n258), .B2(G50), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT8), .A2(G58), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT70), .A2(G58), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT70), .A2(G58), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n262), .B1(new_n266), .B2(KEYINPUT8), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n212), .A2(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n261), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n259), .B1(new_n270), .B2(new_n256), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(new_n251), .A3(G274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(G1), .A2(G13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n251), .A2(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n276), .B1(new_n279), .B2(G226), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT68), .B(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G222), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G77), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n287), .B1(new_n288), .B2(new_n285), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n291), .A2(KEYINPUT69), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n291), .B2(KEYINPUT69), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n280), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(G169), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n271), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n271), .B(KEYINPUT9), .Z(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n296), .A2(G200), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n300), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT13), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n293), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G238), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n275), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT72), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n285), .A2(G226), .A3(new_n286), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G97), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n316), .C1(new_n289), .C2(new_n235), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n294), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n309), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(KEYINPUT73), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n314), .A2(new_n318), .A3(new_n309), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n320), .A2(G179), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n319), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n322), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(G169), .ZN(new_n327));
  INV_X1    g0127(.A(new_n322), .ZN(new_n328));
  OAI21_X1  g0128(.A(G169), .B1(new_n328), .B2(new_n319), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT14), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n323), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT12), .ZN(new_n332));
  INV_X1    g0132(.A(G13), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G1), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G68), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G20), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n332), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n334), .A2(KEYINPUT12), .A3(G20), .A4(new_n336), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n338), .B(new_n339), .C1(new_n258), .C2(new_n336), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT75), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n260), .A2(KEYINPUT74), .A3(G50), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n337), .C1(new_n288), .C2(new_n269), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT74), .B1(new_n260), .B2(G50), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n256), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT11), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n331), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n325), .B2(G200), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n320), .A2(G190), .A3(new_n321), .A4(new_n322), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n257), .B(G77), .C1(G1), .C2(new_n212), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(G77), .B2(new_n252), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G20), .A2(G77), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT8), .B(G58), .Z(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n260), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n354), .B1(new_n269), .B2(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n353), .B1(new_n359), .B2(new_n256), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n282), .A2(new_n284), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G107), .ZN(new_n363));
  INV_X1    g0163(.A(G1698), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT68), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT68), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G1698), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n282), .A2(new_n284), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n363), .B1(new_n235), .B2(new_n368), .C1(new_n289), .C2(new_n312), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n294), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n276), .B1(new_n279), .B2(G244), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n302), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n361), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G169), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n360), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n373), .A2(new_n297), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n379), .A2(new_n380), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n377), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n308), .A2(new_n348), .A3(new_n351), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT81), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n311), .B2(new_n235), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n293), .A2(new_n310), .A3(KEYINPUT81), .A4(G232), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n275), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n282), .A2(new_n284), .A3(G226), .A4(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(new_n392), .C1(new_n368), .C2(new_n290), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n390), .A2(KEYINPUT82), .B1(new_n294), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT83), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT82), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n388), .A2(new_n396), .A3(new_n389), .A4(new_n275), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n394), .A2(new_n395), .A3(new_n297), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT81), .B1(new_n279), .B2(G232), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n389), .A2(new_n275), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT82), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n393), .A2(new_n294), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT83), .B1(new_n403), .B2(new_n378), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n401), .A2(new_n397), .A3(new_n402), .A4(new_n297), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n398), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(G20), .B1(new_n282), .B2(new_n284), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT77), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT7), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT76), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT76), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT7), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n408), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n409), .B1(new_n408), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT78), .B1(new_n418), .B2(new_n336), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n202), .B1(new_n266), .B2(G68), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(new_n212), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n260), .A2(G159), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT79), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n283), .A2(G33), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n212), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n411), .A2(new_n413), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT77), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n408), .A2(new_n409), .A3(new_n414), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n410), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(G68), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n419), .A2(KEYINPUT16), .A3(new_n424), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT16), .ZN(new_n436));
  INV_X1    g0236(.A(new_n423), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n212), .B2(new_n420), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT80), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n282), .B1(new_n426), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n284), .A2(KEYINPUT80), .ZN(new_n441));
  OAI211_X1 g0241(.A(KEYINPUT7), .B(new_n212), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n427), .A2(new_n428), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n336), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n436), .B1(new_n438), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n435), .A2(new_n445), .A3(new_n256), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n267), .A2(new_n258), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n267), .B2(new_n253), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n407), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT84), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT18), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n448), .ZN(new_n452));
  INV_X1    g0252(.A(new_n407), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT18), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(KEYINPUT18), .A3(new_n453), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT84), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n451), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(G200), .B1(new_n394), .B2(new_n397), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n403), .A2(G190), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n446), .B(new_n448), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT17), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n386), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G107), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n442), .B2(new_n443), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT6), .ZN(new_n468));
  XNOR2_X1  g0268(.A(G97), .B(G107), .ZN(new_n469));
  NAND2_X1  g0269(.A1(KEYINPUT6), .A2(G97), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT85), .B1(new_n470), .B2(G107), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(new_n466), .A3(KEYINPUT6), .A4(G97), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n468), .A2(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n474), .A2(new_n212), .B1(new_n288), .B2(new_n358), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n256), .B1(new_n467), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n253), .A2(new_n223), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n251), .A2(G33), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n252), .A2(new_n478), .A3(new_n211), .A4(new_n255), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n479), .B2(new_n223), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT88), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT88), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n476), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n273), .A2(G1), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  AND2_X1   g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(G274), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n488), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n293), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(new_n224), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n282), .A2(new_n284), .A3(G244), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n365), .A2(new_n367), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n494), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n493), .B1(new_n501), .B2(new_n294), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT87), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n502), .A2(KEYINPUT87), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n378), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n297), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n486), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n501), .A2(new_n294), .ZN(new_n509));
  INV_X1    g0309(.A(new_n493), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G190), .A3(new_n503), .ZN(new_n514));
  INV_X1    g0314(.A(new_n482), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT86), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n511), .B2(G200), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n502), .A2(KEYINPUT86), .A3(new_n375), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n514), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n362), .A2(G20), .A3(new_n336), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT19), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n212), .B1(new_n316), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n221), .A2(new_n223), .A3(new_n466), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n521), .B1(new_n316), .B2(G20), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n256), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n355), .A2(new_n253), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n479), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(G87), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n487), .A2(G274), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n487), .A2(new_n222), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n293), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n496), .A2(new_n364), .B1(new_n281), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT89), .B1(new_n368), .B2(new_n312), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT89), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n285), .A2(new_n538), .A3(G238), .A4(new_n286), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G190), .B(new_n534), .C1(new_n540), .C2(new_n293), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n531), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n534), .B1(new_n540), .B2(new_n293), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n378), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n297), .B(new_n534), .C1(new_n540), .C2(new_n293), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n527), .B(new_n528), .C1(new_n355), .C2(new_n479), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n542), .A2(new_n544), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT90), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n508), .A2(new_n519), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n508), .A2(new_n549), .A3(new_n519), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT90), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n334), .A2(G20), .A3(new_n466), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n554), .A2(KEYINPUT25), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(KEYINPUT25), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n466), .C2(new_n479), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n285), .A2(new_n212), .A3(G87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT22), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT22), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n285), .A2(new_n561), .A3(new_n212), .A4(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n281), .A2(new_n535), .A3(G20), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n212), .B2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n466), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(KEYINPUT24), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n256), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT24), .B1(new_n563), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n558), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT94), .B1(new_n368), .B2(new_n222), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT94), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n285), .A2(new_n574), .A3(G250), .A4(new_n286), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G294), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n285), .A2(G257), .A3(G1698), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n573), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n294), .ZN(new_n579));
  INV_X1    g0379(.A(new_n492), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G264), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n490), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n582), .A2(new_n297), .A3(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n578), .A2(new_n294), .B1(G264), .B2(new_n580), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n378), .B1(new_n585), .B2(new_n490), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n572), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT95), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n572), .ZN(new_n590));
  AOI21_X1  g0390(.A(G200), .B1(new_n585), .B2(new_n490), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n585), .A2(new_n490), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(G190), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n572), .B(KEYINPUT95), .C1(new_n584), .C2(new_n586), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n589), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OR3_X1    g0396(.A1(new_n479), .A2(KEYINPUT91), .A3(new_n535), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT91), .B1(new_n479), .B2(new_n535), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n535), .B2(new_n253), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n281), .A2(G97), .ZN(new_n600));
  AOI21_X1  g0400(.A(G20), .B1(new_n600), .B2(new_n500), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n212), .A2(new_n535), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n256), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n362), .A2(G303), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n368), .B2(new_n224), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n285), .A2(G264), .A3(G1698), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n294), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n583), .B1(new_n580), .B2(G270), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n378), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n606), .A2(new_n612), .A3(KEYINPUT21), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT92), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(new_n611), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n606), .A2(new_n614), .A3(new_n616), .A4(G179), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n599), .A2(new_n605), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n610), .A2(new_n611), .A3(G179), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT92), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n613), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n616), .A2(G200), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n615), .A2(G190), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n618), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI211_X1 g0424(.A(KEYINPUT93), .B(KEYINPUT21), .C1(new_n606), .C2(new_n612), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT21), .B1(new_n606), .B2(new_n612), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT93), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n621), .B(new_n624), .C1(new_n625), .C2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n596), .A2(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n465), .A2(new_n551), .A3(new_n553), .A4(new_n630), .ZN(G372));
  NAND4_X1  g0431(.A1(new_n508), .A2(new_n519), .A3(new_n594), .A4(new_n549), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n628), .A2(new_n625), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n621), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n632), .B1(new_n634), .B2(new_n587), .ZN(new_n635));
  INV_X1    g0435(.A(new_n549), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT26), .B1(new_n636), .B2(new_n508), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n548), .A2(new_n545), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n506), .A2(new_n507), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(new_n482), .A3(new_n549), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n637), .B(new_n638), .C1(KEYINPUT26), .C2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n465), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT96), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT96), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n456), .A2(new_n457), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n384), .A2(new_n381), .A3(new_n382), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n351), .B1(new_n331), .B2(new_n347), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n646), .B1(new_n649), .B2(new_n464), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n306), .A2(new_n307), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n300), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n644), .A2(new_n645), .A3(new_n652), .ZN(G369));
  OR3_X1    g0453(.A1(new_n335), .A2(KEYINPUT27), .A3(G20), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT27), .B1(new_n335), .B2(G20), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n634), .A2(new_n606), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n658), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n629), .B1(new_n618), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G330), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n589), .A2(new_n595), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n666), .B(new_n594), .C1(new_n590), .C2(new_n660), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n587), .B2(new_n660), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n634), .A2(new_n658), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n671), .A2(new_n667), .B1(new_n587), .B2(new_n658), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n670), .A2(new_n672), .ZN(G399));
  NOR2_X1   g0473(.A1(new_n208), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G1), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n221), .A2(new_n223), .A3(new_n466), .A4(new_n535), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n676), .A2(new_n677), .B1(new_n216), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n630), .A2(new_n551), .A3(new_n553), .A4(new_n660), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT31), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n504), .A2(new_n505), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n582), .A2(new_n619), .A3(new_n543), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(KEYINPUT30), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n616), .A2(new_n502), .A3(G179), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n685), .A2(new_n543), .A3(new_n592), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT30), .B1(new_n682), .B2(new_n683), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n681), .B1(new_n689), .B2(new_n658), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n680), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n689), .A2(new_n681), .A3(new_n658), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n660), .B1(new_n641), .B2(new_n635), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n638), .B(KEYINPUT97), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n508), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT26), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(new_n703), .A3(new_n549), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT98), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n699), .A2(KEYINPUT98), .A3(new_n704), .A4(new_n700), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n634), .A2(new_n666), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(new_n632), .ZN(new_n708));
  OAI211_X1 g0508(.A(KEYINPUT29), .B(new_n660), .C1(new_n705), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n695), .B1(new_n698), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n679), .B1(new_n710), .B2(G1), .ZN(G364));
  NOR2_X1   g0511(.A1(new_n333), .A2(G20), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G45), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n675), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n714), .A2(KEYINPUT99), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(KEYINPUT99), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n664), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n662), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n211), .B1(G20), .B2(new_n378), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n362), .A2(new_n207), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n245), .A2(G45), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n216), .A2(new_n273), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n285), .A2(new_n207), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT100), .ZN(new_n735));
  XNOR2_X1  g0535(.A(G355), .B(KEYINPUT101), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n735), .A2(new_n736), .B1(new_n535), .B2(new_n208), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT102), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n729), .B1(new_n733), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n212), .A2(G190), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G179), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(KEYINPUT103), .B(G159), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT32), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n297), .A2(new_n375), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n740), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n297), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n740), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G68), .A2(new_n748), .B1(new_n751), .B2(G77), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n212), .A2(new_n302), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n746), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n745), .B(new_n752), .C1(new_n243), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n375), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n740), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n466), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n753), .A2(new_n749), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n758), .B1(new_n266), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n753), .A2(new_n756), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n362), .B1(new_n763), .B2(G87), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n741), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n761), .B(new_n764), .C1(new_n223), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n754), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G326), .A2(new_n769), .B1(new_n760), .B2(G322), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  XOR2_X1   g0571(.A(KEYINPUT33), .B(G317), .Z(new_n772));
  OAI221_X1 g0572(.A(new_n770), .B1(new_n771), .B2(new_n750), .C1(new_n747), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n742), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G303), .A2(new_n763), .B1(new_n774), .B2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(new_n757), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n285), .B1(new_n776), .B2(G283), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n775), .B(new_n777), .C1(new_n778), .C2(new_n767), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n755), .A2(new_n768), .B1(new_n773), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n717), .B1(new_n780), .B2(new_n728), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n739), .A2(new_n781), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n720), .A2(new_n722), .B1(new_n727), .B2(new_n782), .ZN(G396));
  NOR2_X1   g0583(.A1(new_n660), .A2(new_n360), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n647), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n385), .B2(new_n784), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n696), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n695), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n718), .B1(new_n695), .B2(new_n788), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n786), .A2(new_n723), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n728), .A2(G77), .A3(new_n723), .ZN(new_n793));
  INV_X1    g0593(.A(new_n743), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n769), .A2(G137), .B1(new_n751), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G143), .ZN(new_n796));
  INV_X1    g0596(.A(G150), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(new_n796), .B2(new_n759), .C1(new_n797), .C2(new_n747), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT34), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n285), .B1(new_n762), .B2(new_n243), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n757), .A2(new_n336), .B1(new_n742), .B2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n802), .B(new_n804), .C1(new_n266), .C2(new_n766), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n800), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G303), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n754), .A2(new_n807), .B1(new_n750), .B2(new_n535), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G283), .B2(new_n748), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT104), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n362), .B1(new_n759), .B2(new_n778), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G97), .B2(new_n766), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G107), .A2(new_n763), .B1(new_n776), .B2(G87), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(new_n771), .C2(new_n742), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n806), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n717), .B(new_n793), .C1(new_n815), .C2(new_n728), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G384));
  INV_X1    g0618(.A(new_n474), .ZN(new_n819));
  OAI211_X1 g0619(.A(G116), .B(new_n213), .C1(new_n819), .C2(KEYINPUT35), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(KEYINPUT35), .B2(new_n819), .ZN(new_n821));
  XOR2_X1   g0621(.A(KEYINPUT105), .B(KEYINPUT36), .Z(new_n822));
  XNOR2_X1  g0622(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n216), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n824), .B(G77), .C1(new_n336), .C2(new_n265), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n201), .A2(G68), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n251), .B(G13), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n347), .A2(new_n658), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n348), .A2(new_n351), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n351), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n347), .B(new_n658), .C1(new_n831), .C2(new_n331), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n786), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n691), .A2(new_n692), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT40), .ZN(new_n836));
  INV_X1    g0636(.A(new_n656), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n452), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n454), .A2(new_n838), .A3(new_n462), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n435), .A2(new_n256), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n416), .A2(new_n417), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n336), .B1(new_n842), .B2(new_n430), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n438), .B1(new_n843), .B2(new_n433), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT16), .B1(new_n844), .B2(new_n419), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n448), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT106), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n434), .A2(new_n424), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n433), .B1(new_n432), .B2(G68), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n436), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n256), .A3(new_n435), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(KEYINPUT106), .A3(new_n448), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n848), .A2(new_n453), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n848), .A2(new_n837), .A3(new_n853), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n855), .A3(new_n462), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n840), .B1(new_n856), .B2(KEYINPUT37), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n454), .A2(KEYINPUT84), .A3(new_n455), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n450), .B1(new_n449), .B2(KEYINPUT18), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n449), .A2(KEYINPUT18), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n462), .B(KEYINPUT17), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n855), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n857), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n646), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n452), .B(new_n837), .C1(new_n866), .C2(new_n464), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n839), .B(KEYINPUT37), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n836), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(new_n840), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n855), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n459), .B2(new_n464), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT38), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n835), .B1(new_n877), .B2(new_n865), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT107), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(new_n462), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n852), .A2(KEYINPUT106), .A3(new_n448), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT106), .B1(new_n852), .B2(new_n448), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n883), .B1(new_n886), .B2(new_n837), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n882), .B1(new_n887), .B2(new_n854), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n876), .B(KEYINPUT38), .C1(new_n888), .C2(new_n840), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n864), .B1(new_n857), .B2(new_n863), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n834), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT107), .B1(new_n891), .B2(KEYINPUT40), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n871), .B1(new_n881), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n465), .A2(new_n693), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n893), .B(new_n894), .Z(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n663), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n348), .A2(new_n658), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n870), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n889), .A2(new_n890), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT39), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n901), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n648), .A2(new_n660), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n696), .B2(new_n786), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n832), .A2(new_n830), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n904), .A2(new_n908), .B1(new_n646), .B2(new_n837), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n709), .A2(new_n465), .A3(new_n698), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n652), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n910), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n896), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n896), .A2(new_n913), .B1(new_n251), .B2(new_n712), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n828), .B1(new_n915), .B2(new_n916), .ZN(G367));
  OAI211_X1 g0717(.A(new_n508), .B(new_n519), .C1(new_n515), .C2(new_n660), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n639), .A2(new_n482), .A3(new_n658), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OR3_X1    g0721(.A1(new_n669), .A2(new_n671), .A3(new_n921), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n922), .A2(KEYINPUT42), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n508), .B1(new_n921), .B2(new_n666), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n660), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(KEYINPUT42), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n531), .A2(new_n660), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n549), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n638), .B2(new_n928), .ZN(new_n930));
  XNOR2_X1  g0730(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(KEYINPUT43), .B2(new_n930), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n923), .A2(new_n925), .A3(new_n926), .A4(new_n932), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n670), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n936), .B1(new_n937), .B2(new_n921), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n934), .A2(new_n670), .A3(new_n920), .A4(new_n935), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n674), .B(KEYINPUT41), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n669), .A2(new_n671), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n671), .A2(new_n667), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT110), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n671), .A2(new_n667), .A3(KEYINPUT110), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n664), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n710), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n672), .A2(new_n921), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT44), .Z(new_n951));
  NOR2_X1   g0751(.A1(new_n672), .A2(new_n921), .ZN(new_n952));
  XNOR2_X1  g0752(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n951), .A2(new_n937), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n670), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n940), .B1(new_n958), .B2(new_n710), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n713), .A2(G1), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n938), .B(new_n939), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n239), .A2(new_n730), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n729), .B1(new_n207), .B2(new_n355), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n717), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G150), .A2(new_n760), .B1(new_n748), .B2(new_n794), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n776), .A2(G77), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(new_n201), .C2(new_n750), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n767), .A2(new_n336), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n285), .B1(new_n754), .B2(new_n796), .ZN(new_n970));
  INV_X1    g0770(.A(G137), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n762), .A2(new_n265), .B1(new_n742), .B2(new_n971), .ZN(new_n972));
  NOR4_X1   g0772(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT112), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n767), .A2(new_n466), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n762), .A2(new_n535), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n362), .B1(new_n223), .B2(new_n757), .C1(new_n976), .C2(KEYINPUT46), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n975), .B(new_n977), .C1(KEYINPUT46), .C2(new_n976), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G294), .A2(new_n748), .B1(new_n751), .B2(G283), .ZN(new_n979));
  INV_X1    g0779(.A(G317), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(new_n742), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT111), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G311), .A2(new_n769), .B1(new_n760), .B2(G303), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n978), .B(new_n984), .C1(new_n982), .C2(new_n983), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n974), .A2(KEYINPUT47), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n728), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT47), .B1(new_n974), .B2(new_n985), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n965), .B1(new_n987), .B2(new_n988), .C1(new_n930), .C2(new_n726), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n961), .A2(new_n989), .ZN(G387));
  NOR2_X1   g0790(.A1(new_n949), .A2(new_n675), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n710), .B2(new_n947), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n669), .A2(new_n725), .ZN(new_n993));
  INV_X1    g0793(.A(new_n728), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n759), .A2(new_n980), .B1(new_n750), .B2(new_n807), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT115), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(KEYINPUT115), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G322), .A2(new_n769), .B1(new_n748), .B2(G311), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT48), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  INV_X1    g0802(.A(G283), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n767), .A2(new_n1003), .B1(new_n762), .B2(new_n778), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n362), .B1(new_n757), .B2(new_n535), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G326), .B2(new_n774), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n769), .A2(G159), .B1(new_n774), .B2(G150), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n336), .B2(new_n750), .C1(new_n288), .C2(new_n762), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n362), .B(new_n1012), .C1(G97), .C2(new_n776), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n767), .A2(new_n355), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n243), .B2(new_n759), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT114), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1013), .B(new_n1016), .C1(new_n268), .C2(new_n747), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n994), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n236), .A2(G45), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT113), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n356), .A2(new_n243), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT50), .Z(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n677), .C1(G68), .C2(G77), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n730), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n735), .A2(new_n677), .B1(new_n466), .B2(new_n208), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n717), .B(new_n1018), .C1(new_n729), .C2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n947), .A2(new_n960), .B1(new_n993), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n992), .A2(new_n1029), .ZN(G393));
  NAND2_X1  g0830(.A1(new_n957), .A2(new_n955), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n921), .A2(new_n725), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n729), .B1(new_n223), .B2(new_n207), .C1(new_n249), .C2(new_n730), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n718), .A2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n754), .A2(new_n980), .B1(new_n759), .B2(new_n771), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT52), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G303), .A2(new_n748), .B1(new_n774), .B2(G322), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G283), .A2(new_n763), .B1(new_n751), .B2(G294), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n285), .B(new_n758), .C1(G116), .C2(new_n766), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT116), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(G159), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n754), .A2(new_n797), .B1(new_n759), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT51), .Z(new_n1046));
  OAI22_X1  g0846(.A1(new_n762), .A2(new_n336), .B1(new_n742), .B2(new_n796), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n357), .A2(new_n750), .B1(new_n201), .B2(new_n747), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n285), .B1(new_n757), .B2(new_n221), .C1(new_n767), .C2(new_n288), .ZN(new_n1049));
  OR4_X1    g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1043), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1035), .B1(new_n1052), .B2(new_n728), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1032), .A2(new_n960), .B1(new_n1033), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1031), .A2(new_n948), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n958), .A3(new_n674), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(G390));
  INV_X1    g0857(.A(new_n907), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n694), .B2(new_n786), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n660), .B1(new_n705), .B2(new_n708), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n905), .B1(new_n1060), .B2(new_n786), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n835), .A2(G330), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n906), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n465), .A2(G330), .A3(new_n693), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n911), .A2(new_n1065), .A3(new_n652), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1061), .A2(new_n907), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n898), .C1(new_n865), .C2(new_n869), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n908), .A2(new_n898), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n900), .A2(new_n902), .A3(new_n1070), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1069), .A2(new_n1071), .A3(new_n1062), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1062), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1067), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1071), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n897), .B(new_n870), .C1(new_n1061), .C2(new_n907), .ZN(new_n1076));
  OAI211_X1 g0876(.A(G330), .B(new_n835), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1069), .A2(new_n1071), .A3(new_n1062), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1074), .A2(new_n674), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n728), .A2(new_n723), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n717), .B1(new_n268), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(G128), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n285), .B1(new_n754), .B2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT54), .B(G143), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n747), .A2(new_n971), .B1(new_n750), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1085), .B(new_n1087), .C1(G159), .C2(new_n766), .ZN(new_n1088));
  INV_X1    g0888(.A(G125), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n742), .A2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n759), .A2(new_n803), .B1(new_n757), .B2(new_n201), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT53), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n762), .B2(new_n797), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n763), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1090), .B(new_n1091), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n362), .B1(new_n762), .B2(new_n221), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n757), .A2(new_n336), .B1(new_n742), .B2(new_n778), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(G77), .C2(new_n766), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n754), .A2(new_n1003), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n747), .A2(new_n466), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n759), .A2(new_n535), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n750), .A2(new_n223), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1088), .A2(new_n1095), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1083), .B1(new_n1104), .B2(new_n994), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n900), .A2(new_n902), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n723), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n960), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1081), .A2(new_n1109), .ZN(G378));
  INV_X1    g0910(.A(new_n910), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n881), .A2(new_n892), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n871), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n308), .B(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n271), .A2(new_n656), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT55), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1115), .B(new_n1117), .Z(new_n1118));
  AND4_X1   g0918(.A1(G330), .A2(new_n1112), .A3(new_n1113), .A4(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n893), .B2(G330), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1111), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT119), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1112), .A2(G330), .A3(new_n1113), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1118), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n893), .A2(G330), .A3(new_n1118), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n910), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1121), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1125), .A2(KEYINPUT119), .A3(new_n910), .A4(new_n1126), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n960), .A3(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n281), .B(new_n272), .C1(new_n757), .C2(new_n743), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n754), .A2(new_n1089), .B1(new_n747), .B2(new_n803), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n751), .A2(G137), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n1084), .B2(new_n759), .C1(new_n762), .C2(new_n1086), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(G150), .C2(new_n766), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(KEYINPUT59), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1131), .B(new_n1137), .C1(G124), .C2(new_n774), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(KEYINPUT59), .B2(new_n1136), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G116), .A2(new_n769), .B1(new_n776), .B2(new_n266), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n288), .B2(new_n762), .C1(new_n223), .C2(new_n747), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n285), .A2(G41), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n466), .B2(new_n759), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n750), .A2(new_n355), .B1(new_n742), .B2(new_n1003), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1141), .A2(new_n969), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(KEYINPUT58), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(KEYINPUT58), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1142), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(new_n243), .C1(G33), .C2(G41), .ZN(new_n1149));
  AND4_X1   g0949(.A1(new_n1139), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT117), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n994), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1151), .B2(new_n1150), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n717), .B1(new_n201), .B2(new_n1082), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1153), .B(new_n1154), .C1(new_n1118), .C2(new_n724), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1130), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1066), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1080), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1128), .A2(new_n1129), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(KEYINPUT120), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n1080), .B2(new_n1157), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n675), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT120), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1156), .B1(new_n1165), .B2(new_n1166), .ZN(G375));
  OR2_X1    g0967(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1066), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT121), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n940), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n1067), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n960), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G150), .A2(new_n751), .B1(new_n774), .B2(G128), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n1044), .B2(new_n762), .C1(new_n747), .C2(new_n1086), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G132), .A2(new_n769), .B1(new_n760), .B2(G137), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n362), .B1(new_n776), .B2(new_n266), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n243), .C2(new_n767), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G97), .A2(new_n763), .B1(new_n774), .B2(G303), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n466), .B2(new_n750), .C1(new_n778), .C2(new_n754), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G116), .A2(new_n748), .B1(new_n760), .B2(G283), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1182), .A2(new_n1014), .A3(new_n362), .A4(new_n967), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1176), .A2(new_n1179), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n728), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n717), .B1(new_n336), .B2(new_n1082), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n907), .C2(new_n724), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1174), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1172), .A2(new_n1189), .ZN(G381));
  OR2_X1    g0990(.A1(G375), .A2(G378), .ZN(new_n1191));
  INV_X1    g0991(.A(G396), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n992), .A2(new_n1192), .A3(new_n1029), .ZN(new_n1193));
  OR4_X1    g0993(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1193), .ZN(new_n1194));
  OR3_X1    g0994(.A1(new_n1191), .A2(G381), .A3(new_n1194), .ZN(G407));
  OAI211_X1 g0995(.A(G407), .B(G213), .C1(G343), .C2(new_n1191), .ZN(G409));
  NAND2_X1  g0996(.A1(new_n657), .A2(G213), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1128), .A2(new_n1171), .A3(new_n1129), .A4(new_n1158), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1155), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1163), .B2(new_n960), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(G378), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT122), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT122), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1205), .B(G378), .C1(new_n1199), .C2(new_n1201), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G378), .B(new_n1156), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1198), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1067), .A2(KEYINPUT60), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1170), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1169), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n675), .B1(new_n1212), .B2(KEYINPUT60), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G384), .B1(new_n1214), .B2(new_n1189), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n817), .B(new_n1188), .C1(new_n1211), .C2(new_n1213), .ZN(new_n1216));
  OAI211_X1 g1016(.A(G2897), .B(new_n1198), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1189), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n817), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1214), .A2(G384), .A3(new_n1189), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1198), .A2(G2897), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1217), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT63), .B1(new_n1209), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1197), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1209), .A2(KEYINPUT63), .A3(new_n1226), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT61), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G390), .B1(new_n961), .B2(new_n989), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n961), .A2(new_n989), .A3(G390), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(G393), .A2(G396), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1193), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1235), .A2(KEYINPUT123), .A3(new_n1193), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1234), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1233), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1232), .B1(new_n1241), .B2(KEYINPUT125), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT125), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1238), .A2(new_n1239), .B1(new_n1231), .B2(new_n1243), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1240), .A2(KEYINPUT124), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT124), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1234), .A2(new_n1246), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1248), .ZN(new_n1249));
  XOR2_X1   g1049(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1209), .B2(new_n1223), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT127), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT62), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1227), .A2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1209), .A2(new_n1252), .A3(new_n1253), .A4(new_n1226), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1251), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1249), .B1(new_n1259), .B2(new_n1248), .ZN(G405));
  NAND2_X1  g1060(.A1(new_n1240), .A2(KEYINPUT124), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1244), .A2(new_n1242), .ZN(new_n1262));
  AND4_X1   g1062(.A1(new_n1226), .A2(new_n1261), .A3(new_n1247), .A4(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1226), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(G375), .B(G378), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1265), .B(new_n1266), .ZN(G402));
endmodule


