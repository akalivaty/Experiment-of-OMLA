

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U551 ( .A1(n596), .A2(n976), .ZN(n597) );
  NOR2_X2 U552 ( .A1(G164), .A2(G1384), .ZN(n683) );
  NOR2_X1 U553 ( .A1(n665), .A2(n666), .ZN(n641) );
  NOR2_X1 U554 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  AND2_X1 U555 ( .A1(n676), .A2(n675), .ZN(n678) );
  AND2_X1 U556 ( .A1(n683), .A2(n681), .ZN(n615) );
  XNOR2_X1 U557 ( .A(n584), .B(n583), .ZN(n596) );
  NAND2_X1 U558 ( .A1(n680), .A2(n679), .ZN(n687) );
  INV_X1 U559 ( .A(KEYINPUT33), .ZN(n679) );
  NOR2_X1 U560 ( .A1(G543), .A2(G651), .ZN(n780) );
  NOR2_X1 U561 ( .A1(n578), .A2(n577), .ZN(n755) );
  AND2_X1 U562 ( .A1(n686), .A2(n514), .ZN(n513) );
  OR2_X1 U563 ( .A1(n685), .A2(n696), .ZN(n514) );
  XNOR2_X1 U564 ( .A(n580), .B(KEYINPUT26), .ZN(n582) );
  INV_X1 U565 ( .A(KEYINPUT97), .ZN(n583) );
  INV_X1 U566 ( .A(KEYINPUT99), .ZN(n640) );
  NOR2_X1 U567 ( .A1(G168), .A2(n644), .ZN(n645) );
  NAND2_X1 U568 ( .A1(G8), .A2(n655), .ZN(n654) );
  BUF_X1 U569 ( .A(n654), .Z(n696) );
  XNOR2_X1 U570 ( .A(n579), .B(KEYINPUT87), .ZN(n681) );
  INV_X1 U571 ( .A(KEYINPUT64), .ZN(n677) );
  XNOR2_X1 U572 ( .A(n678), .B(n677), .ZN(n680) );
  NOR2_X1 U573 ( .A1(G651), .A2(n533), .ZN(n781) );
  BUF_X1 U574 ( .A(n574), .Z(n878) );
  NOR2_X2 U575 ( .A1(n533), .A2(n532), .ZN(n784) );
  INV_X1 U576 ( .A(KEYINPUT40), .ZN(n753) );
  BUF_X1 U577 ( .A(n755), .Z(G160) );
  INV_X1 U578 ( .A(G651), .ZN(n532) );
  NOR2_X1 U579 ( .A1(G543), .A2(n532), .ZN(n516) );
  XNOR2_X1 U580 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n786) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n533) );
  NAND2_X1 U583 ( .A1(G49), .A2(n781), .ZN(n518) );
  NAND2_X1 U584 ( .A1(G74), .A2(G651), .ZN(n517) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U586 ( .A1(n786), .A2(n519), .ZN(n521) );
  NAND2_X1 U587 ( .A1(n533), .A2(G87), .ZN(n520) );
  NAND2_X1 U588 ( .A1(n521), .A2(n520), .ZN(G288) );
  XOR2_X1 U589 ( .A(KEYINPUT17), .B(n522), .Z(n574) );
  NAND2_X1 U590 ( .A1(G138), .A2(n878), .ZN(n524) );
  INV_X1 U591 ( .A(G2104), .ZN(n525) );
  NOR2_X1 U592 ( .A1(G2105), .A2(n525), .ZN(n569) );
  BUF_X1 U593 ( .A(n569), .Z(n879) );
  NAND2_X1 U594 ( .A1(G102), .A2(n879), .ZN(n523) );
  NAND2_X1 U595 ( .A1(n524), .A2(n523), .ZN(n529) );
  AND2_X1 U596 ( .A1(n525), .A2(G2105), .ZN(n882) );
  NAND2_X1 U597 ( .A1(G126), .A2(n882), .ZN(n527) );
  AND2_X1 U598 ( .A1(G2104), .A2(G2105), .ZN(n883) );
  NAND2_X1 U599 ( .A1(G114), .A2(n883), .ZN(n526) );
  NAND2_X1 U600 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U601 ( .A1(n529), .A2(n528), .ZN(G164) );
  NAND2_X1 U602 ( .A1(G52), .A2(n781), .ZN(n531) );
  NAND2_X1 U603 ( .A1(G64), .A2(n786), .ZN(n530) );
  NAND2_X1 U604 ( .A1(n531), .A2(n530), .ZN(n538) );
  NAND2_X1 U605 ( .A1(G77), .A2(n784), .ZN(n535) );
  NAND2_X1 U606 ( .A1(G90), .A2(n780), .ZN(n534) );
  NAND2_X1 U607 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U608 ( .A(KEYINPUT9), .B(n536), .Z(n537) );
  NOR2_X1 U609 ( .A1(n538), .A2(n537), .ZN(G171) );
  INV_X1 U610 ( .A(G171), .ZN(G301) );
  NAND2_X1 U611 ( .A1(n780), .A2(G89), .ZN(n539) );
  XNOR2_X1 U612 ( .A(n539), .B(KEYINPUT4), .ZN(n541) );
  NAND2_X1 U613 ( .A1(G76), .A2(n784), .ZN(n540) );
  NAND2_X1 U614 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U615 ( .A(n542), .B(KEYINPUT5), .ZN(n547) );
  NAND2_X1 U616 ( .A1(G51), .A2(n781), .ZN(n544) );
  NAND2_X1 U617 ( .A1(G63), .A2(n786), .ZN(n543) );
  NAND2_X1 U618 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U619 ( .A(KEYINPUT6), .B(n545), .Z(n546) );
  NAND2_X1 U620 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U621 ( .A(n548), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U623 ( .A1(G50), .A2(n781), .ZN(n550) );
  NAND2_X1 U624 ( .A1(G62), .A2(n786), .ZN(n549) );
  NAND2_X1 U625 ( .A1(n550), .A2(n549), .ZN(n553) );
  NAND2_X1 U626 ( .A1(n780), .A2(G88), .ZN(n551) );
  XOR2_X1 U627 ( .A(KEYINPUT82), .B(n551), .Z(n552) );
  NOR2_X1 U628 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U629 ( .A1(n784), .A2(G75), .ZN(n554) );
  NAND2_X1 U630 ( .A1(n555), .A2(n554), .ZN(G303) );
  NAND2_X1 U631 ( .A1(G48), .A2(n781), .ZN(n557) );
  NAND2_X1 U632 ( .A1(G61), .A2(n786), .ZN(n556) );
  NAND2_X1 U633 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U634 ( .A1(n784), .A2(G73), .ZN(n558) );
  XOR2_X1 U635 ( .A(KEYINPUT2), .B(n558), .Z(n559) );
  NOR2_X1 U636 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U637 ( .A1(n780), .A2(G86), .ZN(n561) );
  NAND2_X1 U638 ( .A1(n562), .A2(n561), .ZN(G305) );
  NAND2_X1 U639 ( .A1(G47), .A2(n781), .ZN(n564) );
  NAND2_X1 U640 ( .A1(G60), .A2(n786), .ZN(n563) );
  NAND2_X1 U641 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U642 ( .A1(G72), .A2(n784), .ZN(n566) );
  NAND2_X1 U643 ( .A1(G85), .A2(n780), .ZN(n565) );
  NAND2_X1 U644 ( .A1(n566), .A2(n565), .ZN(n567) );
  OR2_X1 U645 ( .A1(n568), .A2(n567), .ZN(G290) );
  NOR2_X1 U646 ( .A1(G1976), .A2(G288), .ZN(n966) );
  NAND2_X1 U647 ( .A1(n569), .A2(G101), .ZN(n570) );
  XOR2_X1 U648 ( .A(n570), .B(KEYINPUT23), .Z(n572) );
  NAND2_X1 U649 ( .A1(n882), .A2(G125), .ZN(n571) );
  NAND2_X1 U650 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U651 ( .A(n573), .B(KEYINPUT66), .ZN(n578) );
  NAND2_X1 U652 ( .A1(G137), .A2(n574), .ZN(n576) );
  NAND2_X1 U653 ( .A1(G113), .A2(n883), .ZN(n575) );
  NAND2_X1 U654 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U655 ( .A1(n755), .A2(G40), .ZN(n579) );
  NAND2_X1 U656 ( .A1(n615), .A2(G1996), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n683), .A2(n681), .ZN(n655) );
  NAND2_X1 U658 ( .A1(G1341), .A2(n655), .ZN(n581) );
  NAND2_X1 U659 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n780), .A2(G81), .ZN(n585) );
  XNOR2_X1 U661 ( .A(KEYINPUT12), .B(n585), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n784), .A2(G68), .ZN(n586) );
  XOR2_X1 U663 ( .A(KEYINPUT73), .B(n586), .Z(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U665 ( .A(KEYINPUT13), .B(n589), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G43), .A2(n781), .ZN(n590) );
  XOR2_X1 U667 ( .A(KEYINPUT74), .B(n590), .Z(n593) );
  NAND2_X1 U668 ( .A1(n786), .A2(G56), .ZN(n591) );
  XOR2_X1 U669 ( .A(KEYINPUT14), .B(n591), .Z(n592) );
  NOR2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n976) );
  XNOR2_X1 U672 ( .A(n597), .B(KEYINPUT65), .ZN(n610) );
  NAND2_X1 U673 ( .A1(G66), .A2(n786), .ZN(n604) );
  NAND2_X1 U674 ( .A1(G92), .A2(n780), .ZN(n599) );
  NAND2_X1 U675 ( .A1(G54), .A2(n781), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n784), .A2(G79), .ZN(n600) );
  XOR2_X1 U678 ( .A(KEYINPUT76), .B(n600), .Z(n601) );
  NOR2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT15), .ZN(n606) );
  XOR2_X2 U682 ( .A(KEYINPUT77), .B(n606), .Z(n977) );
  AND2_X1 U683 ( .A1(n615), .A2(G2067), .ZN(n608) );
  AND2_X1 U684 ( .A1(n655), .A2(G1348), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n611) );
  NOR2_X1 U686 ( .A1(n977), .A2(n611), .ZN(n609) );
  NOR2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n613) );
  AND2_X1 U688 ( .A1(n611), .A2(n977), .ZN(n612) );
  NOR2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n614), .B(KEYINPUT98), .ZN(n628) );
  NAND2_X1 U691 ( .A1(n615), .A2(G2072), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT96), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT27), .ZN(n619) );
  INV_X1 U694 ( .A(G1956), .ZN(n990) );
  INV_X1 U695 ( .A(n655), .ZN(n634) );
  NOR2_X1 U696 ( .A1(n990), .A2(n634), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n629) );
  NAND2_X1 U698 ( .A1(G78), .A2(n784), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G91), .A2(n780), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U701 ( .A1(G65), .A2(n786), .ZN(n622) );
  XOR2_X1 U702 ( .A(KEYINPUT69), .B(n622), .Z(n624) );
  NAND2_X1 U703 ( .A1(n781), .A2(G53), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n971) );
  NAND2_X1 U706 ( .A1(n629), .A2(n971), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n632) );
  NOR2_X1 U708 ( .A1(n629), .A2(n971), .ZN(n630) );
  XOR2_X1 U709 ( .A(n630), .B(KEYINPUT28), .Z(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n633), .B(KEYINPUT29), .ZN(n638) );
  XOR2_X1 U712 ( .A(G2078), .B(KEYINPUT25), .Z(n943) );
  NOR2_X1 U713 ( .A1(n943), .A2(n655), .ZN(n636) );
  XOR2_X1 U714 ( .A(G1961), .B(KEYINPUT95), .Z(n999) );
  NOR2_X1 U715 ( .A1(n634), .A2(n999), .ZN(n635) );
  NOR2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n646) );
  NOR2_X1 U717 ( .A1(G301), .A2(n646), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n651) );
  NOR2_X1 U719 ( .A1(n654), .A2(G1966), .ZN(n639) );
  XNOR2_X1 U720 ( .A(n639), .B(KEYINPUT94), .ZN(n665) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n655), .ZN(n666) );
  XNOR2_X1 U722 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n642), .A2(G8), .ZN(n643) );
  XNOR2_X1 U724 ( .A(n643), .B(KEYINPUT30), .ZN(n644) );
  XNOR2_X1 U725 ( .A(n645), .B(KEYINPUT100), .ZN(n648) );
  AND2_X1 U726 ( .A1(n646), .A2(G301), .ZN(n647) );
  NOR2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n649), .B(KEYINPUT31), .ZN(n650) );
  NOR2_X2 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n652), .B(KEYINPUT101), .ZN(n664) );
  AND2_X1 U731 ( .A1(G286), .A2(G8), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n664), .A2(n653), .ZN(n662) );
  INV_X1 U733 ( .A(G8), .ZN(n660) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n696), .ZN(n657) );
  NOR2_X1 U735 ( .A1(G2090), .A2(n655), .ZN(n656) );
  NOR2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n658), .A2(G303), .ZN(n659) );
  OR2_X1 U738 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U740 ( .A(n663), .B(KEYINPUT32), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n664), .B(KEYINPUT102), .ZN(n669) );
  AND2_X1 U742 ( .A1(n666), .A2(G8), .ZN(n667) );
  NOR2_X1 U743 ( .A1(n665), .A2(n667), .ZN(n668) );
  AND2_X1 U744 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U745 ( .A1(n671), .A2(n670), .ZN(n689) );
  NOR2_X1 U746 ( .A1(n966), .A2(n689), .ZN(n673) );
  OR2_X1 U747 ( .A1(G1971), .A2(G303), .ZN(n964) );
  XOR2_X1 U748 ( .A(n964), .B(KEYINPUT103), .Z(n672) );
  NAND2_X1 U749 ( .A1(n673), .A2(n672), .ZN(n676) );
  INV_X1 U750 ( .A(n696), .ZN(n674) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n965) );
  AND2_X1 U752 ( .A1(n674), .A2(n965), .ZN(n675) );
  XOR2_X1 U753 ( .A(G1981), .B(G305), .Z(n961) );
  INV_X1 U754 ( .A(n681), .ZN(n682) );
  NOR2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n748) );
  XNOR2_X1 U756 ( .A(G1986), .B(G290), .ZN(n973) );
  NAND2_X1 U757 ( .A1(n748), .A2(n973), .ZN(n684) );
  XNOR2_X1 U758 ( .A(KEYINPUT88), .B(n684), .ZN(n688) );
  AND2_X1 U759 ( .A1(n961), .A2(n688), .ZN(n686) );
  NAND2_X1 U760 ( .A1(n966), .A2(KEYINPUT33), .ZN(n685) );
  NAND2_X1 U761 ( .A1(n687), .A2(n513), .ZN(n744) );
  INV_X1 U762 ( .A(n688), .ZN(n700) );
  INV_X1 U763 ( .A(n689), .ZN(n692) );
  NOR2_X1 U764 ( .A1(G2090), .A2(G303), .ZN(n690) );
  NAND2_X1 U765 ( .A1(G8), .A2(n690), .ZN(n691) );
  NAND2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n693) );
  AND2_X1 U767 ( .A1(n693), .A2(n696), .ZN(n698) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n694) );
  XOR2_X1 U769 ( .A(n694), .B(KEYINPUT24), .Z(n695) );
  NOR2_X1 U770 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U771 ( .A1(n698), .A2(n697), .ZN(n699) );
  OR2_X1 U772 ( .A1(n700), .A2(n699), .ZN(n742) );
  NAND2_X1 U773 ( .A1(G129), .A2(n882), .ZN(n702) );
  NAND2_X1 U774 ( .A1(G117), .A2(n883), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n879), .A2(G105), .ZN(n703) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n703), .Z(n704) );
  NOR2_X1 U778 ( .A1(n705), .A2(n704), .ZN(n707) );
  NAND2_X1 U779 ( .A1(n878), .A2(G141), .ZN(n706) );
  NAND2_X1 U780 ( .A1(n707), .A2(n706), .ZN(n894) );
  NOR2_X1 U781 ( .A1(G1996), .A2(n894), .ZN(n914) );
  NAND2_X1 U782 ( .A1(G1996), .A2(n894), .ZN(n708) );
  XNOR2_X1 U783 ( .A(KEYINPUT93), .B(n708), .ZN(n718) );
  NAND2_X1 U784 ( .A1(G119), .A2(n882), .ZN(n710) );
  NAND2_X1 U785 ( .A1(G107), .A2(n883), .ZN(n709) );
  NAND2_X1 U786 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U787 ( .A(KEYINPUT91), .B(n711), .ZN(n715) );
  NAND2_X1 U788 ( .A1(G131), .A2(n878), .ZN(n713) );
  NAND2_X1 U789 ( .A1(G95), .A2(n879), .ZN(n712) );
  AND2_X1 U790 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U791 ( .A1(n715), .A2(n714), .ZN(n872) );
  NAND2_X1 U792 ( .A1(G1991), .A2(n872), .ZN(n716) );
  XOR2_X1 U793 ( .A(KEYINPUT92), .B(n716), .Z(n717) );
  NOR2_X1 U794 ( .A1(n718), .A2(n717), .ZN(n746) );
  INV_X1 U795 ( .A(n746), .ZN(n724) );
  NOR2_X1 U796 ( .A1(G1991), .A2(n872), .ZN(n719) );
  XOR2_X1 U797 ( .A(KEYINPUT105), .B(n719), .Z(n927) );
  NOR2_X1 U798 ( .A1(G1986), .A2(G290), .ZN(n720) );
  XNOR2_X1 U799 ( .A(KEYINPUT104), .B(n720), .ZN(n721) );
  NOR2_X1 U800 ( .A1(n927), .A2(n721), .ZN(n722) );
  XNOR2_X1 U801 ( .A(n722), .B(KEYINPUT106), .ZN(n723) );
  NOR2_X1 U802 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U803 ( .A1(n914), .A2(n725), .ZN(n726) );
  XNOR2_X1 U804 ( .A(KEYINPUT39), .B(n726), .ZN(n738) );
  XNOR2_X1 U805 ( .A(G2067), .B(KEYINPUT37), .ZN(n739) );
  NAND2_X1 U806 ( .A1(G128), .A2(n882), .ZN(n728) );
  NAND2_X1 U807 ( .A1(G116), .A2(n883), .ZN(n727) );
  NAND2_X1 U808 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U809 ( .A(n729), .B(KEYINPUT35), .ZN(n735) );
  XNOR2_X1 U810 ( .A(KEYINPUT34), .B(KEYINPUT89), .ZN(n733) );
  NAND2_X1 U811 ( .A1(G140), .A2(n878), .ZN(n731) );
  NAND2_X1 U812 ( .A1(G104), .A2(n879), .ZN(n730) );
  NAND2_X1 U813 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U814 ( .A(n733), .B(n732), .ZN(n734) );
  NAND2_X1 U815 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U816 ( .A(KEYINPUT36), .B(n736), .Z(n873) );
  OR2_X1 U817 ( .A1(n739), .A2(n873), .ZN(n737) );
  XNOR2_X1 U818 ( .A(n737), .B(KEYINPUT90), .ZN(n747) );
  NAND2_X1 U819 ( .A1(n738), .A2(n747), .ZN(n740) );
  NAND2_X1 U820 ( .A1(n873), .A2(n739), .ZN(n923) );
  NAND2_X1 U821 ( .A1(n740), .A2(n923), .ZN(n741) );
  NAND2_X1 U822 ( .A1(n741), .A2(n748), .ZN(n745) );
  AND2_X1 U823 ( .A1(n742), .A2(n745), .ZN(n743) );
  NAND2_X1 U824 ( .A1(n744), .A2(n743), .ZN(n752) );
  INV_X1 U825 ( .A(n745), .ZN(n750) );
  NAND2_X1 U826 ( .A1(n747), .A2(n746), .ZN(n935) );
  NAND2_X1 U827 ( .A1(n935), .A2(n748), .ZN(n749) );
  OR2_X1 U828 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U829 ( .A1(n752), .A2(n751), .ZN(n754) );
  XNOR2_X1 U830 ( .A(n754), .B(n753), .ZN(G329) );
  NAND2_X1 U831 ( .A1(G123), .A2(n882), .ZN(n756) );
  XNOR2_X1 U832 ( .A(n756), .B(KEYINPUT18), .ZN(n763) );
  NAND2_X1 U833 ( .A1(G135), .A2(n878), .ZN(n758) );
  NAND2_X1 U834 ( .A1(G111), .A2(n883), .ZN(n757) );
  NAND2_X1 U835 ( .A1(n758), .A2(n757), .ZN(n761) );
  NAND2_X1 U836 ( .A1(G99), .A2(n879), .ZN(n759) );
  XNOR2_X1 U837 ( .A(KEYINPUT79), .B(n759), .ZN(n760) );
  NOR2_X1 U838 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U839 ( .A1(n763), .A2(n762), .ZN(n925) );
  XNOR2_X1 U840 ( .A(G2096), .B(n925), .ZN(n764) );
  OR2_X1 U841 ( .A1(G2100), .A2(n764), .ZN(G156) );
  INV_X1 U842 ( .A(G69), .ZN(G235) );
  INV_X1 U843 ( .A(G108), .ZN(G238) );
  INV_X1 U844 ( .A(G120), .ZN(G236) );
  INV_X1 U845 ( .A(G132), .ZN(G219) );
  NAND2_X1 U846 ( .A1(G94), .A2(G452), .ZN(n765) );
  XOR2_X1 U847 ( .A(KEYINPUT68), .B(n765), .Z(G173) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n766) );
  XNOR2_X1 U849 ( .A(n766), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U850 ( .A(G223), .ZN(n820) );
  NAND2_X1 U851 ( .A1(n820), .A2(G567), .ZN(n767) );
  XOR2_X1 U852 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  XNOR2_X1 U853 ( .A(G860), .B(KEYINPUT75), .ZN(n772) );
  OR2_X1 U854 ( .A1(n976), .A2(n772), .ZN(G153) );
  NAND2_X1 U855 ( .A1(G868), .A2(G301), .ZN(n769) );
  OR2_X1 U856 ( .A1(n977), .A2(G868), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(G284) );
  XOR2_X1 U858 ( .A(n971), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U859 ( .A1(G299), .A2(G868), .ZN(n771) );
  INV_X1 U860 ( .A(G868), .ZN(n803) );
  NOR2_X1 U861 ( .A1(G286), .A2(n803), .ZN(n770) );
  NOR2_X1 U862 ( .A1(n771), .A2(n770), .ZN(G297) );
  NAND2_X1 U863 ( .A1(n772), .A2(G559), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n773), .A2(n977), .ZN(n774) );
  XNOR2_X1 U865 ( .A(n774), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U866 ( .A1(G868), .A2(n976), .ZN(n775) );
  XNOR2_X1 U867 ( .A(KEYINPUT78), .B(n775), .ZN(n778) );
  NAND2_X1 U868 ( .A1(G868), .A2(n977), .ZN(n776) );
  NOR2_X1 U869 ( .A1(G559), .A2(n776), .ZN(n777) );
  NOR2_X1 U870 ( .A1(n778), .A2(n777), .ZN(G282) );
  NAND2_X1 U871 ( .A1(G559), .A2(n977), .ZN(n779) );
  XNOR2_X1 U872 ( .A(n976), .B(n779), .ZN(n800) );
  NOR2_X1 U873 ( .A1(n800), .A2(G860), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G93), .A2(n780), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G55), .A2(n781), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G80), .A2(n784), .ZN(n785) );
  XNOR2_X1 U878 ( .A(n785), .B(KEYINPUT80), .ZN(n789) );
  NAND2_X1 U879 ( .A1(G67), .A2(n786), .ZN(n787) );
  XOR2_X1 U880 ( .A(KEYINPUT81), .B(n787), .Z(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n802) );
  XOR2_X1 U883 ( .A(n792), .B(n802), .Z(G145) );
  XNOR2_X1 U884 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n794) );
  XNOR2_X1 U885 ( .A(G288), .B(KEYINPUT84), .ZN(n793) );
  XNOR2_X1 U886 ( .A(n794), .B(n793), .ZN(n795) );
  XOR2_X1 U887 ( .A(n802), .B(n795), .Z(n797) );
  XNOR2_X1 U888 ( .A(G305), .B(G299), .ZN(n796) );
  XNOR2_X1 U889 ( .A(n797), .B(n796), .ZN(n798) );
  XNOR2_X1 U890 ( .A(n798), .B(G303), .ZN(n799) );
  XNOR2_X1 U891 ( .A(n799), .B(G290), .ZN(n898) );
  XOR2_X1 U892 ( .A(n800), .B(n898), .Z(n801) );
  NAND2_X1 U893 ( .A1(n801), .A2(G868), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n805), .A2(n804), .ZN(G295) );
  NAND2_X1 U896 ( .A1(G2084), .A2(G2078), .ZN(n806) );
  XOR2_X1 U897 ( .A(KEYINPUT20), .B(n806), .Z(n807) );
  NAND2_X1 U898 ( .A1(G2090), .A2(n807), .ZN(n808) );
  XNOR2_X1 U899 ( .A(KEYINPUT21), .B(n808), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n809), .A2(G2072), .ZN(n810) );
  XOR2_X1 U901 ( .A(KEYINPUT85), .B(n810), .Z(G158) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U903 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  XNOR2_X1 U904 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  NOR2_X1 U905 ( .A1(G220), .A2(G219), .ZN(n811) );
  XOR2_X1 U906 ( .A(KEYINPUT22), .B(n811), .Z(n812) );
  NOR2_X1 U907 ( .A1(G218), .A2(n812), .ZN(n813) );
  NAND2_X1 U908 ( .A1(G96), .A2(n813), .ZN(n910) );
  NAND2_X1 U909 ( .A1(n910), .A2(G2106), .ZN(n818) );
  NOR2_X1 U910 ( .A1(G237), .A2(G236), .ZN(n815) );
  NOR2_X1 U911 ( .A1(G238), .A2(G235), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U913 ( .A(KEYINPUT86), .B(n816), .ZN(n911) );
  NAND2_X1 U914 ( .A1(n911), .A2(G567), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n912) );
  NAND2_X1 U916 ( .A1(G483), .A2(G661), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n912), .A2(n819), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n820), .ZN(G217) );
  NAND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n821) );
  XNOR2_X1 U921 ( .A(KEYINPUT109), .B(n821), .ZN(n822) );
  NAND2_X1 U922 ( .A1(n822), .A2(G661), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U924 ( .A1(n824), .A2(n823), .ZN(G188) );
  XOR2_X1 U925 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  XOR2_X1 U926 ( .A(G2454), .B(G2435), .Z(n826) );
  XNOR2_X1 U927 ( .A(G2438), .B(G2427), .ZN(n825) );
  XNOR2_X1 U928 ( .A(n826), .B(n825), .ZN(n833) );
  XOR2_X1 U929 ( .A(KEYINPUT107), .B(G2446), .Z(n828) );
  XNOR2_X1 U930 ( .A(G2443), .B(G2430), .ZN(n827) );
  XNOR2_X1 U931 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U932 ( .A(n829), .B(G2451), .Z(n831) );
  XNOR2_X1 U933 ( .A(G1348), .B(G1341), .ZN(n830) );
  XNOR2_X1 U934 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U936 ( .A1(n834), .A2(G14), .ZN(n835) );
  XOR2_X1 U937 ( .A(KEYINPUT108), .B(n835), .Z(G401) );
  XOR2_X1 U938 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n837) );
  XNOR2_X1 U939 ( .A(G2678), .B(KEYINPUT43), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2090), .Z(n839) );
  XNOR2_X1 U942 ( .A(G2072), .B(G2067), .ZN(n838) );
  XNOR2_X1 U943 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U944 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U945 ( .A(G2096), .B(G2100), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U947 ( .A(G2084), .B(G2078), .Z(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1986), .B(G1976), .Z(n847) );
  XNOR2_X1 U950 ( .A(G1961), .B(G1956), .ZN(n846) );
  XNOR2_X1 U951 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U952 ( .A(G1991), .B(G1981), .Z(n849) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1996), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U955 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U956 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n855) );
  XOR2_X1 U958 ( .A(G1971), .B(G2474), .Z(n854) );
  XNOR2_X1 U959 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G112), .A2(n883), .ZN(n856) );
  XNOR2_X1 U961 ( .A(n856), .B(KEYINPUT114), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G124), .A2(n882), .ZN(n857) );
  XNOR2_X1 U963 ( .A(n857), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G136), .A2(n878), .ZN(n861) );
  NAND2_X1 U966 ( .A1(G100), .A2(n879), .ZN(n860) );
  NAND2_X1 U967 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U968 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U969 ( .A1(G130), .A2(n882), .ZN(n865) );
  NAND2_X1 U970 ( .A1(G118), .A2(n883), .ZN(n864) );
  NAND2_X1 U971 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G142), .A2(n878), .ZN(n867) );
  NAND2_X1 U973 ( .A1(G106), .A2(n879), .ZN(n866) );
  NAND2_X1 U974 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U975 ( .A(n868), .B(KEYINPUT45), .Z(n869) );
  NOR2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U977 ( .A(n871), .B(n925), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n872), .B(G162), .ZN(n875) );
  XOR2_X1 U979 ( .A(G160), .B(n873), .Z(n874) );
  XNOR2_X1 U980 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n877), .B(n876), .ZN(n896) );
  NAND2_X1 U982 ( .A1(G139), .A2(n878), .ZN(n881) );
  NAND2_X1 U983 ( .A1(G103), .A2(n879), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U985 ( .A1(G127), .A2(n882), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G115), .A2(n883), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n886), .Z(n887) );
  NOR2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n916) );
  XNOR2_X1 U990 ( .A(G164), .B(n916), .ZN(n892) );
  XOR2_X1 U991 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n890) );
  XNOR2_X1 U992 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n889) );
  XNOR2_X1 U993 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U994 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U997 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U998 ( .A(KEYINPUT117), .B(n898), .Z(n900) );
  XNOR2_X1 U999 ( .A(G171), .B(n977), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(G286), .B(n901), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n902), .B(n976), .ZN(n903) );
  NOR2_X1 U1003 ( .A1(n903), .A2(G37), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n904), .B(KEYINPUT118), .ZN(G397) );
  OR2_X1 U1005 ( .A1(n912), .A2(G401), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n909) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(G225) );
  XNOR2_X1 U1011 ( .A(KEYINPUT119), .B(G225), .ZN(G308) );
  NOR2_X1 U1013 ( .A1(n911), .A2(n910), .ZN(G325) );
  INV_X1 U1014 ( .A(G325), .ZN(G261) );
  INV_X1 U1015 ( .A(n912), .ZN(G319) );
  INV_X1 U1016 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1017 ( .A(G2090), .B(G162), .Z(n913) );
  NOR2_X1 U1018 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1019 ( .A(KEYINPUT51), .B(n915), .Z(n933) );
  XOR2_X1 U1020 ( .A(G2072), .B(n916), .Z(n917) );
  XNOR2_X1 U1021 ( .A(KEYINPUT121), .B(n917), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(G164), .B(G2078), .ZN(n918) );
  XNOR2_X1 U1023 ( .A(n918), .B(KEYINPUT122), .ZN(n919) );
  NAND2_X1 U1024 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1025 ( .A(n921), .B(KEYINPUT50), .ZN(n922) );
  XNOR2_X1 U1026 ( .A(n922), .B(KEYINPUT123), .ZN(n924) );
  NAND2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(G160), .B(G2084), .ZN(n926) );
  NAND2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1031 ( .A(KEYINPUT120), .B(n929), .Z(n930) );
  NOR2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n936), .ZN(n937) );
  INV_X1 U1036 ( .A(KEYINPUT55), .ZN(n957) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n957), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n938), .A2(G29), .ZN(n1019) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n952) );
  XOR2_X1 U1040 ( .A(G1991), .B(G25), .Z(n939) );
  NAND2_X1 U1041 ( .A1(n939), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G2072), .B(G33), .ZN(n941) );
  XNOR2_X1 U1043 ( .A(G26), .B(G2067), .ZN(n940) );
  NOR2_X1 U1044 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1045 ( .A(KEYINPUT124), .B(n942), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(n943), .B(G27), .ZN(n945) );
  XNOR2_X1 U1047 ( .A(G32), .B(G1996), .ZN(n944) );
  NOR2_X1 U1048 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n950), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n953) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n953), .ZN(n954) );
  NAND2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1056 ( .A(n957), .B(n956), .ZN(n959) );
  INV_X1 U1057 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n960), .ZN(n1017) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n989) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G168), .ZN(n962) );
  NAND2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1063 ( .A(n963), .B(KEYINPUT57), .ZN(n987) );
  NAND2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(KEYINPUT127), .B(n966), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n967) );
  NAND2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n975) );
  XOR2_X1 U1069 ( .A(n971), .B(G1956), .Z(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n985) );
  XOR2_X1 U1072 ( .A(n976), .B(G1341), .Z(n983) );
  XNOR2_X1 U1073 ( .A(n977), .B(G1348), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(n978), .B(KEYINPUT125), .ZN(n980) );
  XOR2_X1 U1075 ( .A(G1961), .B(G171), .Z(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(KEYINPUT126), .B(n981), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n1015) );
  INV_X1 U1082 ( .A(G16), .ZN(n1013) );
  XNOR2_X1 U1083 ( .A(G20), .B(n990), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1088 ( .A(KEYINPUT59), .B(G1348), .Z(n995) );
  XNOR2_X1 U1089 ( .A(G4), .B(n995), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n998), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n999), .B(G5), .ZN(n1000) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(G24), .B(G1986), .ZN(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XOR2_X1 U1099 ( .A(G1976), .B(G23), .Z(n1006) );
  NAND2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1020), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

