

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(n726), .ZN(n705) );
  NAND2_X2 U554 ( .A1(n676), .A2(n675), .ZN(n726) );
  NOR2_X1 U555 ( .A1(n972), .A2(n689), .ZN(n695) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n703) );
  XNOR2_X1 U557 ( .A(n704), .B(n703), .ZN(n709) );
  XOR2_X1 U558 ( .A(KEYINPUT17), .B(n533), .Z(n866) );
  NOR2_X1 U559 ( .A1(G651), .A2(G543), .ZN(n636) );
  NAND2_X1 U560 ( .A1(G89), .A2(n636), .ZN(n518) );
  XNOR2_X1 U561 ( .A(n518), .B(KEYINPUT72), .ZN(n519) );
  XNOR2_X1 U562 ( .A(n519), .B(KEYINPUT4), .ZN(n522) );
  INV_X1 U563 ( .A(G651), .ZN(n524) );
  XOR2_X1 U564 ( .A(KEYINPUT0), .B(G543), .Z(n616) );
  OR2_X1 U565 ( .A1(n524), .A2(n616), .ZN(n520) );
  XNOR2_X1 U566 ( .A(KEYINPUT65), .B(n520), .ZN(n635) );
  NAND2_X1 U567 ( .A1(G76), .A2(n635), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U569 ( .A(n523), .B(KEYINPUT5), .ZN(n531) );
  NOR2_X1 U570 ( .A1(G543), .A2(n524), .ZN(n525) );
  XOR2_X1 U571 ( .A(KEYINPUT1), .B(n525), .Z(n640) );
  NAND2_X1 U572 ( .A1(G63), .A2(n640), .ZN(n528) );
  NOR2_X1 U573 ( .A1(G651), .A2(n616), .ZN(n526) );
  XNOR2_X1 U574 ( .A(KEYINPUT64), .B(n526), .ZN(n644) );
  NAND2_X1 U575 ( .A1(G51), .A2(n644), .ZN(n527) );
  NAND2_X1 U576 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U577 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U579 ( .A(n532), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U580 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U581 ( .A(G2105), .ZN(n536) );
  AND2_X1 U582 ( .A1(n536), .A2(G2104), .ZN(n865) );
  NAND2_X1 U583 ( .A1(G102), .A2(n865), .ZN(n535) );
  NOR2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  NAND2_X1 U585 ( .A1(G138), .A2(n866), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n540) );
  NOR2_X1 U587 ( .A1(G2104), .A2(n536), .ZN(n869) );
  NAND2_X1 U588 ( .A1(G126), .A2(n869), .ZN(n538) );
  AND2_X1 U589 ( .A1(G2105), .A2(G2104), .ZN(n870) );
  NAND2_X1 U590 ( .A1(G114), .A2(n870), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U592 ( .A1(n540), .A2(n539), .ZN(G164) );
  XNOR2_X1 U593 ( .A(KEYINPUT9), .B(KEYINPUT69), .ZN(n544) );
  NAND2_X1 U594 ( .A1(G90), .A2(n636), .ZN(n542) );
  NAND2_X1 U595 ( .A1(G77), .A2(n635), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U597 ( .A(n544), .B(n543), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n640), .A2(G64), .ZN(n545) );
  XNOR2_X1 U599 ( .A(n545), .B(KEYINPUT68), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G52), .A2(n644), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U602 ( .A1(n549), .A2(n548), .ZN(G171) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U604 ( .A(G132), .ZN(G219) );
  INV_X1 U605 ( .A(G82), .ZN(G220) );
  INV_X1 U606 ( .A(G57), .ZN(G237) );
  INV_X1 U607 ( .A(G108), .ZN(G238) );
  INV_X1 U608 ( .A(G120), .ZN(G236) );
  NAND2_X1 U609 ( .A1(n869), .A2(G125), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G101), .A2(n865), .ZN(n550) );
  XOR2_X1 U611 ( .A(KEYINPUT23), .B(n550), .Z(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G113), .A2(n870), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G137), .A2(n866), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U616 ( .A1(n556), .A2(n555), .ZN(G160) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U619 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n559) );
  INV_X1 U620 ( .A(G223), .ZN(n810) );
  NAND2_X1 U621 ( .A1(G567), .A2(n810), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n559), .B(n558), .ZN(G234) );
  NAND2_X1 U623 ( .A1(G56), .A2(n640), .ZN(n560) );
  XOR2_X1 U624 ( .A(KEYINPUT14), .B(n560), .Z(n566) );
  NAND2_X1 U625 ( .A1(n636), .A2(G81), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G68), .A2(n635), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT13), .B(n564), .Z(n565) );
  NOR2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U631 ( .A1(G43), .A2(n644), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n972) );
  INV_X1 U633 ( .A(G860), .ZN(n586) );
  OR2_X1 U634 ( .A1(n972), .A2(n586), .ZN(G153) );
  XNOR2_X1 U635 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G868), .A2(G301), .ZN(n577) );
  NAND2_X1 U637 ( .A1(G92), .A2(n636), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G66), .A2(n640), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G79), .A2(n635), .ZN(n572) );
  NAND2_X1 U641 ( .A1(G54), .A2(n644), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U644 ( .A(KEYINPUT15), .B(n575), .Z(n960) );
  OR2_X1 U645 ( .A1(n960), .A2(G868), .ZN(n576) );
  NAND2_X1 U646 ( .A1(n577), .A2(n576), .ZN(G284) );
  NAND2_X1 U647 ( .A1(G65), .A2(n640), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G53), .A2(n644), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G91), .A2(n636), .ZN(n581) );
  NAND2_X1 U651 ( .A1(G78), .A2(n635), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n951) );
  INV_X1 U654 ( .A(n951), .ZN(G299) );
  INV_X1 U655 ( .A(G868), .ZN(n657) );
  NOR2_X1 U656 ( .A1(G286), .A2(n657), .ZN(n585) );
  NOR2_X1 U657 ( .A1(G868), .A2(G299), .ZN(n584) );
  NOR2_X1 U658 ( .A1(n585), .A2(n584), .ZN(G297) );
  NAND2_X1 U659 ( .A1(n586), .A2(G559), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n587), .A2(n960), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n588), .B(KEYINPUT16), .ZN(n589) );
  XOR2_X1 U662 ( .A(KEYINPUT73), .B(n589), .Z(G148) );
  NOR2_X1 U663 ( .A1(G868), .A2(n972), .ZN(n590) );
  XNOR2_X1 U664 ( .A(KEYINPUT74), .B(n590), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G868), .A2(n960), .ZN(n591) );
  NOR2_X1 U666 ( .A1(G559), .A2(n591), .ZN(n592) );
  NOR2_X1 U667 ( .A1(n593), .A2(n592), .ZN(G282) );
  NAND2_X1 U668 ( .A1(G111), .A2(n870), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G99), .A2(n865), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G135), .A2(n866), .ZN(n596) );
  XNOR2_X1 U672 ( .A(n596), .B(KEYINPUT76), .ZN(n600) );
  XOR2_X1 U673 ( .A(KEYINPUT75), .B(KEYINPUT18), .Z(n598) );
  NAND2_X1 U674 ( .A1(G123), .A2(n869), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n598), .B(n597), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n986) );
  XNOR2_X1 U678 ( .A(n986), .B(G2096), .ZN(n604) );
  INV_X1 U679 ( .A(G2100), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(G156) );
  NAND2_X1 U681 ( .A1(n960), .A2(G559), .ZN(n647) );
  XNOR2_X1 U682 ( .A(n972), .B(n647), .ZN(n605) );
  NOR2_X1 U683 ( .A1(n605), .A2(G860), .ZN(n612) );
  NAND2_X1 U684 ( .A1(G93), .A2(n636), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G67), .A2(n640), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G80), .A2(n635), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G55), .A2(n644), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n610) );
  OR2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n656) );
  XOR2_X1 U691 ( .A(n612), .B(n656), .Z(G145) );
  NAND2_X1 U692 ( .A1(G651), .A2(G74), .ZN(n614) );
  NAND2_X1 U693 ( .A1(G49), .A2(n644), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U695 ( .A1(n640), .A2(n615), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n616), .A2(G87), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(G288) );
  NAND2_X1 U698 ( .A1(G62), .A2(n640), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G50), .A2(n644), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U701 ( .A(KEYINPUT78), .B(n621), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G88), .A2(n636), .ZN(n622) );
  XNOR2_X1 U703 ( .A(KEYINPUT79), .B(n622), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n635), .A2(G75), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(G303) );
  INV_X1 U707 ( .A(G303), .ZN(G166) );
  NAND2_X1 U708 ( .A1(n640), .A2(G61), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G86), .A2(n636), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G48), .A2(n644), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n635), .A2(G73), .ZN(n629) );
  XOR2_X1 U713 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U716 ( .A(KEYINPUT77), .B(n634), .Z(G305) );
  NAND2_X1 U717 ( .A1(n635), .A2(G72), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n636), .A2(G85), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U720 ( .A(KEYINPUT66), .B(n639), .ZN(n643) );
  NAND2_X1 U721 ( .A1(G60), .A2(n640), .ZN(n641) );
  XNOR2_X1 U722 ( .A(KEYINPUT67), .B(n641), .ZN(n642) );
  NOR2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G47), .A2(n644), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(G290) );
  XOR2_X1 U726 ( .A(KEYINPUT80), .B(n647), .Z(n654) );
  XNOR2_X1 U727 ( .A(KEYINPUT19), .B(n656), .ZN(n648) );
  XNOR2_X1 U728 ( .A(G288), .B(n648), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n951), .B(n649), .ZN(n652) );
  XNOR2_X1 U730 ( .A(G166), .B(n972), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n650), .B(G305), .ZN(n651) );
  XNOR2_X1 U732 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n653), .B(G290), .ZN(n879) );
  XNOR2_X1 U734 ( .A(n654), .B(n879), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n655), .A2(G868), .ZN(n659) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U744 ( .A1(G236), .A2(G238), .ZN(n664) );
  NAND2_X1 U745 ( .A1(G69), .A2(n664), .ZN(n665) );
  NOR2_X1 U746 ( .A1(n665), .A2(G237), .ZN(n666) );
  XNOR2_X1 U747 ( .A(n666), .B(KEYINPUT81), .ZN(n816) );
  NAND2_X1 U748 ( .A1(n816), .A2(G567), .ZN(n671) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U751 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U752 ( .A1(G96), .A2(n669), .ZN(n817) );
  NAND2_X1 U753 ( .A1(n817), .A2(G2106), .ZN(n670) );
  NAND2_X1 U754 ( .A1(n671), .A2(n670), .ZN(n818) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U756 ( .A1(n818), .A2(n672), .ZN(n813) );
  NAND2_X1 U757 ( .A1(n813), .A2(G36), .ZN(G176) );
  NOR2_X2 U758 ( .A1(G164), .A2(G1384), .ZN(n676) );
  NAND2_X1 U759 ( .A1(G160), .A2(G40), .ZN(n674) );
  NOR2_X1 U760 ( .A1(n676), .A2(n674), .ZN(n806) );
  XNOR2_X1 U761 ( .A(G1986), .B(G290), .ZN(n958) );
  NAND2_X1 U762 ( .A1(n806), .A2(n958), .ZN(n673) );
  XOR2_X1 U763 ( .A(KEYINPUT82), .B(n673), .Z(n761) );
  INV_X1 U764 ( .A(n674), .ZN(n675) );
  NAND2_X1 U765 ( .A1(G8), .A2(n726), .ZN(n752) );
  NOR2_X1 U766 ( .A1(G1981), .A2(G305), .ZN(n677) );
  XOR2_X1 U767 ( .A(n677), .B(KEYINPUT89), .Z(n678) );
  XNOR2_X1 U768 ( .A(KEYINPUT24), .B(n678), .ZN(n744) );
  XOR2_X1 U769 ( .A(KEYINPUT96), .B(G1981), .Z(n679) );
  XNOR2_X1 U770 ( .A(G305), .B(n679), .ZN(n963) );
  NAND2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n949) );
  NAND2_X1 U772 ( .A1(n963), .A2(n949), .ZN(n742) );
  NOR2_X1 U773 ( .A1(G2084), .A2(n726), .ZN(n710) );
  NAND2_X1 U774 ( .A1(G8), .A2(n710), .ZN(n724) );
  NOR2_X1 U775 ( .A1(G1966), .A2(n752), .ZN(n722) );
  NAND2_X1 U776 ( .A1(G2072), .A2(n705), .ZN(n680) );
  XNOR2_X1 U777 ( .A(n680), .B(KEYINPUT90), .ZN(n681) );
  XNOR2_X1 U778 ( .A(KEYINPUT27), .B(n681), .ZN(n683) );
  AND2_X1 U779 ( .A1(n726), .A2(G1956), .ZN(n682) );
  NOR2_X1 U780 ( .A1(n683), .A2(n682), .ZN(n698) );
  NOR2_X1 U781 ( .A1(n951), .A2(n698), .ZN(n685) );
  XNOR2_X1 U782 ( .A(KEYINPUT28), .B(KEYINPUT91), .ZN(n684) );
  XNOR2_X1 U783 ( .A(n685), .B(n684), .ZN(n702) );
  AND2_X1 U784 ( .A1(n705), .A2(G1996), .ZN(n686) );
  XOR2_X1 U785 ( .A(n686), .B(KEYINPUT26), .Z(n688) );
  NAND2_X1 U786 ( .A1(n726), .A2(G1341), .ZN(n687) );
  NAND2_X1 U787 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U788 ( .A1(n960), .A2(n695), .ZN(n694) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n726), .ZN(n691) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n705), .ZN(n690) );
  NAND2_X1 U791 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U792 ( .A(KEYINPUT92), .B(n692), .ZN(n693) );
  NAND2_X1 U793 ( .A1(n694), .A2(n693), .ZN(n697) );
  OR2_X1 U794 ( .A1(n960), .A2(n695), .ZN(n696) );
  NAND2_X1 U795 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n951), .A2(n698), .ZN(n699) );
  NAND2_X1 U797 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n704) );
  INV_X1 U799 ( .A(G1961), .ZN(n923) );
  NAND2_X1 U800 ( .A1(n726), .A2(n923), .ZN(n707) );
  XNOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .ZN(n907) );
  NAND2_X1 U802 ( .A1(n705), .A2(n907), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n714) );
  NAND2_X1 U804 ( .A1(n714), .A2(G171), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n720) );
  NOR2_X1 U806 ( .A1(n722), .A2(n710), .ZN(n711) );
  NAND2_X1 U807 ( .A1(G8), .A2(n711), .ZN(n712) );
  XNOR2_X1 U808 ( .A(KEYINPUT30), .B(n712), .ZN(n713) );
  NOR2_X1 U809 ( .A1(G168), .A2(n713), .ZN(n717) );
  NOR2_X1 U810 ( .A1(G171), .A2(n714), .ZN(n715) );
  XOR2_X1 U811 ( .A(KEYINPUT93), .B(n715), .Z(n716) );
  NOR2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U813 ( .A(KEYINPUT31), .B(n718), .Z(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n725) );
  INV_X1 U815 ( .A(n725), .ZN(n721) );
  NOR2_X1 U816 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n736) );
  NAND2_X1 U818 ( .A1(n725), .A2(G286), .ZN(n731) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n752), .ZN(n728) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n726), .ZN(n727) );
  NOR2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U822 ( .A1(n729), .A2(G303), .ZN(n730) );
  NAND2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U824 ( .A(KEYINPUT94), .B(n732), .ZN(n733) );
  NAND2_X1 U825 ( .A1(n733), .A2(G8), .ZN(n734) );
  XNOR2_X1 U826 ( .A(n734), .B(KEYINPUT32), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n748) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n737) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n948) );
  NOR2_X1 U830 ( .A1(n737), .A2(n948), .ZN(n738) );
  NAND2_X1 U831 ( .A1(n748), .A2(n738), .ZN(n740) );
  NOR2_X1 U832 ( .A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U836 ( .A1(n752), .A2(n745), .ZN(n759) );
  NAND2_X1 U837 ( .A1(G8), .A2(G166), .ZN(n746) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n746), .ZN(n747) );
  XNOR2_X1 U839 ( .A(n747), .B(KEYINPUT97), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U841 ( .A1(n750), .A2(n752), .ZN(n757) );
  XNOR2_X1 U842 ( .A(KEYINPUT95), .B(n948), .ZN(n751) );
  NOR2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n754) );
  INV_X1 U844 ( .A(n963), .ZN(n753) );
  NOR2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U846 ( .A1(KEYINPUT33), .A2(n755), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n793) );
  XNOR2_X1 U850 ( .A(G2067), .B(KEYINPUT37), .ZN(n762) );
  XOR2_X1 U851 ( .A(n762), .B(KEYINPUT83), .Z(n803) );
  NAND2_X1 U852 ( .A1(G128), .A2(n869), .ZN(n764) );
  NAND2_X1 U853 ( .A1(G116), .A2(n870), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U855 ( .A(n765), .B(KEYINPUT35), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G104), .A2(n865), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G140), .A2(n866), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U859 ( .A(KEYINPUT34), .B(n768), .Z(n769) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U861 ( .A(n771), .B(KEYINPUT36), .Z(n862) );
  OR2_X1 U862 ( .A1(n803), .A2(n862), .ZN(n987) );
  NAND2_X1 U863 ( .A1(G129), .A2(n869), .ZN(n773) );
  NAND2_X1 U864 ( .A1(G141), .A2(n866), .ZN(n772) );
  NAND2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n865), .A2(G105), .ZN(n774) );
  XOR2_X1 U867 ( .A(KEYINPUT38), .B(n774), .Z(n775) );
  NOR2_X1 U868 ( .A1(n776), .A2(n775), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n870), .A2(G117), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n853) );
  NAND2_X1 U871 ( .A1(G1996), .A2(n853), .ZN(n779) );
  XNOR2_X1 U872 ( .A(n779), .B(KEYINPUT86), .ZN(n788) );
  XOR2_X1 U873 ( .A(KEYINPUT85), .B(G1991), .Z(n908) );
  NAND2_X1 U874 ( .A1(G95), .A2(n865), .ZN(n780) );
  XNOR2_X1 U875 ( .A(n780), .B(KEYINPUT84), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n870), .A2(G107), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U878 ( .A1(G119), .A2(n869), .ZN(n784) );
  NAND2_X1 U879 ( .A1(G131), .A2(n866), .ZN(n783) );
  NAND2_X1 U880 ( .A1(n784), .A2(n783), .ZN(n785) );
  OR2_X1 U881 ( .A1(n786), .A2(n785), .ZN(n857) );
  NAND2_X1 U882 ( .A1(n908), .A2(n857), .ZN(n787) );
  NAND2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U884 ( .A(KEYINPUT87), .B(n789), .Z(n797) );
  INV_X1 U885 ( .A(n797), .ZN(n992) );
  NAND2_X1 U886 ( .A1(n987), .A2(n992), .ZN(n790) );
  NAND2_X1 U887 ( .A1(n790), .A2(n806), .ZN(n791) );
  XNOR2_X1 U888 ( .A(n791), .B(KEYINPUT88), .ZN(n792) );
  NAND2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n808) );
  OR2_X1 U890 ( .A1(n908), .A2(n857), .ZN(n794) );
  XNOR2_X1 U891 ( .A(n794), .B(KEYINPUT99), .ZN(n990) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n795) );
  XNOR2_X1 U893 ( .A(KEYINPUT98), .B(n795), .ZN(n796) );
  NOR2_X1 U894 ( .A1(n990), .A2(n796), .ZN(n798) );
  NOR2_X1 U895 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n853), .ZN(n996) );
  NOR2_X1 U897 ( .A1(n799), .A2(n996), .ZN(n800) );
  XNOR2_X1 U898 ( .A(n800), .B(KEYINPUT39), .ZN(n801) );
  XNOR2_X1 U899 ( .A(n801), .B(KEYINPUT100), .ZN(n802) );
  NAND2_X1 U900 ( .A1(n802), .A2(n987), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n803), .A2(n862), .ZN(n1005) );
  NAND2_X1 U902 ( .A1(n804), .A2(n1005), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U905 ( .A(KEYINPUT40), .B(n809), .ZN(G329) );
  NAND2_X1 U906 ( .A1(n810), .A2(G2106), .ZN(n811) );
  XNOR2_X1 U907 ( .A(n811), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n812) );
  NAND2_X1 U909 ( .A1(G661), .A2(n812), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G3), .A2(G1), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U912 ( .A(KEYINPUT105), .B(n815), .Z(G188) );
  XOR2_X1 U913 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  NOR2_X1 U915 ( .A1(n817), .A2(n816), .ZN(G325) );
  INV_X1 U916 ( .A(G325), .ZN(G261) );
  INV_X1 U917 ( .A(n818), .ZN(G319) );
  XOR2_X1 U918 ( .A(G2100), .B(G2096), .Z(n820) );
  XNOR2_X1 U919 ( .A(KEYINPUT42), .B(G2678), .ZN(n819) );
  XNOR2_X1 U920 ( .A(n820), .B(n819), .ZN(n824) );
  XOR2_X1 U921 ( .A(KEYINPUT43), .B(G2090), .Z(n822) );
  XNOR2_X1 U922 ( .A(G2067), .B(G2072), .ZN(n821) );
  XNOR2_X1 U923 ( .A(n822), .B(n821), .ZN(n823) );
  XOR2_X1 U924 ( .A(n824), .B(n823), .Z(n826) );
  XNOR2_X1 U925 ( .A(G2078), .B(G2084), .ZN(n825) );
  XNOR2_X1 U926 ( .A(n826), .B(n825), .ZN(G227) );
  XOR2_X1 U927 ( .A(G1976), .B(G1971), .Z(n828) );
  XNOR2_X1 U928 ( .A(G1986), .B(G1966), .ZN(n827) );
  XNOR2_X1 U929 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U930 ( .A(G1981), .B(G1956), .Z(n830) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n829) );
  XNOR2_X1 U932 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U933 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U934 ( .A(G2474), .B(KEYINPUT41), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U936 ( .A(KEYINPUT107), .B(n835), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n836), .B(n923), .ZN(G229) );
  NAND2_X1 U938 ( .A1(G124), .A2(n869), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n837), .B(KEYINPUT108), .ZN(n838) );
  XNOR2_X1 U940 ( .A(KEYINPUT44), .B(n838), .ZN(n841) );
  NAND2_X1 U941 ( .A1(G100), .A2(n865), .ZN(n839) );
  XOR2_X1 U942 ( .A(KEYINPUT109), .B(n839), .Z(n840) );
  NAND2_X1 U943 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U944 ( .A1(G112), .A2(n870), .ZN(n843) );
  NAND2_X1 U945 ( .A1(G136), .A2(n866), .ZN(n842) );
  NAND2_X1 U946 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U947 ( .A1(n845), .A2(n844), .ZN(G162) );
  NAND2_X1 U948 ( .A1(G130), .A2(n869), .ZN(n847) );
  NAND2_X1 U949 ( .A1(G118), .A2(n870), .ZN(n846) );
  NAND2_X1 U950 ( .A1(n847), .A2(n846), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G106), .A2(n865), .ZN(n849) );
  NAND2_X1 U952 ( .A1(G142), .A2(n866), .ZN(n848) );
  NAND2_X1 U953 ( .A1(n849), .A2(n848), .ZN(n850) );
  XOR2_X1 U954 ( .A(n850), .B(KEYINPUT45), .Z(n851) );
  NOR2_X1 U955 ( .A1(n852), .A2(n851), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n861) );
  XNOR2_X1 U957 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT46), .ZN(n856) );
  XOR2_X1 U959 ( .A(n856), .B(G160), .Z(n859) );
  XOR2_X1 U960 ( .A(n857), .B(G164), .Z(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U962 ( .A(n861), .B(n860), .Z(n864) );
  XOR2_X1 U963 ( .A(n862), .B(G162), .Z(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n877) );
  NAND2_X1 U965 ( .A1(G103), .A2(n865), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G139), .A2(n866), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n875) );
  NAND2_X1 U968 ( .A1(G127), .A2(n869), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G115), .A2(n870), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n873), .Z(n874) );
  NOR2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n1001) );
  XNOR2_X1 U973 ( .A(n1001), .B(n986), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n878) );
  NOR2_X1 U975 ( .A1(G37), .A2(n878), .ZN(G395) );
  XNOR2_X1 U976 ( .A(n960), .B(G286), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n881), .B(G171), .ZN(n882) );
  NOR2_X1 U979 ( .A1(G37), .A2(n882), .ZN(G397) );
  XOR2_X1 U980 ( .A(KEYINPUT103), .B(G2446), .Z(n884) );
  XNOR2_X1 U981 ( .A(KEYINPUT101), .B(G2451), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U983 ( .A(n885), .B(G2430), .Z(n887) );
  XNOR2_X1 U984 ( .A(G1341), .B(G1348), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n891) );
  XOR2_X1 U986 ( .A(G2438), .B(G2435), .Z(n889) );
  XNOR2_X1 U987 ( .A(KEYINPUT102), .B(G2454), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U989 ( .A(n891), .B(n890), .Z(n893) );
  XNOR2_X1 U990 ( .A(G2443), .B(G2427), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n894) );
  NAND2_X1 U992 ( .A1(n894), .A2(G14), .ZN(n901) );
  NAND2_X1 U993 ( .A1(G319), .A2(n901), .ZN(n898) );
  NOR2_X1 U994 ( .A1(G227), .A2(G229), .ZN(n895) );
  XOR2_X1 U995 ( .A(KEYINPUT49), .B(n895), .Z(n896) );
  XNOR2_X1 U996 ( .A(n896), .B(KEYINPUT111), .ZN(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n900) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n899) );
  NAND2_X1 U999 ( .A1(n900), .A2(n899), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(G69), .ZN(G235) );
  INV_X1 U1002 ( .A(n901), .ZN(G401) );
  XNOR2_X1 U1003 ( .A(KEYINPUT54), .B(G34), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n902), .B(KEYINPUT115), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(G2084), .B(n903), .ZN(n919) );
  XNOR2_X1 U1006 ( .A(G2090), .B(G35), .ZN(n917) );
  XOR2_X1 U1007 ( .A(G2072), .B(G33), .Z(n904) );
  NAND2_X1 U1008 ( .A1(n904), .A2(G28), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(G2067), .B(G26), .ZN(n906) );
  XNOR2_X1 U1010 ( .A(G1996), .B(G32), .ZN(n905) );
  NOR2_X1 U1011 ( .A1(n906), .A2(n905), .ZN(n912) );
  XOR2_X1 U1012 ( .A(n907), .B(G27), .Z(n910) );
  XNOR2_X1 U1013 ( .A(n908), .B(G25), .ZN(n909) );
  NOR2_X1 U1014 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1015 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(KEYINPUT53), .B(n915), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n920), .B(KEYINPUT116), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n921), .B(KEYINPUT55), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(G29), .A2(n922), .ZN(n983) );
  XNOR2_X1 U1023 ( .A(G5), .B(n923), .ZN(n943) );
  XOR2_X1 U1024 ( .A(G1981), .B(G6), .Z(n926) );
  XNOR2_X1 U1025 ( .A(G1956), .B(G20), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(n924), .B(KEYINPUT123), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(G19), .B(G1341), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT124), .B(n929), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(G1348), .B(KEYINPUT59), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(n930), .B(G4), .ZN(n931) );
  NAND2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(n933), .B(KEYINPUT60), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(G1986), .B(G24), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(G23), .B(G1976), .ZN(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(G1971), .B(KEYINPUT125), .ZN(n936) );
  XNOR2_X1 U1039 ( .A(n936), .B(G22), .ZN(n937) );
  NAND2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1041 ( .A(KEYINPUT58), .B(n939), .ZN(n940) );
  NOR2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(G21), .B(G1966), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1046 ( .A(KEYINPUT61), .B(n946), .Z(n947) );
  NOR2_X1 U1047 ( .A1(G16), .A2(n947), .ZN(n979) );
  XOR2_X1 U1048 ( .A(G16), .B(KEYINPUT56), .Z(n977) );
  XNOR2_X1 U1049 ( .A(KEYINPUT119), .B(n948), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(G166), .B(G1971), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(n951), .B(G1956), .ZN(n952) );
  NAND2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1055 ( .A(KEYINPUT120), .B(n956), .Z(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1057 ( .A(KEYINPUT121), .B(n959), .Z(n971) );
  XNOR2_X1 U1058 ( .A(n960), .B(G1348), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(G171), .B(G1961), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G168), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(n965), .B(KEYINPUT57), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n966) );
  XNOR2_X1 U1065 ( .A(n967), .B(n966), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G1341), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(n975), .B(KEYINPUT122), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(KEYINPUT126), .B(n980), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(G11), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(n984), .B(KEYINPUT127), .ZN(n1014) );
  INV_X1 U1077 ( .A(G29), .ZN(n1012) );
  XOR2_X1 U1078 ( .A(G2084), .B(G160), .Z(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(KEYINPUT112), .B(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(KEYINPUT113), .ZN(n1000) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n995) );
  XNOR2_X1 U1086 ( .A(KEYINPUT114), .B(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1088 ( .A(KEYINPUT51), .B(n998), .Z(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1008) );
  XOR2_X1 U1090 ( .A(G2072), .B(n1001), .Z(n1003) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(n1004), .B(KEYINPUT50), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1009), .Z(n1010) );
  NOR2_X1 U1097 ( .A1(KEYINPUT55), .A2(n1010), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(KEYINPUT62), .B(n1015), .ZN(G311) );
  INV_X1 U1101 ( .A(G311), .ZN(G150) );
endmodule

