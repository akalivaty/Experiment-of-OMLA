//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907;
  INV_X1    g000(.A(G64gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G57gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT95), .B(G57gat), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n205), .B2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n207), .B(new_n209), .C1(new_n213), .C2(new_n210), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT7), .ZN(new_n217));
  INV_X1    g016(.A(G99gat), .ZN(new_n218));
  INV_X1    g017(.A(G106gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT8), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n220), .C1(G85gat), .C2(G92gat), .ZN(new_n221));
  XOR2_X1   g020(.A(G99gat), .B(G106gat), .Z(new_n222));
  OAI21_X1  g021(.A(KEYINPUT99), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n221), .B(new_n222), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n215), .A2(KEYINPUT10), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n226), .A2(KEYINPUT10), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G230gat), .A2(G233gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n229), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT100), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n231), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G120gat), .B(G148gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(G176gat), .B(G204gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT102), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n237), .A2(new_n241), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT101), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G43gat), .B(G50gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT15), .ZN(new_n249));
  NAND2_X1  g048(.A1(G29gat), .A2(G36gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(G29gat), .A2(G36gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT14), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n249), .A2(new_n250), .A3(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n248), .A2(KEYINPUT15), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT90), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n254), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT90), .B1(new_n251), .B2(new_n252), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n250), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n249), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n256), .A2(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT17), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT93), .ZN(new_n265));
  XNOR2_X1  g064(.A(G15gat), .B(G22gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT16), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n266), .B1(new_n267), .B2(G1gat), .ZN(new_n268));
  INV_X1    g067(.A(G8gat), .ZN(new_n269));
  OAI221_X1 g068(.A(new_n268), .B1(KEYINPUT91), .B2(new_n269), .C1(G1gat), .C2(new_n266), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n269), .A2(KEYINPUT91), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT92), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n263), .A2(KEYINPUT17), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n272), .A2(KEYINPUT92), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n265), .A2(new_n273), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G229gat), .A2(G233gat), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n272), .A2(new_n263), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT18), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT94), .ZN(new_n282));
  XNOR2_X1  g081(.A(G113gat), .B(G141gat), .ZN(new_n283));
  INV_X1    g082(.A(G197gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(KEYINPUT11), .B(G169gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n287), .B(KEYINPUT12), .Z(new_n288));
  XNOR2_X1  g087(.A(new_n272), .B(new_n263), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n277), .B(KEYINPUT13), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n279), .A2(new_n280), .ZN(new_n292));
  AND4_X1   g091(.A1(new_n282), .A2(new_n288), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n281), .A2(KEYINPUT94), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n288), .B(KEYINPUT89), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n291), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n296), .B1(new_n297), .B2(new_n281), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n247), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT27), .B(G183gat), .ZN(new_n302));
  INV_X1    g101(.A(G190gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(KEYINPUT28), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n305));
  AND2_X1   g104(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT27), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(KEYINPUT27), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n310), .ZN(new_n319));
  AOI21_X1  g118(.A(G190gat), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n320), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n304), .B1(new_n313), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n322), .A2(new_n323), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT71), .B(G120gat), .ZN(new_n332));
  MUX2_X1   g131(.A(G120gat), .B(new_n332), .S(G113gat), .Z(new_n333));
  XOR2_X1   g132(.A(G127gat), .B(G134gat), .Z(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(KEYINPUT1), .ZN(new_n335));
  XNOR2_X1  g134(.A(G113gat), .B(G120gat), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n336), .A2(KEYINPUT1), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n333), .A2(new_n335), .B1(new_n337), .B2(new_n334), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n315), .A2(new_n303), .ZN(new_n341));
  NAND3_X1  g140(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n343), .A2(KEYINPUT65), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n327), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n343), .A2(KEYINPUT65), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n351), .A2(KEYINPUT66), .A3(new_n327), .A4(new_n346), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n344), .A2(new_n349), .A3(new_n350), .A4(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n347), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT68), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n340), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n316), .A2(new_n317), .ZN(new_n360));
  INV_X1    g159(.A(new_n323), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n360), .A2(new_n303), .B1(KEYINPUT24), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n357), .A2(KEYINPUT25), .A3(new_n363), .A4(new_n351), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n331), .A2(new_n338), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT72), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n331), .A2(new_n365), .ZN(new_n368));
  INV_X1    g167(.A(new_n338), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n331), .A2(new_n371), .A3(new_n338), .A4(new_n365), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G15gat), .B(G43gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G71gat), .B(G99gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n373), .A2(new_n375), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n376), .A2(KEYINPUT32), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT34), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n376), .A2(KEYINPUT32), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n376), .B2(KEYINPUT32), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT32), .ZN(new_n391));
  AOI211_X1 g190(.A(new_n391), .B(KEYINPUT34), .C1(new_n373), .C2(new_n375), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n390), .A2(new_n392), .A3(new_n383), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n382), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT31), .B(G50gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT73), .B(G204gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(new_n284), .ZN(new_n398));
  AND2_X1   g197(.A1(G211gat), .A2(G218gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(KEYINPUT22), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G211gat), .B(G218gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT74), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n400), .B(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n396), .B1(new_n403), .B2(KEYINPUT29), .ZN(new_n404));
  NAND2_X1  g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT2), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT78), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G148gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G141gat), .ZN(new_n410));
  INV_X1    g209(.A(G141gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(G148gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n405), .A2(KEYINPUT78), .A3(KEYINPUT2), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n408), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(G155gat), .A2(G162gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n405), .A2(KEYINPUT77), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT77), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(G155gat), .A3(G162gat), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G155gat), .B(G162gat), .ZN(new_n422));
  AND2_X1   g221(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n424));
  INV_X1    g223(.A(G155gat), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT2), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n413), .B(new_n422), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n404), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G78gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n421), .A2(new_n428), .A3(new_n396), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n421), .A2(new_n428), .A3(KEYINPUT81), .A4(new_n396), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n403), .B1(new_n437), .B2(KEYINPUT29), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n431), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n431), .B1(new_n430), .B2(new_n438), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n395), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n443), .B(G22gat), .Z(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(G106gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n438), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(G78gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n395), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n439), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n442), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n445), .B1(new_n442), .B2(new_n449), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n386), .A2(new_n388), .A3(new_n384), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n383), .B1(new_n390), .B2(new_n392), .ZN(new_n454));
  INV_X1    g253(.A(new_n382), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n394), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(G226gat), .ZN(new_n458));
  INV_X1    g257(.A(G233gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT75), .ZN(new_n462));
  INV_X1    g261(.A(new_n304), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT70), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n306), .A2(new_n307), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n310), .B1(new_n465), .B2(KEYINPUT27), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n305), .B(new_n312), .C1(new_n466), .C2(G190gat), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n468), .A2(new_n361), .A3(new_n329), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n355), .A2(new_n364), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n331), .A2(KEYINPUT75), .A3(new_n365), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n460), .A2(KEYINPUT29), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n368), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n403), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n331), .A2(new_n460), .A3(new_n365), .ZN(new_n479));
  INV_X1    g278(.A(new_n403), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G8gat), .B(G36gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(G64gat), .B(G92gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(KEYINPUT76), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT76), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n477), .B2(new_n481), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(KEYINPUT30), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n481), .A3(new_n485), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(KEYINPUT30), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n489), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT86), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n494), .A2(new_n493), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n492), .A4(new_n489), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n457), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n338), .B(new_n429), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n507));
  OR2_X1    g306(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(G155gat), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n510), .A2(KEYINPUT2), .B1(new_n410), .B2(new_n412), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n511), .A2(new_n422), .B1(new_n415), .B2(new_n420), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n507), .B1(new_n512), .B2(new_n396), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n429), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n513), .A2(new_n514), .B1(new_n434), .B2(new_n435), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT4), .B1(new_n369), .B2(new_n429), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n338), .A2(new_n517), .A3(new_n512), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n515), .A2(new_n369), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n506), .B1(new_n519), .B2(new_n503), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n513), .A2(new_n514), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(new_n369), .A3(new_n436), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n518), .ZN(new_n523));
  AND4_X1   g322(.A1(new_n503), .A2(new_n522), .A3(new_n523), .A4(new_n506), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n505), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G1gat), .B(G29gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G85gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT0), .B(G57gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n527), .B(new_n528), .Z(new_n529));
  NOR2_X1   g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT85), .B1(new_n530), .B2(KEYINPUT6), .ZN(new_n531));
  INV_X1    g330(.A(new_n506), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n522), .A2(new_n523), .ZN(new_n533));
  INV_X1    g332(.A(new_n503), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n503), .A3(new_n506), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n504), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n529), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT85), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT6), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n531), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT83), .B1(new_n537), .B2(new_n538), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT83), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n525), .A2(new_n545), .A3(new_n529), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n544), .A2(new_n546), .A3(new_n541), .A4(new_n539), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT35), .B1(new_n500), .B2(new_n548), .ZN(new_n549));
  AND4_X1   g348(.A1(KEYINPUT35), .A2(new_n394), .A3(new_n452), .A4(new_n456), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n546), .A3(new_n541), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT84), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n544), .A2(new_n546), .A3(KEYINPUT84), .A4(new_n541), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n539), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n495), .B1(new_n555), .B2(new_n543), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n549), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n543), .ZN(new_n560));
  INV_X1    g359(.A(new_n495), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n452), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n564));
  INV_X1    g363(.A(new_n456), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n455), .B1(new_n453), .B2(new_n454), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n394), .A2(KEYINPUT36), .A3(new_n456), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n562), .A2(new_n563), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n482), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT37), .B1(new_n477), .B2(new_n481), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT38), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n543), .A2(new_n547), .A3(new_n573), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n482), .A2(KEYINPUT38), .A3(new_n485), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n478), .A2(new_n479), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n403), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n469), .A2(new_n470), .A3(new_n462), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT75), .B1(new_n331), .B2(new_n365), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n460), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n475), .A3(new_n480), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(KEYINPUT37), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT88), .ZN(new_n583));
  INV_X1    g382(.A(new_n572), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT88), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n577), .A2(new_n581), .A3(new_n586), .A4(KEYINPUT37), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n575), .B1(new_n588), .B2(new_n485), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n574), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n533), .A2(new_n534), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT87), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT39), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n591), .B(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n593), .B1(new_n501), .B2(new_n503), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n594), .A2(new_n598), .A3(new_n529), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n599), .A2(KEYINPUT40), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n530), .B1(new_n599), .B2(KEYINPUT40), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n496), .A2(new_n499), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n590), .A2(new_n602), .A3(new_n452), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n569), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n559), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n215), .A2(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n272), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G183gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n215), .A2(KEYINPUT21), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G211gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  NAND3_X1  g416(.A1(new_n265), .A2(new_n225), .A3(new_n274), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n225), .A2(new_n263), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G190gat), .B(G218gat), .Z(new_n622));
  OAI211_X1 g421(.A(new_n618), .B(new_n621), .C1(KEYINPUT97), .C2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n623), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(KEYINPUT97), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT96), .B(KEYINPUT98), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n627), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AND4_X1   g431(.A1(new_n301), .A2(new_n605), .A3(new_n617), .A4(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n560), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g435(.A1(new_n496), .A2(new_n499), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n267), .A2(new_n269), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT42), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n639), .A2(new_n269), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT103), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(G1325gat));
  NOR2_X1   g445(.A1(new_n565), .A2(new_n566), .ZN(new_n647));
  AOI21_X1  g446(.A(G15gat), .B1(new_n633), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n567), .A2(new_n568), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n650), .A2(G15gat), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n648), .B1(new_n633), .B2(new_n651), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n563), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT43), .B(G22gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  XNOR2_X1  g454(.A(new_n615), .B(new_n616), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n301), .ZN(new_n657));
  AOI211_X1 g456(.A(new_n632), .B(new_n657), .C1(new_n559), .C2(new_n604), .ZN(new_n658));
  INV_X1    g457(.A(G29gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n634), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT104), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT45), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n549), .B2(new_n558), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n394), .A2(new_n452), .A3(new_n456), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n637), .A3(new_n548), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT35), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(KEYINPUT106), .A3(new_n557), .ZN(new_n670));
  AND4_X1   g469(.A1(new_n496), .A2(new_n499), .A3(new_n600), .A4(new_n601), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n452), .B1(new_n574), .B2(new_n589), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n568), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT36), .B1(new_n394), .B2(new_n456), .ZN(new_n675));
  OAI22_X1  g474(.A1(new_n674), .A2(new_n675), .B1(new_n556), .B2(new_n452), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT105), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n569), .A2(new_n603), .A3(new_n678), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n665), .A2(new_n670), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n663), .B1(new_n680), .B2(new_n632), .ZN(new_n681));
  INV_X1    g480(.A(new_n657), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n605), .A2(KEYINPUT44), .A3(new_n631), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685), .B2(new_n560), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n662), .A2(new_n686), .ZN(G1328gat));
  OAI21_X1  g486(.A(G36gat), .B1(new_n685), .B2(new_n637), .ZN(new_n688));
  INV_X1    g487(.A(G36gat), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n658), .A2(new_n689), .A3(new_n638), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT46), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(G1329gat));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n693), .A2(KEYINPUT108), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(KEYINPUT108), .ZN(new_n695));
  OAI21_X1  g494(.A(G43gat), .B1(new_n685), .B2(new_n649), .ZN(new_n696));
  INV_X1    g495(.A(G43gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n658), .A2(new_n697), .A3(new_n647), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT107), .ZN(new_n699));
  AOI211_X1 g498(.A(new_n694), .B(new_n695), .C1(new_n696), .C2(new_n699), .ZN(new_n700));
  AND4_X1   g499(.A1(KEYINPUT108), .A2(new_n696), .A3(new_n693), .A4(new_n699), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(G1330gat));
  NAND3_X1  g501(.A1(new_n684), .A2(G50gat), .A3(new_n563), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n658), .A2(new_n563), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(G50gat), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g505(.A1(new_n243), .A2(new_n246), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n617), .A2(new_n300), .A3(new_n632), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n680), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n634), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n205), .ZN(G1332gat));
  AOI21_X1  g510(.A(new_n637), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT109), .Z(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT110), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1333gat));
  INV_X1    g516(.A(G71gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n709), .A2(new_n718), .A3(new_n647), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n709), .A2(new_n650), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(new_n718), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g521(.A1(new_n709), .A2(new_n563), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G78gat), .ZN(G1335gat));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n680), .B2(new_n632), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n617), .A2(new_n299), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT106), .B1(new_n669), .B2(new_n557), .ZN(new_n728));
  AOI221_X4 g527(.A(new_n664), .B1(new_n550), .B2(new_n556), .C1(new_n667), .C2(new_n668), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n673), .A2(new_n676), .A3(KEYINPUT105), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n678), .B1(new_n569), .B2(new_n603), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n728), .A2(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(KEYINPUT111), .A3(new_n631), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n726), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n726), .A2(new_n733), .A3(KEYINPUT51), .A4(new_n727), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n560), .A2(G85gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n247), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n681), .A2(new_n247), .A3(new_n683), .A4(new_n727), .ZN(new_n741));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n560), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT112), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n740), .A2(new_n745), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(G1336gat));
  NOR2_X1   g546(.A1(new_n637), .A2(G92gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n738), .A2(new_n247), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G92gat), .B1(new_n741), .B2(new_n637), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(KEYINPUT52), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  INV_X1    g552(.A(new_n748), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n707), .B(new_n754), .C1(new_n736), .C2(new_n737), .ZN(new_n755));
  INV_X1    g554(.A(new_n750), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n752), .A2(new_n757), .ZN(G1337gat));
  NAND3_X1  g557(.A1(new_n247), .A2(new_n218), .A3(new_n647), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT115), .Z(new_n760));
  NAND2_X1  g559(.A1(new_n738), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n741), .A2(new_n649), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT114), .Z(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(new_n218), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n247), .A2(new_n219), .A3(new_n563), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT116), .Z(new_n766));
  NAND2_X1  g565(.A1(new_n738), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G106gat), .B1(new_n741), .B2(new_n452), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n767), .B(new_n768), .C1(new_n771), .C2(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1339gat));
  NOR2_X1   g574(.A1(new_n708), .A2(new_n247), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n289), .A2(new_n290), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT118), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n276), .A2(new_n278), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(G229gat), .A3(G233gat), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n287), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n293), .B2(new_n294), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n247), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n240), .B1(new_n230), .B2(KEYINPUT54), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n228), .A2(new_n229), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(KEYINPUT54), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n785), .B1(new_n787), .B2(new_n230), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n788), .A2(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(KEYINPUT55), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n246), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n300), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n632), .B1(new_n784), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n782), .A2(new_n631), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT119), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n791), .A2(KEYINPUT119), .A3(new_n794), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n776), .B1(new_n798), .B2(new_n656), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n799), .A2(new_n638), .A3(new_n457), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n634), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n801), .A2(new_n300), .B1(KEYINPUT120), .B2(G113gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(KEYINPUT120), .A2(G113gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT121), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n802), .B(new_n804), .ZN(G1340gat));
  INV_X1    g604(.A(new_n801), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n332), .A3(new_n247), .ZN(new_n807));
  OAI21_X1  g606(.A(G120gat), .B1(new_n801), .B2(new_n707), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT122), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n811), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1341gat));
  NAND2_X1  g612(.A1(new_n806), .A2(new_n617), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g614(.A1(new_n806), .A2(new_n631), .ZN(new_n816));
  OR3_X1    g615(.A1(new_n816), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(G134gat), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT56), .B1(new_n816), .B2(G134gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(G1343gat));
  OAI21_X1  g619(.A(KEYINPUT57), .B1(new_n799), .B2(new_n452), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n796), .A2(new_n797), .ZN(new_n822));
  INV_X1    g621(.A(new_n792), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n631), .B1(new_n823), .B2(new_n783), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n656), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n776), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n563), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n650), .A2(new_n560), .A3(new_n638), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n821), .A2(new_n829), .A3(new_n299), .A4(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(G141gat), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n827), .A2(new_n563), .A3(new_n830), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n833), .A2(new_n411), .A3(new_n299), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT58), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n821), .A2(new_n829), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n836), .A2(new_n837), .A3(new_n299), .A4(new_n830), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(KEYINPUT123), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n838), .A2(G141gat), .A3(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n834), .A2(KEYINPUT58), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n835), .B1(new_n840), .B2(new_n841), .ZN(G1344gat));
  NAND3_X1  g641(.A1(new_n833), .A2(new_n409), .A3(new_n247), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n836), .A2(new_n247), .A3(new_n830), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n844), .A2(new_n845), .A3(G148gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n617), .B1(new_n793), .B2(new_n795), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n828), .B(new_n563), .C1(new_n847), .C2(new_n776), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n821), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n830), .B(KEYINPUT124), .Z(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n247), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n845), .B1(new_n851), .B2(G148gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n843), .B1(new_n846), .B2(new_n852), .ZN(G1345gat));
  AOI21_X1  g652(.A(G155gat), .B1(new_n833), .B2(new_n617), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n836), .A2(new_n830), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n656), .A2(new_n425), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(G1346gat));
  NAND2_X1  g656(.A1(new_n508), .A2(new_n509), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n632), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n833), .A2(new_n631), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n855), .A2(new_n859), .B1(new_n858), .B2(new_n860), .ZN(G1347gat));
  NAND4_X1  g660(.A1(new_n827), .A2(new_n560), .A3(new_n638), .A4(new_n666), .ZN(new_n862));
  OAI21_X1  g661(.A(G169gat), .B1(new_n862), .B2(new_n300), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n862), .A2(KEYINPUT125), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(KEYINPUT125), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n300), .A2(G169gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(G1348gat));
  INV_X1    g667(.A(G176gat), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n862), .A2(new_n869), .A3(new_n707), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n864), .A2(new_n247), .A3(new_n865), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n869), .ZN(G1349gat));
  INV_X1    g671(.A(new_n862), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n302), .A3(new_n617), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n465), .B1(new_n862), .B2(new_n656), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(new_n631), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(G190gat), .ZN(new_n880));
  AOI211_X1 g679(.A(KEYINPUT61), .B(new_n303), .C1(new_n873), .C2(new_n631), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n631), .A2(new_n303), .ZN(new_n882));
  OAI22_X1  g681(.A1(new_n880), .A2(new_n881), .B1(new_n866), .B2(new_n882), .ZN(G1351gat));
  NAND3_X1  g682(.A1(new_n827), .A2(new_n560), .A3(new_n638), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n452), .A3(new_n650), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n284), .A3(new_n299), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n650), .A2(new_n634), .A3(new_n637), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n849), .A2(new_n299), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n886), .B1(new_n888), .B2(new_n284), .ZN(G1352gat));
  XOR2_X1   g688(.A(KEYINPUT126), .B(G204gat), .Z(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n885), .A2(new_n247), .A3(new_n891), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT62), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(KEYINPUT62), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n849), .A2(new_n247), .A3(new_n887), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n893), .B(new_n894), .C1(new_n891), .C2(new_n895), .ZN(G1353gat));
  INV_X1    g695(.A(G211gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n885), .A2(new_n897), .A3(new_n617), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n849), .A2(new_n617), .A3(new_n887), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n899), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT63), .B1(new_n899), .B2(G211gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(G1354gat));
  INV_X1    g701(.A(G218gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n903), .A3(new_n631), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n821), .A2(new_n631), .A3(new_n848), .A4(new_n887), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G218gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


