

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738;

  XNOR2_X1 U366 ( .A(G110), .B(G104), .ZN(n455) );
  XNOR2_X1 U367 ( .A(n455), .B(G107), .ZN(n507) );
  AND2_X1 U368 ( .A1(n422), .A2(n593), .ZN(n529) );
  XNOR2_X1 U369 ( .A(n436), .B(n433), .ZN(n714) );
  NOR2_X1 U370 ( .A1(n669), .A2(n361), .ZN(n526) );
  INV_X2 U371 ( .A(G953), .ZN(n725) );
  AND2_X4 U372 ( .A1(n345), .A2(n344), .ZN(n390) );
  XNOR2_X2 U373 ( .A(n346), .B(KEYINPUT64), .ZN(n345) );
  INV_X2 U374 ( .A(G128), .ZN(n397) );
  NAND2_X2 U375 ( .A1(n370), .A2(n368), .ZN(n568) );
  NAND2_X2 U376 ( .A1(n437), .A2(n621), .ZN(n544) );
  XNOR2_X1 U377 ( .A(n508), .B(n509), .ZN(n692) );
  INV_X1 U378 ( .A(n683), .ZN(n344) );
  NOR2_X1 U379 ( .A1(n680), .A2(n679), .ZN(n683) );
  NAND2_X1 U380 ( .A1(n563), .A2(n565), .ZN(n642) );
  NOR2_X1 U381 ( .A1(G902), .A2(n608), .ZN(n502) );
  XNOR2_X1 U382 ( .A(n401), .B(G131), .ZN(n494) );
  INV_X1 U383 ( .A(KEYINPUT16), .ZN(n435) );
  XNOR2_X1 U384 ( .A(G119), .B(G116), .ZN(n452) );
  INV_X1 U385 ( .A(KEYINPUT3), .ZN(n451) );
  NAND2_X1 U386 ( .A1(n392), .A2(n394), .ZN(n347) );
  AND2_X1 U387 ( .A1(n587), .A2(n408), .ZN(n592) );
  NOR2_X1 U388 ( .A1(n737), .A2(n539), .ZN(n540) );
  XNOR2_X1 U389 ( .A(n522), .B(KEYINPUT101), .ZN(n737) );
  XNOR2_X1 U390 ( .A(n421), .B(n528), .ZN(n734) );
  NOR2_X1 U391 ( .A1(n384), .A2(n387), .ZN(n636) );
  XNOR2_X1 U392 ( .A(n375), .B(KEYINPUT39), .ZN(n560) );
  XNOR2_X1 U393 ( .A(n426), .B(KEYINPUT75), .ZN(n628) );
  XNOR2_X1 U394 ( .A(n445), .B(n444), .ZN(n575) );
  XNOR2_X1 U395 ( .A(n374), .B(n351), .ZN(n563) );
  XNOR2_X1 U396 ( .A(n484), .B(n415), .ZN(n534) );
  NOR2_X2 U397 ( .A1(n462), .A2(n603), .ZN(n465) );
  XNOR2_X1 U398 ( .A(n507), .B(n434), .ZN(n433) );
  XNOR2_X1 U399 ( .A(n454), .B(n453), .ZN(n436) );
  XNOR2_X1 U400 ( .A(n490), .B(G134), .ZN(n496) );
  XNOR2_X1 U401 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U402 ( .A(n435), .B(G122), .ZN(n434) );
  XNOR2_X1 U403 ( .A(n404), .B(G146), .ZN(n364) );
  XNOR2_X1 U404 ( .A(n452), .B(n451), .ZN(n454) );
  INV_X1 U405 ( .A(KEYINPUT66), .ZN(n401) );
  INV_X1 U406 ( .A(G125), .ZN(n404) );
  NAND2_X1 U407 ( .A1(n708), .A2(n724), .ZN(n680) );
  XNOR2_X2 U408 ( .A(n396), .B(KEYINPUT45), .ZN(n708) );
  NAND2_X1 U409 ( .A1(n347), .A2(n391), .ZN(n346) );
  BUF_X1 U410 ( .A(n708), .Z(n348) );
  NAND2_X2 U411 ( .A1(n557), .A2(n659), .ZN(n591) );
  XNOR2_X2 U412 ( .A(n465), .B(n464), .ZN(n557) );
  XNOR2_X2 U413 ( .A(n591), .B(KEYINPUT19), .ZN(n583) );
  AND2_X1 U414 ( .A1(n724), .A2(n446), .ZN(n393) );
  AND2_X1 U415 ( .A1(n372), .A2(n371), .ZN(n370) );
  NAND2_X1 U416 ( .A1(n510), .A2(n381), .ZN(n369) );
  XNOR2_X1 U417 ( .A(n568), .B(KEYINPUT1), .ZN(n593) );
  XNOR2_X1 U418 ( .A(n418), .B(n416), .ZN(n695) );
  XNOR2_X1 U419 ( .A(n481), .B(n417), .ZN(n416) );
  NOR2_X1 U420 ( .A1(G902), .A2(G237), .ZN(n463) );
  NOR2_X1 U421 ( .A1(G953), .A2(G237), .ZN(n501) );
  INV_X1 U422 ( .A(KEYINPUT71), .ZN(n498) );
  XOR2_X1 U423 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n499) );
  XNOR2_X1 U424 ( .A(G902), .B(KEYINPUT15), .ZN(n602) );
  XNOR2_X1 U425 ( .A(n413), .B(n412), .ZN(n533) );
  INV_X1 U426 ( .A(G478), .ZN(n412) );
  NAND2_X1 U427 ( .A1(n382), .A2(n381), .ZN(n413) );
  AND2_X1 U428 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U429 ( .A(n410), .B(n409), .ZN(n516) );
  INV_X1 U430 ( .A(KEYINPUT8), .ZN(n409) );
  NAND2_X1 U431 ( .A1(n725), .A2(G234), .ZN(n410) );
  XNOR2_X1 U432 ( .A(KEYINPUT10), .B(G140), .ZN(n427) );
  XNOR2_X1 U433 ( .A(KEYINPUT73), .B(KEYINPUT91), .ZN(n511) );
  XOR2_X1 U434 ( .A(KEYINPUT92), .B(KEYINPUT24), .Z(n512) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n423) );
  XNOR2_X1 U436 ( .A(G110), .B(G119), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n514), .B(n450), .ZN(n378) );
  XNOR2_X1 U438 ( .A(G128), .B(G137), .ZN(n514) );
  XNOR2_X1 U439 ( .A(G116), .B(G122), .ZN(n485) );
  XNOR2_X1 U440 ( .A(n380), .B(G107), .ZN(n486) );
  INV_X1 U441 ( .A(KEYINPUT7), .ZN(n380) );
  NAND2_X1 U442 ( .A1(n446), .A2(n395), .ZN(n394) );
  INV_X1 U443 ( .A(KEYINPUT79), .ZN(n395) );
  XOR2_X1 U444 ( .A(G140), .B(KEYINPUT89), .Z(n505) );
  AND2_X1 U445 ( .A1(n575), .A2(n660), .ZN(n376) );
  NAND2_X1 U446 ( .A1(n400), .A2(KEYINPUT36), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n403), .B(KEYINPUT102), .ZN(n594) );
  NOR2_X1 U448 ( .A1(n705), .A2(G902), .ZN(n374) );
  AND2_X1 U449 ( .A1(n569), .A2(n568), .ZN(n582) );
  INV_X1 U450 ( .A(G475), .ZN(n415) );
  NAND2_X1 U451 ( .A1(n373), .A2(G902), .ZN(n371) );
  XNOR2_X1 U452 ( .A(KEYINPUT90), .B(KEYINPUT23), .ZN(n450) );
  XOR2_X1 U453 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n480) );
  XNOR2_X1 U454 ( .A(n476), .B(n477), .ZN(n419) );
  XNOR2_X1 U455 ( .A(G113), .B(G143), .ZN(n476) );
  XNOR2_X1 U456 ( .A(G122), .B(G104), .ZN(n477) );
  XNOR2_X1 U457 ( .A(n494), .B(n478), .ZN(n417) );
  XOR2_X1 U458 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n478) );
  AND2_X1 U459 ( .A1(n604), .A2(n447), .ZN(n446) );
  NAND2_X1 U460 ( .A1(n602), .A2(KEYINPUT79), .ZN(n447) );
  NAND2_X1 U461 ( .A1(G237), .A2(G234), .ZN(n468) );
  XNOR2_X1 U462 ( .A(n558), .B(n599), .ZN(n660) );
  XOR2_X1 U463 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n473) );
  XNOR2_X1 U464 ( .A(n508), .B(n448), .ZN(n608) );
  XNOR2_X1 U465 ( .A(n500), .B(n354), .ZN(n449) );
  INV_X1 U466 ( .A(n639), .ZN(n438) );
  BUF_X1 U467 ( .A(n557), .Z(n599) );
  INV_X1 U468 ( .A(KEYINPUT30), .ZN(n444) );
  NAND2_X1 U469 ( .A1(n651), .A2(n659), .ZN(n445) );
  INV_X1 U470 ( .A(n662), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n399), .B(n515), .ZN(n705) );
  XNOR2_X1 U472 ( .A(n423), .B(n517), .ZN(n399) );
  XNOR2_X1 U473 ( .A(n489), .B(n383), .ZN(n702) );
  XNOR2_X1 U474 ( .A(n491), .B(n349), .ZN(n383) );
  XOR2_X1 U475 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n488) );
  XNOR2_X1 U476 ( .A(n695), .B(n694), .ZN(n696) );
  INV_X1 U477 ( .A(n707), .ZN(n366) );
  XNOR2_X1 U478 ( .A(n572), .B(KEYINPUT42), .ZN(n736) );
  XNOR2_X1 U479 ( .A(n561), .B(KEYINPUT40), .ZN(n735) );
  NAND2_X1 U480 ( .A1(n385), .A2(n353), .ZN(n384) );
  NAND2_X1 U481 ( .A1(n389), .A2(n411), .ZN(n388) );
  NAND2_X1 U482 ( .A1(n402), .A2(n352), .ZN(n522) );
  INV_X1 U483 ( .A(n521), .ZN(n402) );
  XNOR2_X1 U484 ( .A(n689), .B(n405), .ZN(G75) );
  XNOR2_X1 U485 ( .A(n406), .B(KEYINPUT118), .ZN(n405) );
  INV_X1 U486 ( .A(KEYINPUT53), .ZN(n406) );
  XOR2_X1 U487 ( .A(n486), .B(n485), .Z(n349) );
  AND2_X1 U488 ( .A1(n367), .A2(n366), .ZN(n350) );
  XNOR2_X1 U489 ( .A(KEYINPUT25), .B(n519), .ZN(n351) );
  NOR2_X1 U490 ( .A1(n407), .A2(n520), .ZN(n352) );
  AND2_X1 U491 ( .A1(n407), .A2(n386), .ZN(n353) );
  AND2_X1 U492 ( .A1(n501), .A2(G210), .ZN(n354) );
  AND2_X1 U493 ( .A1(n520), .A2(n643), .ZN(n355) );
  XOR2_X1 U494 ( .A(n636), .B(KEYINPUT82), .Z(n356) );
  AND2_X1 U495 ( .A1(n640), .A2(n438), .ZN(n357) );
  INV_X1 U496 ( .A(KEYINPUT36), .ZN(n411) );
  XOR2_X1 U497 ( .A(n461), .B(n460), .Z(n358) );
  NOR2_X1 U498 ( .A1(n602), .A2(KEYINPUT79), .ZN(n359) );
  INV_X1 U499 ( .A(n641), .ZN(n360) );
  NOR2_X1 U500 ( .A1(n643), .A2(n563), .ZN(n541) );
  BUF_X1 U501 ( .A(n531), .Z(n361) );
  XNOR2_X1 U502 ( .A(n428), .B(KEYINPUT0), .ZN(n531) );
  INV_X1 U503 ( .A(n400), .ZN(n389) );
  BUF_X1 U504 ( .A(n593), .Z(n407) );
  INV_X1 U505 ( .A(n407), .ZN(n643) );
  XNOR2_X1 U506 ( .A(n524), .B(n525), .ZN(n669) );
  NOR2_X1 U507 ( .A1(n594), .A2(n388), .ZN(n387) );
  NAND2_X1 U508 ( .A1(n594), .A2(KEYINPUT36), .ZN(n385) );
  XNOR2_X1 U509 ( .A(n722), .B(n419), .ZN(n418) );
  NAND2_X1 U510 ( .A1(n362), .A2(n541), .ZN(n542) );
  XNOR2_X1 U511 ( .A(n362), .B(KEYINPUT83), .ZN(n521) );
  AND2_X2 U512 ( .A1(n363), .A2(n588), .ZN(n362) );
  AND2_X1 U513 ( .A1(n363), .A2(n355), .ZN(n543) );
  XNOR2_X1 U514 ( .A(n442), .B(KEYINPUT22), .ZN(n363) );
  XNOR2_X1 U515 ( .A(n364), .B(n459), .ZN(n432) );
  XNOR2_X1 U516 ( .A(n364), .B(n427), .ZN(n722) );
  XNOR2_X1 U517 ( .A(n365), .B(KEYINPUT122), .ZN(G66) );
  NOR2_X2 U518 ( .A1(n706), .A2(n707), .ZN(n365) );
  XNOR2_X1 U519 ( .A(n605), .B(n358), .ZN(n367) );
  NOR2_X2 U520 ( .A1(n698), .A2(n707), .ZN(n700) );
  NOR2_X2 U521 ( .A1(n613), .A2(n707), .ZN(n615) );
  NAND2_X1 U522 ( .A1(n708), .A2(n393), .ZN(n392) );
  NAND2_X1 U523 ( .A1(n390), .A2(G217), .ZN(n704) );
  NAND2_X1 U524 ( .A1(n692), .A2(n373), .ZN(n372) );
  OR2_X1 U525 ( .A1(n692), .A2(n369), .ZN(n368) );
  INV_X1 U526 ( .A(n510), .ZN(n373) );
  NAND2_X1 U527 ( .A1(n379), .A2(n708), .ZN(n391) );
  INV_X1 U528 ( .A(n642), .ZN(n422) );
  NAND2_X1 U529 ( .A1(n560), .A2(n627), .ZN(n561) );
  NAND2_X1 U530 ( .A1(n576), .A2(n376), .ZN(n375) );
  XNOR2_X1 U531 ( .A(n556), .B(KEYINPUT72), .ZN(n576) );
  AND2_X1 U532 ( .A1(n724), .A2(n359), .ZN(n379) );
  INV_X1 U533 ( .A(G902), .ZN(n381) );
  INV_X1 U534 ( .A(n702), .ZN(n382) );
  NAND2_X1 U535 ( .A1(n390), .A2(G210), .ZN(n605) );
  NAND2_X1 U536 ( .A1(n390), .A2(G472), .ZN(n612) );
  NAND2_X1 U537 ( .A1(n390), .A2(G475), .ZN(n697) );
  NAND2_X1 U538 ( .A1(n390), .A2(G478), .ZN(n701) );
  NAND2_X1 U539 ( .A1(n390), .A2(G469), .ZN(n690) );
  NAND2_X1 U540 ( .A1(n734), .A2(KEYINPUT44), .ZN(n420) );
  NAND2_X1 U541 ( .A1(n440), .A2(n441), .ZN(n396) );
  XNOR2_X2 U542 ( .A(n397), .B(G143), .ZN(n490) );
  XNOR2_X1 U543 ( .A(n690), .B(n398), .ZN(n693) );
  XNOR2_X1 U544 ( .A(n692), .B(n691), .ZN(n398) );
  AND2_X1 U545 ( .A1(n586), .A2(n356), .ZN(n408) );
  NOR2_X1 U546 ( .A1(n589), .A2(n566), .ZN(n567) );
  NOR2_X1 U547 ( .A1(n425), .A2(n424), .ZN(n584) );
  BUF_X1 U548 ( .A(n591), .Z(n400) );
  NAND2_X1 U549 ( .A1(n590), .A2(n627), .ZN(n403) );
  XNOR2_X1 U550 ( .A(n429), .B(n714), .ZN(n462) );
  XNOR2_X1 U551 ( .A(n432), .B(n458), .ZN(n431) );
  AND2_X2 U552 ( .A1(n439), .A2(n357), .ZN(n724) );
  NAND2_X1 U553 ( .A1(n414), .A2(n565), .ZN(n443) );
  NAND2_X1 U554 ( .A1(n533), .A2(n534), .ZN(n662) );
  NAND2_X1 U555 ( .A1(n420), .A2(n538), .ZN(n539) );
  NAND2_X1 U556 ( .A1(n527), .A2(n577), .ZN(n421) );
  AND2_X1 U557 ( .A1(n628), .A2(n665), .ZN(n424) );
  XNOR2_X1 U558 ( .A(n628), .B(KEYINPUT47), .ZN(n425) );
  NAND2_X1 U559 ( .A1(n582), .A2(n583), .ZN(n426) );
  XNOR2_X2 U560 ( .A(n720), .B(n497), .ZN(n508) );
  XNOR2_X2 U561 ( .A(n496), .B(n495), .ZN(n720) );
  NAND2_X1 U562 ( .A1(n583), .A2(n471), .ZN(n428) );
  XNOR2_X1 U563 ( .A(n431), .B(n430), .ZN(n429) );
  XNOR2_X1 U564 ( .A(n490), .B(n492), .ZN(n430) );
  XNOR2_X1 U565 ( .A(n592), .B(KEYINPUT48), .ZN(n439) );
  XNOR2_X1 U566 ( .A(n449), .B(n436), .ZN(n448) );
  XNOR2_X1 U567 ( .A(n437), .B(G119), .ZN(n733) );
  XNOR2_X2 U568 ( .A(n542), .B(KEYINPUT32), .ZN(n437) );
  XNOR2_X1 U569 ( .A(n540), .B(KEYINPUT84), .ZN(n440) );
  NAND2_X1 U570 ( .A1(n549), .A2(n548), .ZN(n441) );
  NOR2_X2 U571 ( .A1(n531), .A2(n443), .ZN(n442) );
  INV_X1 U572 ( .A(n496), .ZN(n491) );
  INV_X1 U573 ( .A(n676), .ZN(n469) );
  INV_X1 U574 ( .A(n563), .ZN(n520) );
  INV_X1 U575 ( .A(KEYINPUT44), .ZN(n545) );
  XNOR2_X1 U576 ( .A(n499), .B(n498), .ZN(n500) );
  NOR2_X1 U577 ( .A1(n555), .A2(n562), .ZN(n556) );
  XNOR2_X1 U578 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U579 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U580 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U581 ( .A1(G952), .A2(n725), .ZN(n707) );
  XOR2_X1 U582 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n461) );
  XOR2_X1 U583 ( .A(KEYINPUT68), .B(G113), .Z(n453) );
  XOR2_X1 U584 ( .A(KEYINPUT74), .B(KEYINPUT17), .Z(n457) );
  XNOR2_X1 U585 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n456) );
  XNOR2_X1 U586 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U587 ( .A1(G224), .A2(n725), .ZN(n459) );
  XOR2_X1 U588 ( .A(G101), .B(KEYINPUT65), .Z(n492) );
  XNOR2_X1 U589 ( .A(n462), .B(KEYINPUT86), .ZN(n460) );
  INV_X1 U590 ( .A(n602), .ZN(n603) );
  XOR2_X1 U591 ( .A(KEYINPUT70), .B(n463), .Z(n466) );
  NAND2_X1 U592 ( .A1(G210), .A2(n466), .ZN(n464) );
  NAND2_X1 U593 ( .A1(n466), .A2(G214), .ZN(n659) );
  XNOR2_X1 U594 ( .A(G898), .B(KEYINPUT88), .ZN(n710) );
  NOR2_X1 U595 ( .A1(n725), .A2(n710), .ZN(n716) );
  NAND2_X1 U596 ( .A1(n716), .A2(G902), .ZN(n467) );
  NAND2_X1 U597 ( .A1(G952), .A2(n725), .ZN(n551) );
  NAND2_X1 U598 ( .A1(n467), .A2(n551), .ZN(n470) );
  XOR2_X1 U599 ( .A(n468), .B(KEYINPUT14), .Z(n676) );
  NAND2_X1 U600 ( .A1(G234), .A2(n602), .ZN(n472) );
  XNOR2_X1 U601 ( .A(n473), .B(n472), .ZN(n518) );
  NAND2_X1 U602 ( .A1(n518), .A2(G221), .ZN(n474) );
  XNOR2_X1 U603 ( .A(n474), .B(KEYINPUT21), .ZN(n475) );
  XOR2_X1 U604 ( .A(KEYINPUT94), .B(n475), .Z(n565) );
  INV_X1 U605 ( .A(n565), .ZN(n645) );
  NAND2_X1 U606 ( .A1(G214), .A2(n501), .ZN(n479) );
  XNOR2_X1 U607 ( .A(n480), .B(n479), .ZN(n481) );
  NOR2_X1 U608 ( .A1(G902), .A2(n695), .ZN(n483) );
  XNOR2_X1 U609 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n482) );
  XNOR2_X1 U610 ( .A(n483), .B(n482), .ZN(n484) );
  NAND2_X1 U611 ( .A1(G217), .A2(n516), .ZN(n487) );
  XNOR2_X1 U612 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U613 ( .A(G146), .B(n492), .Z(n497) );
  XNOR2_X1 U614 ( .A(G137), .B(KEYINPUT4), .ZN(n493) );
  XNOR2_X2 U615 ( .A(G472), .B(n502), .ZN(n566) );
  INV_X1 U616 ( .A(KEYINPUT6), .ZN(n503) );
  XNOR2_X1 U617 ( .A(n566), .B(n503), .ZN(n588) );
  INV_X1 U618 ( .A(n588), .ZN(n523) );
  NAND2_X1 U619 ( .A1(G227), .A2(n725), .ZN(n504) );
  XNOR2_X1 U620 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U621 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U622 ( .A(KEYINPUT67), .B(G469), .ZN(n510) );
  XNOR2_X1 U623 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U624 ( .A(n513), .B(n722), .ZN(n515) );
  NAND2_X1 U625 ( .A1(G221), .A2(n516), .ZN(n517) );
  NAND2_X1 U626 ( .A1(n518), .A2(G217), .ZN(n519) );
  XOR2_X1 U627 ( .A(KEYINPUT81), .B(KEYINPUT35), .Z(n528) );
  XNOR2_X1 U628 ( .A(KEYINPUT87), .B(KEYINPUT33), .ZN(n525) );
  NAND2_X1 U629 ( .A1(n529), .A2(n523), .ZN(n524) );
  XNOR2_X1 U630 ( .A(n526), .B(KEYINPUT34), .ZN(n527) );
  NOR2_X1 U631 ( .A1(n533), .A2(n534), .ZN(n577) );
  INV_X1 U632 ( .A(n566), .ZN(n651) );
  NAND2_X1 U633 ( .A1(n651), .A2(n529), .ZN(n653) );
  NOR2_X1 U634 ( .A1(n361), .A2(n653), .ZN(n530) );
  XNOR2_X1 U635 ( .A(n530), .B(KEYINPUT31), .ZN(n633) );
  NAND2_X1 U636 ( .A1(n422), .A2(n568), .ZN(n555) );
  NOR2_X1 U637 ( .A1(n361), .A2(n555), .ZN(n532) );
  NAND2_X1 U638 ( .A1(n532), .A2(n566), .ZN(n617) );
  NAND2_X1 U639 ( .A1(n633), .A2(n617), .ZN(n537) );
  INV_X1 U640 ( .A(n533), .ZN(n535) );
  NOR2_X1 U641 ( .A1(n535), .A2(n534), .ZN(n627) );
  NAND2_X1 U642 ( .A1(n535), .A2(n534), .ZN(n634) );
  INV_X1 U643 ( .A(n634), .ZN(n622) );
  XNOR2_X1 U644 ( .A(KEYINPUT100), .B(n622), .ZN(n559) );
  NOR2_X1 U645 ( .A1(n627), .A2(n559), .ZN(n665) );
  INV_X1 U646 ( .A(n665), .ZN(n536) );
  NAND2_X1 U647 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U648 ( .A1(n543), .A2(n566), .ZN(n621) );
  XNOR2_X2 U649 ( .A(n544), .B(KEYINPUT85), .ZN(n546) );
  XNOR2_X1 U650 ( .A(n546), .B(n545), .ZN(n549) );
  BUF_X1 U651 ( .A(n546), .Z(n547) );
  NAND2_X1 U652 ( .A1(n547), .A2(n734), .ZN(n548) );
  NOR2_X1 U653 ( .A1(G900), .A2(n725), .ZN(n550) );
  NAND2_X1 U654 ( .A1(n550), .A2(G902), .ZN(n552) );
  NAND2_X1 U655 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U656 ( .A1(n553), .A2(n469), .ZN(n554) );
  XNOR2_X1 U657 ( .A(KEYINPUT76), .B(n554), .ZN(n562) );
  XNOR2_X1 U658 ( .A(KEYINPUT38), .B(KEYINPUT69), .ZN(n558) );
  AND2_X1 U659 ( .A1(n559), .A2(n560), .ZN(n639) );
  NOR2_X1 U660 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U661 ( .A1(n565), .A2(n564), .ZN(n589) );
  XNOR2_X1 U662 ( .A(KEYINPUT28), .B(n567), .ZN(n569) );
  NAND2_X1 U663 ( .A1(n660), .A2(n659), .ZN(n664) );
  NOR2_X1 U664 ( .A1(n662), .A2(n664), .ZN(n571) );
  XNOR2_X1 U665 ( .A(KEYINPUT41), .B(KEYINPUT105), .ZN(n570) );
  XNOR2_X1 U666 ( .A(n571), .B(n570), .ZN(n657) );
  NAND2_X1 U667 ( .A1(n582), .A2(n657), .ZN(n572) );
  NAND2_X1 U668 ( .A1(n735), .A2(n736), .ZN(n574) );
  INV_X1 U669 ( .A(KEYINPUT46), .ZN(n573) );
  XNOR2_X1 U670 ( .A(n574), .B(n573), .ZN(n587) );
  NAND2_X1 U671 ( .A1(KEYINPUT47), .A2(n665), .ZN(n580) );
  AND2_X1 U672 ( .A1(n576), .A2(n575), .ZN(n579) );
  AND2_X1 U673 ( .A1(n599), .A2(n577), .ZN(n578) );
  NAND2_X1 U674 ( .A1(n579), .A2(n578), .ZN(n626) );
  NAND2_X1 U675 ( .A1(n580), .A2(n626), .ZN(n581) );
  XNOR2_X1 U676 ( .A(KEYINPUT78), .B(n581), .ZN(n585) );
  NOR2_X1 U677 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U678 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U679 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n597) );
  NOR2_X1 U680 ( .A1(n594), .A2(n407), .ZN(n595) );
  NAND2_X1 U681 ( .A1(n595), .A2(n659), .ZN(n596) );
  XNOR2_X1 U682 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U683 ( .A(n598), .B(KEYINPUT103), .ZN(n601) );
  INV_X1 U684 ( .A(n599), .ZN(n600) );
  NAND2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n640) );
  NAND2_X1 U686 ( .A1(KEYINPUT2), .A2(n603), .ZN(n604) );
  INV_X1 U687 ( .A(KEYINPUT2), .ZN(n679) );
  INV_X1 U688 ( .A(KEYINPUT119), .ZN(n606) );
  XNOR2_X1 U689 ( .A(n606), .B(KEYINPUT56), .ZN(n607) );
  XNOR2_X1 U690 ( .A(n350), .B(n607), .ZN(G51) );
  INV_X1 U691 ( .A(n608), .ZN(n610) );
  XOR2_X1 U692 ( .A(KEYINPUT62), .B(KEYINPUT106), .Z(n609) );
  XNOR2_X1 U693 ( .A(KEYINPUT63), .B(KEYINPUT107), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n615), .B(n614), .ZN(G57) );
  INV_X1 U695 ( .A(n627), .ZN(n631) );
  NOR2_X1 U696 ( .A1(n631), .A2(n617), .ZN(n616) );
  XOR2_X1 U697 ( .A(G104), .B(n616), .Z(G6) );
  NOR2_X1 U698 ( .A1(n634), .A2(n617), .ZN(n619) );
  XNOR2_X1 U699 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n618) );
  XNOR2_X1 U700 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U701 ( .A(G107), .B(n620), .ZN(G9) );
  XNOR2_X1 U702 ( .A(G110), .B(n621), .ZN(G12) );
  XOR2_X1 U703 ( .A(KEYINPUT109), .B(KEYINPUT29), .Z(n624) );
  NAND2_X1 U704 ( .A1(n628), .A2(n622), .ZN(n623) );
  XNOR2_X1 U705 ( .A(n624), .B(n623), .ZN(n625) );
  XOR2_X1 U706 ( .A(G128), .B(n625), .Z(G30) );
  XNOR2_X1 U707 ( .A(G143), .B(n626), .ZN(G45) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U709 ( .A(n629), .B(KEYINPUT110), .ZN(n630) );
  XNOR2_X1 U710 ( .A(G146), .B(n630), .ZN(G48) );
  NOR2_X1 U711 ( .A1(n631), .A2(n633), .ZN(n632) );
  XOR2_X1 U712 ( .A(G113), .B(n632), .Z(G15) );
  NOR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U714 ( .A(G116), .B(n635), .Z(G18) );
  XOR2_X1 U715 ( .A(KEYINPUT37), .B(KEYINPUT111), .Z(n638) );
  XNOR2_X1 U716 ( .A(G125), .B(n636), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n638), .B(n637), .ZN(G27) );
  XOR2_X1 U718 ( .A(G134), .B(n639), .Z(G36) );
  XNOR2_X1 U719 ( .A(G140), .B(n640), .ZN(G42) );
  INV_X1 U720 ( .A(n669), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n641), .A2(n657), .ZN(n688) );
  NAND2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U723 ( .A(KEYINPUT50), .B(n644), .ZN(n649) );
  XOR2_X1 U724 ( .A(KEYINPUT49), .B(KEYINPUT112), .Z(n647) );
  NAND2_X1 U725 ( .A1(n520), .A2(n645), .ZN(n646) );
  XNOR2_X1 U726 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U727 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U728 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n652), .B(KEYINPUT113), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n656) );
  XOR2_X1 U731 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n655) );
  XNOR2_X1 U732 ( .A(n656), .B(n655), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n672) );
  NOR2_X1 U734 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U735 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U736 ( .A(KEYINPUT115), .B(n663), .Z(n667) );
  NOR2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U739 ( .A1(n360), .A2(n668), .ZN(n670) );
  XOR2_X1 U740 ( .A(KEYINPUT116), .B(n670), .Z(n671) );
  NAND2_X1 U741 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U742 ( .A(KEYINPUT52), .B(n673), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n674), .A2(G952), .ZN(n675) );
  NOR2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n677), .B(KEYINPUT117), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n725), .A2(n678), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U748 ( .A(KEYINPUT77), .B(n681), .ZN(n682) );
  NOR2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U750 ( .A(KEYINPUT80), .B(n684), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U753 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n691) );
  NOR2_X1 U754 ( .A1(n707), .A2(n693), .ZN(G54) );
  XOR2_X1 U755 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n694) );
  XOR2_X1 U756 ( .A(KEYINPUT60), .B(KEYINPUT121), .Z(n699) );
  XNOR2_X1 U757 ( .A(n700), .B(n699), .ZN(G60) );
  XNOR2_X1 U758 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U759 ( .A1(n707), .A2(n703), .ZN(G63) );
  XNOR2_X1 U760 ( .A(n704), .B(n705), .ZN(n706) );
  NAND2_X1 U761 ( .A1(n725), .A2(n348), .ZN(n713) );
  NAND2_X1 U762 ( .A1(G953), .A2(G224), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n709), .B(KEYINPUT61), .ZN(n711) );
  NAND2_X1 U764 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n719) );
  XOR2_X1 U766 ( .A(n714), .B(G101), .Z(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U768 ( .A(KEYINPUT123), .B(n717), .Z(n718) );
  XNOR2_X1 U769 ( .A(n719), .B(n718), .ZN(G69) );
  BUF_X1 U770 ( .A(n720), .Z(n721) );
  XOR2_X1 U771 ( .A(n722), .B(n721), .Z(n723) );
  XOR2_X1 U772 ( .A(KEYINPUT124), .B(n723), .Z(n727) );
  XOR2_X1 U773 ( .A(n727), .B(n724), .Z(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n732) );
  XNOR2_X1 U775 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(G900), .ZN(n729) );
  XOR2_X1 U777 ( .A(KEYINPUT125), .B(n729), .Z(n730) );
  NAND2_X1 U778 ( .A1(G953), .A2(n730), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n732), .A2(n731), .ZN(G72) );
  XNOR2_X1 U780 ( .A(n733), .B(KEYINPUT126), .ZN(G21) );
  XOR2_X1 U781 ( .A(n734), .B(G122), .Z(G24) );
  XNOR2_X1 U782 ( .A(n735), .B(G131), .ZN(G33) );
  XNOR2_X1 U783 ( .A(G137), .B(n736), .ZN(G39) );
  XOR2_X1 U784 ( .A(n737), .B(G101), .Z(n738) );
  XNOR2_X1 U785 ( .A(KEYINPUT108), .B(n738), .ZN(G3) );
endmodule

