//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910;
  XNOR2_X1  g000(.A(G141gat), .B(G148gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  AND2_X1   g002(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT80), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G155gat), .B2(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n211), .A2(KEYINPUT81), .A3(new_n203), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT81), .B1(new_n211), .B2(new_n203), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n202), .A2(KEYINPUT82), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n206), .A2(new_n207), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n203), .B1(new_n216), .B2(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT82), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n214), .A2(new_n222), .A3(new_n219), .ZN(new_n223));
  XNOR2_X1  g022(.A(G113gat), .B(G120gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XOR2_X1   g024(.A(G127gat), .B(G134gat), .Z(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G225gat), .A2(G233gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n214), .A3(new_n219), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT4), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n227), .A2(new_n214), .A3(KEYINPUT4), .A4(new_n219), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n229), .A2(new_n230), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT83), .ZN(new_n236));
  OR3_X1    g035(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT5), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n235), .B2(KEYINPUT5), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT5), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n228), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n231), .ZN(new_n242));
  INV_X1    g041(.A(new_n230), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n235), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G1gat), .B(G29gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT0), .ZN(new_n248));
  XNOR2_X1  g047(.A(G57gat), .B(G85gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n233), .A3(new_n234), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n243), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n254), .B(KEYINPUT39), .C1(new_n243), .C2(new_n242), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n250), .B1(new_n254), .B2(KEYINPUT39), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n256), .A2(KEYINPUT88), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(KEYINPUT88), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT40), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n252), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n260), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT89), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT89), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n264), .A3(new_n260), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G8gat), .B(G36gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT78), .ZN(new_n268));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271));
  INV_X1    g070(.A(G211gat), .ZN(new_n272));
  INV_X1    g071(.A(G218gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n271), .B1(KEYINPUT22), .B2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G211gat), .B(G218gat), .Z(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT25), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n281));
  INV_X1    g080(.A(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n283), .A2(KEYINPUT23), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n290), .A2(new_n291), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n289), .B(new_n292), .C1(new_n293), .C2(KEYINPUT24), .ZN(new_n294));
  NAND2_X1  g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n284), .A2(new_n282), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n280), .B1(new_n288), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT66), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT65), .ZN(new_n302));
  INV_X1    g101(.A(new_n299), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT25), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n293), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT24), .B1(new_n307), .B2(KEYINPUT67), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(KEYINPUT67), .B2(new_n307), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n289), .A2(KEYINPUT68), .B1(new_n290), .B2(new_n291), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n309), .B(new_n310), .C1(KEYINPUT68), .C2(new_n289), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT25), .B1(new_n297), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(new_n297), .B2(new_n296), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n301), .A2(new_n306), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT26), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n297), .A2(new_n316), .A3(new_n295), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n317), .B(new_n307), .C1(new_n316), .C2(new_n297), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT72), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT69), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(G183gat), .ZN(new_n324));
  AOI21_X1  g123(.A(G190gat), .B1(new_n323), .B2(G183gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n290), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n331), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n290), .A2(KEYINPUT27), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n325), .A2(KEYINPUT28), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n321), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n327), .A2(new_n331), .A3(new_n328), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n331), .B1(new_n327), .B2(new_n328), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n321), .B(new_n335), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n320), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT73), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT71), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n339), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n320), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n315), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n279), .B1(new_n348), .B2(KEYINPUT29), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n311), .A2(new_n314), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n300), .A2(KEYINPUT66), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n304), .A2(new_n305), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n341), .ZN(new_n355));
  INV_X1    g154(.A(new_n279), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n350), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(KEYINPUT77), .B(new_n279), .C1(new_n348), .C2(KEYINPUT29), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n278), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n347), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n356), .A3(new_n354), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(new_n364), .A3(new_n279), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n277), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n270), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n346), .B1(new_n345), .B2(new_n320), .ZN(new_n368));
  AOI211_X1 g167(.A(KEYINPUT73), .B(new_n319), .C1(new_n344), .C2(new_n339), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n354), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n364), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n357), .B1(new_n371), .B2(new_n279), .ZN(new_n372));
  AOI211_X1 g171(.A(new_n350), .B(new_n356), .C1(new_n370), .C2(new_n364), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n277), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n366), .ZN(new_n375));
  INV_X1    g174(.A(new_n270), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n374), .A2(KEYINPUT30), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n356), .B1(new_n370), .B2(new_n364), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n360), .B1(new_n378), .B2(new_n357), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n366), .B1(new_n379), .B2(new_n277), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT30), .B1(new_n380), .B2(new_n376), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n367), .B(new_n377), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  AOI211_X1 g182(.A(new_n366), .B(new_n270), .C1(new_n379), .C2(new_n277), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n384), .A2(KEYINPUT79), .A3(KEYINPUT30), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n266), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n277), .A2(KEYINPUT85), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n275), .A2(new_n276), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n387), .B(new_n364), .C1(KEYINPUT85), .C2(new_n388), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n389), .A2(new_n222), .B1(new_n214), .B2(new_n219), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n278), .B1(new_n364), .B2(new_n223), .ZN(new_n391));
  INV_X1    g190(.A(G228gat), .ZN(new_n392));
  INV_X1    g191(.A(G233gat), .ZN(new_n393));
  OAI22_X1  g192(.A1(new_n390), .A2(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n222), .B1(new_n277), .B2(KEYINPUT29), .ZN(new_n395));
  AOI211_X1 g194(.A(new_n392), .B(new_n393), .C1(new_n395), .C2(new_n220), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n396), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n391), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(KEYINPUT86), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n394), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G22gat), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n394), .B(new_n403), .C1(new_n398), .C2(new_n400), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT87), .B1(new_n401), .B2(G22gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(G50gat), .ZN(new_n408));
  XOR2_X1   g207(.A(G78gat), .B(G106gat), .Z(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n405), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n402), .A2(KEYINPUT87), .A3(new_n404), .A4(new_n410), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT37), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n374), .A2(new_n415), .A3(new_n375), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n270), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n380), .A2(new_n415), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT38), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n237), .A2(new_n238), .B1(new_n235), .B2(new_n244), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT6), .B1(new_n420), .B2(new_n250), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n252), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n246), .A2(KEYINPUT6), .A3(new_n251), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(new_n384), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n363), .A2(new_n277), .A3(new_n365), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT90), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n360), .B(new_n278), .C1(new_n378), .C2(new_n357), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT37), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT38), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n430), .A2(new_n431), .A3(new_n270), .A4(new_n416), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n419), .A2(new_n425), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n386), .A2(new_n414), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n367), .A2(new_n377), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT79), .B1(new_n384), .B2(KEYINPUT30), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n380), .A2(new_n376), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n382), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n435), .A2(new_n436), .A3(new_n439), .A4(new_n424), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n412), .A2(new_n413), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  XNOR2_X1  g242(.A(G15gat), .B(G43gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT75), .ZN(new_n445));
  XNOR2_X1  g244(.A(G71gat), .B(G99gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n227), .B1(new_n362), .B2(new_n354), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n228), .B(new_n315), .C1(new_n342), .C2(new_n347), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT74), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n455), .A3(KEYINPUT32), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n370), .A2(new_n228), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n362), .A2(new_n227), .A3(new_n354), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n448), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT32), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT74), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n454), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(new_n458), .A3(new_n448), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT76), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT34), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n463), .B2(new_n464), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n452), .B(KEYINPUT32), .C1(new_n453), .C2(new_n447), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n462), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n462), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n443), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n462), .A2(new_n469), .ZN(new_n473));
  INV_X1    g272(.A(new_n468), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n462), .A2(new_n468), .A3(new_n469), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(KEYINPUT36), .A3(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n434), .A2(new_n442), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT91), .B(new_n414), .C1(new_n470), .C2(new_n471), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(new_n440), .ZN(new_n482));
  AND4_X1   g281(.A1(new_n424), .A2(new_n435), .A3(new_n436), .A4(new_n439), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n441), .B1(new_n475), .B2(new_n476), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT91), .A4(KEYINPUT35), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n479), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT16), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(G1gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(G1gat), .B2(new_n487), .ZN(new_n490));
  INV_X1    g289(.A(G8gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(G29gat), .A2(G36gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT14), .ZN(new_n494));
  NAND2_X1  g293(.A1(G29gat), .A2(G36gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT92), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n497), .A2(KEYINPUT93), .B1(KEYINPUT15), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(KEYINPUT15), .B2(new_n498), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n500), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n501), .A2(KEYINPUT17), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT17), .B1(new_n501), .B2(new_n502), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n492), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n492), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(new_n501), .A3(new_n502), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n501), .A2(new_n502), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n492), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n508), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n506), .B(KEYINPUT13), .Z(new_n513));
  AOI22_X1  g312(.A1(new_n509), .A2(KEYINPUT18), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT94), .B1(new_n509), .B2(KEYINPUT18), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n514), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G197gat), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT11), .B(G169gat), .Z(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(KEYINPUT12), .Z(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n525), .B1(new_n516), .B2(new_n518), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n514), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(KEYINPUT95), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT95), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n520), .A2(new_n530), .A3(new_n525), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT9), .ZN(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(G71gat), .A2(G78gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT96), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  OR3_X1    g340(.A1(new_n537), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n539), .B1(new_n537), .B2(new_n541), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G127gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(KEYINPUT99), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n507), .B1(new_n554), .B2(KEYINPUT21), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n550), .B(new_n555), .Z(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT98), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G155gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT100), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n559), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n556), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT102), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(KEYINPUT102), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(KEYINPUT7), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT103), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT104), .B(G85gat), .Z(new_n573));
  XOR2_X1   g372(.A(KEYINPUT105), .B(G92gat), .Z(new_n574));
  OAI221_X1 g373(.A(new_n566), .B1(new_n571), .B2(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G99gat), .B(G106gat), .Z(new_n576));
  OR2_X1    g375(.A1(new_n567), .A2(KEYINPUT7), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  OR3_X1    g377(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n576), .B1(new_n575), .B2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(KEYINPUT106), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(KEYINPUT106), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n582), .B(new_n583), .C1(new_n503), .C2(new_n504), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT107), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n510), .A2(new_n581), .ZN(new_n588));
  AND2_X1   g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(KEYINPUT41), .B2(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n584), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n587), .B1(new_n584), .B2(new_n590), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(KEYINPUT41), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT101), .Z(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OR3_X1    g396(.A1(new_n591), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n591), .B2(new_n592), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n564), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT109), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n579), .A2(new_n580), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n545), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n581), .A2(new_n544), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT10), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND4_X1   g405(.A1(KEYINPUT10), .A2(new_n603), .A3(new_n551), .A4(new_n553), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT108), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n602), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  OAI211_X1 g411(.A(KEYINPUT109), .B(new_n612), .C1(new_n606), .C2(new_n607), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n604), .A2(new_n605), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n612), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n610), .B(KEYINPUT110), .Z(new_n623));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n620), .B1(new_n624), .B2(new_n616), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AND4_X1   g426(.A1(new_n486), .A2(new_n533), .A3(new_n601), .A4(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n424), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g430(.A1(new_n383), .A2(new_n385), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT16), .B(G8gat), .Z(new_n635));
  AND2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n634), .A2(new_n491), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT42), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(KEYINPUT42), .B2(new_n636), .ZN(G1325gat));
  INV_X1    g438(.A(G15gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n475), .A2(new_n476), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n628), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n478), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n628), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n644), .B2(new_n640), .ZN(G1326gat));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n441), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT43), .B(G22gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1327gat));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n486), .B2(new_n600), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n600), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n485), .A2(new_n482), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n479), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n563), .A2(new_n532), .A3(new_n626), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G29gat), .B1(new_n659), .B2(new_n424), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(new_n658), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n424), .A2(G29gat), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n661), .A2(KEYINPUT111), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT45), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT111), .B1(new_n661), .B2(new_n662), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n663), .B2(new_n665), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n660), .B1(new_n666), .B2(new_n667), .ZN(G1328gat));
  NOR3_X1   g467(.A1(new_n661), .A2(G36gat), .A3(new_n632), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT46), .ZN(new_n670));
  OAI21_X1  g469(.A(G36gat), .B1(new_n659), .B2(new_n632), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(G1329gat));
  INV_X1    g471(.A(new_n658), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n651), .B2(new_n656), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(G43gat), .A3(new_n643), .ZN(new_n675));
  INV_X1    g474(.A(G43gat), .ZN(new_n676));
  INV_X1    g475(.A(new_n641), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n661), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT47), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT47), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n675), .A2(new_n681), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(G1330gat));
  OAI21_X1  g482(.A(G50gat), .B1(new_n659), .B2(new_n414), .ZN(new_n684));
  INV_X1    g483(.A(new_n661), .ZN(new_n685));
  INV_X1    g484(.A(G50gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n441), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT113), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n684), .A2(KEYINPUT48), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT48), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n686), .B1(new_n674), .B2(new_n441), .ZN(new_n692));
  INV_X1    g491(.A(new_n689), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n694), .ZN(G1331gat));
  NAND3_X1  g494(.A1(new_n601), .A2(new_n532), .A3(new_n626), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n653), .B2(new_n479), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n629), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g498(.A(new_n632), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT114), .ZN(new_n702));
  NOR2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1333gat));
  NAND2_X1  g503(.A1(new_n697), .A2(new_n643), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n677), .A2(G71gat), .ZN(new_n706));
  AOI22_X1  g505(.A1(new_n705), .A2(G71gat), .B1(new_n697), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g507(.A1(new_n697), .A2(new_n441), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g509(.A1(new_n533), .A2(new_n563), .A3(new_n627), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n657), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n573), .B1(new_n712), .B2(new_n424), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT115), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n533), .A2(new_n563), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n654), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n654), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n715), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n627), .A2(new_n424), .A3(new_n573), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n713), .A2(new_n723), .ZN(G1336gat));
  NOR3_X1   g523(.A1(new_n632), .A2(G92gat), .A3(new_n627), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n717), .A2(KEYINPUT116), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n654), .B2(new_n715), .ZN(new_n727));
  AND4_X1   g526(.A1(new_n486), .A2(new_n600), .A3(new_n715), .A4(new_n726), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT117), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT117), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n731), .B(new_n725), .C1(new_n727), .C2(new_n728), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n486), .A2(new_n600), .A3(new_n655), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n633), .B(new_n711), .C1(new_n733), .C2(new_n650), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n574), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n730), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT52), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n725), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n739), .A3(new_n735), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n712), .B2(new_n478), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n677), .A2(G99gat), .A3(new_n627), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n721), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1338gat));
  NOR3_X1   g544(.A1(new_n627), .A2(new_n414), .A3(G106gat), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n721), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n441), .B(new_n711), .C1(new_n733), .C2(new_n650), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G106gat), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n727), .A2(new_n728), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n752), .A2(new_n746), .B1(new_n748), .B2(G106gat), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n747), .A2(new_n751), .B1(new_n753), .B2(new_n750), .ZN(G1339gat));
  INV_X1    g553(.A(new_n484), .ZN(new_n755));
  INV_X1    g554(.A(new_n623), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n606), .B2(new_n607), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n620), .B1(new_n757), .B2(KEYINPUT54), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n608), .B2(new_n623), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n758), .B1(new_n614), .B2(new_n760), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n761), .A2(KEYINPUT55), .B1(new_n614), .B2(new_n621), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT10), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n615), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n607), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n766), .A3(new_n623), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT54), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n611), .B2(new_n613), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n763), .B1(new_n769), .B2(new_n758), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n762), .A2(new_n529), .A3(new_n531), .A4(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n512), .B2(new_n513), .ZN(new_n773));
  INV_X1    g572(.A(new_n513), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n511), .A2(KEYINPUT118), .A3(new_n508), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n506), .B1(new_n505), .B2(new_n508), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n524), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n626), .A2(new_n780), .A3(new_n528), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n600), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n770), .A2(new_n600), .A3(new_n780), .A4(new_n528), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n761), .A2(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n622), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n564), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n601), .A2(new_n532), .A3(new_n627), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n755), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n629), .A3(new_n632), .ZN(new_n790));
  INV_X1    g589(.A(G113gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n790), .A2(new_n791), .A3(new_n532), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n424), .B1(new_n787), .B2(new_n788), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(new_n484), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(new_n632), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n533), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n792), .B1(new_n796), .B2(new_n791), .ZN(G1340gat));
  NOR2_X1   g596(.A1(new_n627), .A2(G120gat), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT120), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G120gat), .B1(new_n790), .B2(new_n627), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1341gat));
  INV_X1    g601(.A(G127gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n795), .A2(new_n803), .A3(new_n563), .ZN(new_n804));
  OAI21_X1  g603(.A(G127gat), .B1(new_n790), .B2(new_n564), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1342gat));
  INV_X1    g607(.A(G134gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n632), .A2(new_n600), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT122), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n812), .A2(KEYINPUT56), .ZN(new_n813));
  OAI21_X1  g612(.A(G134gat), .B1(new_n790), .B2(new_n652), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(KEYINPUT56), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(G1343gat));
  INV_X1    g615(.A(G141gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n529), .A2(new_n770), .A3(new_n531), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n781), .B1(new_n818), .B2(new_n785), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n786), .B1(new_n819), .B2(new_n652), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n788), .B1(new_n820), .B2(new_n563), .ZN(new_n821));
  AND4_X1   g620(.A1(new_n629), .A2(new_n821), .A3(new_n441), .A4(new_n478), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n632), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n817), .B1(new_n823), .B2(new_n532), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n414), .B1(new_n787), .B2(new_n788), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT57), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n643), .A2(new_n633), .A3(new_n424), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n532), .A2(new_n817), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n824), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(G1344gat));
  INV_X1    g632(.A(new_n823), .ZN(new_n834));
  INV_X1    g633(.A(G148gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n626), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n826), .A2(new_n827), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT59), .B(new_n835), .C1(new_n837), .C2(new_n626), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n821), .A2(KEYINPUT57), .A3(new_n441), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(KEYINPUT123), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n825), .B2(KEYINPUT57), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n819), .A2(new_n652), .ZN(new_n844));
  INV_X1    g643(.A(new_n786), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(KEYINPUT124), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n782), .B2(new_n786), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n848), .A3(new_n564), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n414), .B1(new_n849), .B2(new_n788), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n841), .A2(new_n843), .B1(new_n850), .B2(KEYINPUT57), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n626), .A3(new_n827), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n839), .B1(new_n852), .B2(G148gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n836), .B1(new_n838), .B2(new_n853), .ZN(G1345gat));
  OAI21_X1  g653(.A(G155gat), .B1(new_n828), .B2(new_n564), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n834), .A2(new_n206), .A3(new_n563), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1346gat));
  OAI21_X1  g656(.A(G162gat), .B1(new_n828), .B2(new_n652), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n822), .A2(new_n207), .A3(new_n811), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1347gat));
  NOR2_X1   g659(.A1(new_n632), .A2(new_n629), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n789), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(new_n284), .A3(new_n532), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n629), .B1(new_n787), .B2(new_n788), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n755), .A2(new_n632), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n533), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n863), .B1(new_n284), .B2(new_n868), .ZN(G1348gat));
  OAI21_X1  g668(.A(new_n282), .B1(new_n866), .B2(new_n627), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n283), .A2(new_n285), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n626), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n862), .B2(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT125), .Z(G1349gat));
  OAI21_X1  g673(.A(G183gat), .B1(new_n862), .B2(new_n564), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n323), .A2(G183gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n563), .A2(new_n334), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n866), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g678(.A1(new_n867), .A2(new_n291), .A3(new_n600), .ZN(new_n880));
  OAI21_X1  g679(.A(G190gat), .B1(new_n862), .B2(new_n652), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(KEYINPUT61), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(KEYINPUT61), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(G1351gat));
  NOR3_X1   g683(.A1(new_n643), .A2(new_n414), .A3(new_n632), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(KEYINPUT126), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(KEYINPUT126), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n864), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(KEYINPUT127), .B(G197gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n533), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n851), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n478), .A2(new_n861), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n532), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n894), .B2(new_n890), .ZN(G1352gat));
  NOR3_X1   g694(.A1(new_n888), .A2(G204gat), .A3(new_n627), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n892), .A2(new_n627), .A3(new_n893), .ZN(new_n900));
  INV_X1    g699(.A(G204gat), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n898), .B(new_n899), .C1(new_n900), .C2(new_n901), .ZN(G1353gat));
  NAND3_X1  g701(.A1(new_n889), .A2(new_n272), .A3(new_n563), .ZN(new_n903));
  INV_X1    g702(.A(new_n893), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n851), .A2(new_n563), .A3(new_n904), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n905), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT63), .B1(new_n905), .B2(G211gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G1354gat));
  NAND3_X1  g707(.A1(new_n889), .A2(new_n273), .A3(new_n600), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n892), .A2(new_n652), .A3(new_n893), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n273), .ZN(G1355gat));
endmodule


