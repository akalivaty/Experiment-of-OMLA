//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT64), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n461), .A2(KEYINPUT65), .A3(G101), .A4(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  OAI211_X1 g051(.A(G137), .B(new_n461), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT66), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n474), .A2(new_n480), .A3(new_n477), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n469), .B1(new_n479), .B2(new_n481), .ZN(G160));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g059(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G112), .B2(new_n461), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n466), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  AOI21_X1  g064(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OAI221_X1 g066(.A(new_n486), .B1(new_n487), .B2(new_n488), .C1(new_n489), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NOR2_X1   g068(.A1(new_n461), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n497), .A2(new_n461), .A3(KEYINPUT4), .A4(G138), .ZN(new_n498));
  NAND2_X1  g073(.A1(G126), .A2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n500), .B2(new_n466), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n461), .C1(new_n475), .C2(new_n476), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(KEYINPUT68), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT69), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT69), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n513), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n515), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(G166));
  NAND2_X1  g101(.A1(new_n520), .A2(KEYINPUT70), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n521), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n517), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(G168));
  NAND3_X1  g117(.A1(new_n527), .A2(new_n532), .A3(G64), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n524), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n514), .A2(G52), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n547), .B2(new_n521), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n533), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n524), .B1(new_n552), .B2(KEYINPUT71), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n553), .B1(KEYINPUT71), .B2(new_n552), .ZN(new_n554));
  INV_X1    g129(.A(new_n521), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G81), .B1(G43), .B2(new_n514), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n539), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n514), .A2(new_n563), .A3(new_n566), .A4(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n530), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n565), .A2(new_n567), .B1(G651), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n555), .A2(KEYINPUT73), .A3(G91), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n521), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n571), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  NAND3_X1  g155(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n521), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n533), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n583), .B1(new_n585), .B2(G651), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G288));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n518), .B2(new_n519), .ZN(new_n589));
  AND2_X1   g164(.A1(G73), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n517), .A2(new_n520), .A3(G86), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n555), .A2(G85), .B1(G47), .B2(new_n514), .ZN(new_n595));
  INV_X1    g170(.A(G60), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n533), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n595), .B1(new_n598), .B2(new_n524), .ZN(G290));
  AND3_X1   g174(.A1(new_n517), .A2(G92), .A3(new_n520), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT74), .B(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n530), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G321));
  NOR2_X1   g185(.A1(G286), .A2(new_n607), .ZN(new_n611));
  XNOR2_X1  g186(.A(G299), .B(KEYINPUT75), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n607), .ZN(G297));
  XOR2_X1   g188(.A(G297), .B(KEYINPUT76), .Z(G280));
  INV_X1    g189(.A(new_n606), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n554), .A2(new_n556), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n607), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n606), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n607), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g197(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n623));
  NOR3_X1   g198(.A1(new_n462), .A2(new_n463), .A3(G2105), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n623), .B(new_n624), .Z(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n490), .A2(G135), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n461), .A2(G111), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G123), .ZN(new_n634));
  OAI221_X1 g209(.A(new_n631), .B1(new_n632), .B2(new_n633), .C1(new_n634), .C2(new_n488), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT79), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT80), .ZN(new_n652));
  OAI21_X1  g227(.A(G14), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  AOI21_X1  g234(.A(new_n657), .B1(new_n656), .B2(KEYINPUT81), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(KEYINPUT81), .B2(new_n656), .ZN(new_n661));
  INV_X1    g236(.A(new_n655), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n656), .B(KEYINPUT17), .Z(new_n663));
  INV_X1    g238(.A(new_n657), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n661), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n655), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n659), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT82), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT83), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g256(.A(new_n681), .B(new_n680), .S(new_n673), .Z(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT85), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT84), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n694), .A2(G33), .ZN(new_n695));
  AND3_X1   g270(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT25), .ZN(new_n697));
  INV_X1    g272(.A(G139), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n491), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT91), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(new_n461), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n695), .B1(new_n704), .B2(G29), .ZN(new_n705));
  INV_X1    g280(.A(G2072), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NOR2_X1   g284(.A1(G168), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n709), .B2(G21), .ZN(new_n711));
  INV_X1    g286(.A(G1966), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G34), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(KEYINPUT24), .ZN(new_n715));
  AOI21_X1  g290(.A(G29), .B1(new_n714), .B2(KEYINPUT24), .ZN(new_n716));
  AOI22_X1  g291(.A1(G160), .A2(G29), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(G2084), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n705), .B2(new_n706), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n709), .A2(G5), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G171), .B2(new_n709), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(G1961), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n694), .A2(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n694), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2078), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n722), .B1(KEYINPUT95), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT30), .B(G28), .ZN(new_n727));
  OR2_X1    g302(.A1(KEYINPUT31), .A2(G11), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n727), .A2(new_n694), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n635), .B2(new_n694), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n711), .B2(new_n712), .ZN(new_n732));
  AND4_X1   g307(.A1(new_n713), .A2(new_n719), .A3(new_n726), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n694), .A2(G32), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n475), .A2(new_n476), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n461), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G129), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT93), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT26), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n739), .B(new_n741), .C1(G141), .C2(new_n490), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n738), .A2(KEYINPUT94), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(KEYINPUT94), .B1(new_n738), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n734), .B1(new_n745), .B2(new_n694), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n721), .A2(G1961), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n725), .B2(KEYINPUT95), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G2084), .B2(new_n717), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n708), .A2(new_n733), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(KEYINPUT96), .ZN(new_n753));
  NOR2_X1   g328(.A1(G16), .A2(G19), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n557), .B2(G16), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1341), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n694), .A2(G35), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G162), .B2(new_n694), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2090), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT97), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n615), .A2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G4), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n694), .A2(G26), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT28), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n736), .A2(G128), .B1(G140), .B2(new_n490), .ZN(new_n771));
  OAI21_X1  g346(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NOR3_X1   g348(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n774));
  OAI221_X1 g349(.A(G2104), .B1(G116), .B2(new_n461), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n767), .A2(new_n768), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n756), .A2(new_n763), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n760), .A2(new_n761), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n709), .A2(G20), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT23), .Z(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G299), .B2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G1956), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(KEYINPUT98), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(KEYINPUT98), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n781), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n752), .A2(KEYINPUT96), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n753), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT99), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(KEYINPUT99), .ZN(new_n796));
  NOR2_X1   g371(.A1(G6), .A2(G16), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT32), .ZN(new_n800));
  INV_X1    g375(.A(G1981), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n709), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n709), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT88), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(KEYINPUT88), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n709), .A2(G23), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n586), .B2(new_n709), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT33), .B(G1976), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n802), .A2(new_n807), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n815));
  MUX2_X1   g390(.A(G24), .B(G290), .S(G16), .Z(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1986), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n694), .A2(G25), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n490), .A2(G131), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n461), .A2(G107), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n821));
  INV_X1    g396(.A(G119), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n819), .B1(new_n820), .B2(new_n821), .C1(new_n822), .C2(new_n488), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(KEYINPUT86), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(KEYINPUT86), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n818), .B1(new_n827), .B2(new_n694), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT35), .B(G1991), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT87), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n814), .A2(new_n815), .A3(new_n817), .A4(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT89), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n834), .B1(new_n832), .B2(new_n833), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n832), .A2(new_n833), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n795), .A2(new_n796), .B1(new_n837), .B2(new_n838), .ZN(G311));
  NAND2_X1  g414(.A1(new_n795), .A2(new_n796), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n835), .B2(new_n836), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(G150));
  NAND2_X1  g417(.A1(new_n615), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n514), .A2(G55), .ZN(new_n845));
  INV_X1    g420(.A(G93), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n521), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n533), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n847), .B1(new_n850), .B2(G651), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n554), .B2(new_n556), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n554), .A2(new_n556), .A3(new_n851), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n844), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  INV_X1    g434(.A(new_n851), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT100), .Z(G145));
  XNOR2_X1  g439(.A(G160), .B(new_n492), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n635), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n776), .B(new_n507), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n738), .A2(new_n742), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n704), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n743), .B2(new_n744), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT94), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n738), .A2(KEYINPUT94), .A3(new_n742), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(KEYINPUT101), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n868), .B(new_n870), .C1(new_n877), .C2(new_n704), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n736), .A2(G130), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n490), .A2(G142), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n826), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n824), .B2(new_n825), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n625), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n625), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n885), .B2(new_n887), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n704), .B1(new_n872), .B2(new_n876), .ZN(new_n893));
  INV_X1    g468(.A(new_n870), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n867), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n878), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n878), .A2(new_n895), .ZN(new_n899));
  INV_X1    g474(.A(new_n892), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n897), .A3(new_n900), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n866), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G37), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n896), .A2(new_n866), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n892), .B1(new_n878), .B2(new_n895), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT103), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n866), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n907), .B1(new_n897), .B2(new_n896), .ZN(new_n911));
  INV_X1    g486(.A(new_n903), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n908), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n909), .A2(new_n916), .A3(KEYINPUT40), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT40), .B1(new_n909), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(G395));
  NOR2_X1   g494(.A1(new_n855), .A2(new_n620), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n855), .A2(new_n620), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n615), .A2(G299), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n571), .A2(new_n576), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n606), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n924), .B1(new_n923), .B2(new_n606), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR3_X1    g503(.A1(new_n920), .A2(new_n921), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT41), .B1(new_n926), .B2(new_n927), .ZN(new_n930));
  INV_X1    g505(.A(new_n927), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n922), .A4(new_n925), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n921), .B2(new_n920), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n937));
  XNOR2_X1  g512(.A(G166), .B(KEYINPUT105), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(G305), .ZN(new_n939));
  XNOR2_X1  g514(.A(G290), .B(new_n586), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n939), .B(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n929), .A2(new_n935), .A3(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n937), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n937), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g520(.A(G868), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(G868), .B2(new_n851), .ZN(G295));
  OAI21_X1  g522(.A(new_n946), .B1(G868), .B2(new_n851), .ZN(G331));
  OAI21_X1  g523(.A(KEYINPUT106), .B1(new_n545), .B2(new_n548), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n545), .A2(KEYINPUT106), .A3(new_n548), .ZN(new_n951));
  OAI21_X1  g526(.A(G286), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n951), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(G168), .A3(new_n949), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n853), .A3(new_n854), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n554), .A2(new_n556), .A3(new_n851), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n954), .B(new_n952), .C1(new_n957), .C2(new_n852), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n955), .A2(new_n853), .A3(KEYINPUT107), .A4(new_n854), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n934), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n956), .B(new_n958), .C1(new_n927), .C2(new_n926), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n941), .A3(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n964), .A2(new_n905), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  INV_X1    g542(.A(new_n941), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n928), .B1(new_n960), .B2(new_n961), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n930), .A2(new_n933), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n956), .B2(new_n958), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n968), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n972), .A2(new_n967), .A3(new_n964), .A4(new_n905), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n964), .A2(new_n905), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n941), .B1(new_n962), .B2(new_n963), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT43), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n972), .A2(new_n905), .A3(new_n964), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n982), .B2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g558(.A(new_n977), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n965), .A2(new_n967), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT109), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n983), .A2(KEYINPUT109), .A3(new_n985), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n981), .B1(new_n986), .B2(new_n987), .ZN(G397));
  INV_X1    g563(.A(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n467), .A2(new_n468), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G2105), .ZN(new_n991));
  INV_X1    g566(.A(new_n481), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n480), .B1(new_n474), .B2(new_n477), .ZN(new_n993));
  OAI211_X1 g568(.A(G40), .B(new_n991), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n494), .A2(new_n495), .ZN(new_n996));
  INV_X1    g571(.A(new_n499), .ZN(new_n997));
  INV_X1    g572(.A(G138), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(G2105), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n504), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n996), .B1(new_n1000), .B2(new_n735), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n504), .B1(new_n490), .B2(G138), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n995), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n994), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1996), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n745), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n776), .A2(G2067), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n771), .A2(new_n778), .A3(new_n775), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(G1996), .B2(new_n869), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n826), .B(new_n830), .Z(new_n1014));
  OAI21_X1  g589(.A(new_n1006), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(G290), .A2(G1986), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G290), .A2(G1986), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1006), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT110), .Z(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT116), .B(KEYINPUT63), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n994), .A2(new_n1003), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT112), .B1(new_n586), .B2(G1976), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n585), .A2(G651), .ZN(new_n1027));
  INV_X1    g602(.A(new_n583), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1976), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1025), .B(new_n1026), .C1(KEYINPUT52), .C2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n501), .B2(new_n506), .ZN(new_n1031));
  NAND3_X1  g606(.A1(G160), .A2(G40), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1026), .A2(new_n1032), .A3(G8), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(G8), .A3(new_n1029), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n801), .B1(new_n591), .B2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1039), .A2(G305), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(G305), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT114), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n593), .A2(new_n592), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1044), .B(new_n591), .C1(new_n1038), .C2(new_n801), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1039), .A2(G305), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT49), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1032), .B(G8), .C1(new_n1051), .C2(new_n1037), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1030), .A2(new_n1036), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1031), .A2(KEYINPUT45), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1005), .A2(G160), .A3(new_n1055), .A4(G40), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n805), .ZN(new_n1057));
  INV_X1    g632(.A(G40), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1058), .B(new_n469), .C1(new_n479), .C2(new_n481), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n507), .A2(new_n1061), .A3(new_n995), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1059), .A2(new_n761), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1024), .B1(new_n1057), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(G166), .B2(new_n1024), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1065), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT45), .B1(new_n507), .B2(new_n995), .ZN(new_n1073));
  AOI211_X1 g648(.A(new_n1004), .B(G1384), .C1(new_n501), .C2(new_n506), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n994), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1063), .B1(new_n1075), .B2(G1971), .ZN(new_n1076));
  AND4_X1   g651(.A1(new_n1072), .A2(new_n1076), .A3(G8), .A4(new_n1069), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1072), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1054), .B(new_n1071), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1060), .A2(G160), .A3(G40), .A4(new_n1062), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1075), .A2(G1966), .B1(new_n1080), .B2(G2084), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(G286), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1022), .B1(new_n1079), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1076), .A2(new_n1069), .A3(G8), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT111), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1064), .A2(new_n1072), .A3(new_n1069), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1087), .A2(new_n1088), .B1(new_n1070), .B2(new_n1065), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1054), .A4(new_n1083), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G288), .A2(G1976), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1047), .B(KEYINPUT114), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1052), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n798), .A2(new_n801), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT115), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1092), .A2(new_n1054), .B1(new_n1098), .B2(new_n1025), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1085), .A2(new_n1091), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1056), .B2(G2078), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(G2078), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1075), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1961), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1080), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1102), .A2(new_n1104), .A3(G301), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT54), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1059), .A2(KEYINPUT123), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n994), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1103), .A4(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1108), .B1(G171), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1079), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(KEYINPUT51), .B(G8), .C1(new_n1081), .C2(G286), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1056), .A2(new_n712), .ZN(new_n1120));
  INV_X1    g695(.A(G2084), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1059), .A2(new_n1121), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1024), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G168), .A2(new_n1024), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT121), .B(KEYINPUT51), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1124), .A2(KEYINPUT51), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1082), .A2(KEYINPUT122), .A3(new_n1127), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1119), .A2(new_n1125), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1081), .A2(new_n1124), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(G301), .A4(new_n1113), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT124), .B1(new_n1114), .B2(G171), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1102), .A2(new_n1106), .A3(new_n1104), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(G171), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1116), .A2(new_n1133), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1080), .A2(new_n786), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT56), .B(G2072), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1110), .A2(new_n1059), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1144), .A2(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1032), .A2(G2067), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1080), .A2(new_n766), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n606), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1144), .A2(new_n1146), .A3(new_n1149), .A4(new_n1148), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1150), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT118), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT61), .B1(new_n1150), .B2(KEYINPUT118), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT119), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT119), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1161), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1153), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1168), .A2(new_n615), .A3(new_n1151), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT60), .B1(new_n1169), .B2(new_n1154), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT58), .B(G1341), .Z(new_n1171));
  AOI22_X1  g746(.A1(new_n1075), .A2(new_n1007), .B1(new_n1032), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(KEYINPUT117), .B(KEYINPUT59), .C1(new_n1172), .C2(new_n618), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1032), .A2(new_n1171), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(G1996), .B2(new_n1056), .ZN(new_n1175));
  NAND2_X1  g750(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1175), .A2(new_n557), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1168), .A2(new_n1151), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1173), .A2(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1182), .A2(new_n1183), .A3(new_n1155), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1182), .B2(new_n1155), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1170), .B(new_n1180), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1156), .B1(new_n1167), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1100), .B1(new_n1143), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1133), .A2(KEYINPUT62), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1131), .A2(new_n1190), .A3(new_n1132), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1079), .A2(new_n1139), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1021), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n827), .A2(new_n830), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT125), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1010), .B1(new_n1196), .B2(new_n1013), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n1006), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1017), .A2(new_n1006), .ZN(new_n1199));
  XOR2_X1   g774(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1200));
  XNOR2_X1  g775(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1015), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1198), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1204), .A2(KEYINPUT46), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(KEYINPUT46), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1011), .A2(new_n869), .ZN(new_n1207));
  AOI22_X1  g782(.A1(new_n1205), .A2(new_n1206), .B1(new_n1006), .B2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1203), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n989), .B1(new_n1194), .B2(new_n1211), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1085), .A2(new_n1091), .A3(new_n1099), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1156), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1186), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1166), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1165), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1214), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1116), .A2(new_n1133), .A3(new_n1142), .ZN(new_n1220));
  OAI211_X1 g795(.A(new_n1193), .B(new_n1213), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1221), .A2(new_n1020), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1222), .A2(KEYINPUT127), .A3(new_n1210), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1212), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g799(.A1(G227), .A2(new_n459), .ZN(new_n1226));
  OAI211_X1 g800(.A(new_n1226), .B(new_n692), .C1(new_n652), .C2(new_n653), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n909), .B2(new_n916), .ZN(new_n1228));
  AND2_X1   g802(.A1(new_n1228), .A2(new_n979), .ZN(G308));
  NAND2_X1  g803(.A1(new_n1228), .A2(new_n979), .ZN(G225));
endmodule


