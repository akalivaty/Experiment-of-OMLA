//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G97), .A2(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G58), .C2(G232), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G1), .B2(G20), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR3_X1   g0019(.A1(new_n218), .A2(new_n219), .A3(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT0), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n219), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n221), .A2(new_n222), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n223), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n217), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n208), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(G200), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n218), .B1(G41), .B2(G45), .ZN(new_n255));
  AND2_X1   g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT67), .B1(new_n256), .B2(new_n227), .ZN(new_n257));
  AND2_X1   g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI211_X1 g0061(.A(new_n254), .B(new_n255), .C1(new_n257), .C2(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G222), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n267), .B1(new_n247), .B2(new_n265), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n256), .A2(new_n227), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n262), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n257), .B2(new_n261), .ZN(new_n276));
  XOR2_X1   g0076(.A(KEYINPUT68), .B(G226), .Z(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n253), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n272), .A2(new_n278), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n279), .B1(G190), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n218), .A2(G13), .A3(G20), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  XOR2_X1   g0083(.A(KEYINPUT8), .B(G58), .Z(new_n284));
  INV_X1    g0084(.A(KEYINPUT69), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G20), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n219), .A2(KEYINPUT69), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT70), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n203), .A2(G20), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n294), .B1(new_n284), .B2(new_n289), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n295), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n227), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n283), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n218), .B2(G20), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G50), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n304), .B1(new_n303), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n281), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(KEYINPUT72), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n303), .A2(new_n306), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT9), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n310), .A2(KEYINPUT72), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n310), .A2(KEYINPUT72), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n315), .A2(new_n317), .A3(new_n319), .A4(new_n281), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n311), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n265), .A2(G226), .A3(new_n266), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n265), .A2(G232), .A3(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G97), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n322), .B(new_n323), .C1(new_n286), .C2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n262), .B1(new_n325), .B2(new_n271), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n276), .A2(G238), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n327), .B1(new_n326), .B2(new_n328), .ZN(new_n331));
  OAI21_X1  g0131(.A(G200), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n326), .A2(new_n328), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT13), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(G190), .A3(new_n329), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n289), .A2(G77), .B1(G50), .B2(new_n291), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n219), .B2(G68), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n302), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT11), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(KEYINPUT11), .A3(new_n302), .ZN(new_n341));
  INV_X1    g0141(.A(new_n282), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n212), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT12), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n305), .A2(G68), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT73), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n340), .A2(new_n341), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n332), .A2(new_n335), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n332), .A2(new_n335), .A3(KEYINPUT74), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n280), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n312), .C1(G179), .C2(new_n355), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n359));
  INV_X1    g0159(.A(G107), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n359), .B1(new_n360), .B2(new_n265), .C1(new_n268), .C2(new_n213), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n271), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n256), .A2(KEYINPUT67), .A3(new_n227), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n259), .B1(new_n258), .B2(new_n260), .ZN(new_n364));
  OAI211_X1 g0164(.A(G274), .B(new_n275), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n276), .A2(G244), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G190), .ZN(new_n369));
  XOR2_X1   g0169(.A(KEYINPUT15), .B(G87), .Z(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n371));
  INV_X1    g0171(.A(new_n284), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n292), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n302), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT71), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(KEYINPUT71), .A3(new_n302), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n376), .A2(new_n377), .B1(new_n247), .B2(new_n342), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n367), .A2(G200), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n305), .A2(G77), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n369), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n321), .A2(new_n354), .A3(new_n358), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G179), .ZN(new_n383));
  AND2_X1   g0183(.A1(KEYINPUT3), .A2(G33), .ZN(new_n384));
  NOR2_X1   g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  OAI211_X1 g0185(.A(G226), .B(G1698), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT75), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n265), .A2(KEYINPUT75), .A3(G226), .A4(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n265), .A2(G223), .A3(new_n266), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n388), .A2(new_n389), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n271), .ZN(new_n393));
  OAI211_X1 g0193(.A(G232), .B(new_n255), .C1(new_n363), .C2(new_n364), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n365), .A2(new_n394), .A3(KEYINPUT76), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT76), .B1(new_n365), .B2(new_n394), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n383), .B(new_n393), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT77), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n236), .B(new_n275), .C1(new_n257), .C2(new_n261), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n262), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n365), .A2(new_n394), .A3(KEYINPUT76), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n404), .A2(KEYINPUT77), .A3(new_n383), .A4(new_n393), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n393), .A2(new_n365), .A3(new_n394), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n356), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT78), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT78), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n399), .A2(new_n405), .A3(new_n410), .A4(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n384), .A2(new_n385), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT7), .B1(new_n413), .B2(new_n219), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n384), .A2(new_n385), .A3(new_n415), .A4(G20), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G159), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n292), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G58), .A2(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n219), .B1(new_n224), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT16), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n263), .A2(new_n219), .A3(new_n264), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n415), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n413), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n422), .B1(new_n430), .B2(G68), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT16), .A3(new_n420), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n426), .A2(new_n432), .A3(new_n302), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n305), .A2(new_n284), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n372), .A2(new_n342), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n412), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT79), .B(KEYINPUT18), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n434), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT16), .B1(new_n431), .B2(new_n420), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n212), .B1(new_n428), .B2(new_n429), .ZN(new_n442));
  NOR4_X1   g0242(.A1(new_n442), .A2(new_n425), .A3(new_n419), .A4(new_n422), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n444), .B2(new_n302), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT17), .ZN(new_n446));
  INV_X1    g0246(.A(G190), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n404), .A2(new_n447), .A3(new_n393), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n406), .A2(new_n253), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n445), .A2(new_n446), .A3(new_n450), .A4(new_n435), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n402), .A2(new_n403), .B1(new_n271), .B2(new_n392), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(new_n447), .B1(new_n406), .B2(new_n253), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT17), .B1(new_n436), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n409), .B2(new_n411), .ZN(new_n457));
  INV_X1    g0257(.A(new_n438), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n439), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT14), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n334), .A2(new_n329), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(G169), .ZN(new_n463));
  AOI211_X1 g0263(.A(KEYINPUT14), .B(new_n356), .C1(new_n334), .C2(new_n329), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(new_n383), .ZN(new_n465));
  OR3_X1    g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n347), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n378), .A2(new_n380), .B1(new_n383), .B2(new_n368), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n367), .A2(new_n356), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n382), .A2(new_n460), .A3(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(new_n266), .C1(new_n384), .C2(new_n385), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT83), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n265), .A2(KEYINPUT83), .A3(G257), .A4(new_n266), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n413), .A2(G303), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n265), .A2(G264), .A3(G1698), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n475), .A2(new_n476), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n271), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n274), .A2(G1), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n257), .A2(new_n261), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n254), .B1(new_n257), .B2(new_n261), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n482), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(G270), .A2(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G283), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n219), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT80), .B(G97), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n286), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n207), .A2(G20), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n302), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n491), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n324), .A2(KEYINPUT80), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT80), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n497), .B1(new_n501), .B2(G33), .ZN(new_n502));
  INV_X1    g0302(.A(new_n495), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT20), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n282), .A2(G116), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n301), .A2(new_n227), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n218), .A2(G33), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(new_n282), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n207), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n488), .A2(new_n513), .A3(G169), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n506), .B(new_n511), .C1(new_n496), .C2(new_n504), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n480), .A2(G190), .A3(new_n487), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n484), .A2(new_n486), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n485), .B(G270), .C1(new_n364), .C2(new_n363), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n271), .B2(new_n479), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n517), .B(new_n518), .C1(new_n522), .C2(new_n253), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(G179), .A3(new_n513), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n488), .A2(new_n513), .A3(KEYINPUT21), .A4(G169), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n516), .A2(new_n523), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n219), .A2(G33), .A3(G116), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n219), .A2(KEYINPUT23), .A3(G107), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT23), .B1(new_n219), .B2(G107), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(KEYINPUT84), .B(KEYINPUT23), .C1(new_n219), .C2(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n219), .B(G87), .C1(new_n384), .C2(new_n385), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n534), .A2(KEYINPUT22), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n534), .A2(KEYINPUT22), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n527), .B(new_n533), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT24), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n534), .B(KEYINPUT22), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(new_n527), .A4(new_n533), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n302), .ZN(new_n543));
  INV_X1    g0343(.A(new_n510), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT25), .B1(new_n342), .B2(new_n360), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n342), .A2(KEYINPUT25), .A3(new_n360), .ZN(new_n547));
  AOI22_X1  g0347(.A1(G107), .A2(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(KEYINPUT85), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT85), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n508), .B1(new_n538), .B2(new_n541), .ZN(new_n551));
  INV_X1    g0351(.A(new_n548), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(G257), .B(G1698), .C1(new_n384), .C2(new_n385), .ZN(new_n555));
  OAI211_X1 g0355(.A(G250), .B(new_n266), .C1(new_n384), .C2(new_n385), .ZN(new_n556));
  INV_X1    g0356(.A(G294), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n555), .B(new_n556), .C1(new_n286), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n271), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n483), .A2(G264), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n519), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G169), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n383), .B2(new_n561), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n526), .B1(new_n554), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n253), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n558), .A2(new_n271), .B1(new_n483), .B2(G264), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n447), .A3(new_n519), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n543), .A2(new_n548), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n282), .A2(G97), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n510), .A2(new_n324), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n360), .B1(new_n428), .B2(new_n429), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n360), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT6), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n324), .A2(new_n360), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G97), .A2(G107), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n219), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n292), .A2(new_n247), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n574), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n571), .B(new_n573), .C1(new_n582), .C2(new_n508), .ZN(new_n583));
  OAI211_X1 g0383(.A(G244), .B(new_n266), .C1(new_n384), .C2(new_n385), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT4), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .A4(new_n266), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n490), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n271), .ZN(new_n590));
  AOI22_X1  g0390(.A1(G257), .A2(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n356), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n383), .A3(new_n591), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n583), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n370), .A2(new_n282), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  INV_X1    g0397(.A(new_n289), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(new_n501), .ZN(new_n599));
  INV_X1    g0399(.A(G87), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n501), .A2(new_n600), .A3(new_n360), .ZN(new_n601));
  NAND3_X1  g0401(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n219), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n265), .A2(new_n219), .A3(G68), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n596), .B1(new_n606), .B2(new_n302), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n544), .A2(new_n370), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(G244), .B(G1698), .C1(new_n384), .C2(new_n385), .ZN(new_n610));
  OAI211_X1 g0410(.A(G238), .B(new_n266), .C1(new_n384), .C2(new_n385), .ZN(new_n611));
  NAND2_X1  g0411(.A1(G33), .A2(G116), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT82), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT82), .A4(new_n612), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n271), .A3(new_n616), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n259), .A2(new_n274), .A3(new_n254), .A4(G1), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n482), .B1(new_n257), .B2(new_n261), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(G250), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n356), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n383), .A3(new_n620), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n609), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n510), .A2(new_n600), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n596), .B(new_n625), .C1(new_n606), .C2(new_n302), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(G200), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n617), .A2(G190), .A3(new_n620), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n569), .A2(new_n595), .A3(new_n624), .A4(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT81), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n592), .B2(new_n447), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n590), .A2(KEYINPUT81), .A3(new_n591), .A4(G190), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n592), .A2(G200), .ZN(new_n635));
  INV_X1    g0435(.A(new_n583), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n472), .A2(new_n564), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g0439(.A(new_n639), .B(KEYINPUT86), .Z(G372));
  INV_X1    g0440(.A(KEYINPUT18), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n456), .A2(new_n408), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n399), .A2(new_n405), .A3(new_n407), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT18), .B1(new_n643), .B2(new_n436), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n332), .A2(new_n335), .A3(new_n348), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n455), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n471), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n311), .A2(new_n320), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n358), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT87), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n638), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT87), .B1(new_n630), .B2(new_n637), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n516), .A2(new_n524), .A3(new_n525), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n563), .B1(new_n551), .B2(new_n552), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n653), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n624), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n624), .A2(new_n629), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n595), .ZN(new_n663));
  INV_X1    g0463(.A(new_n595), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n664), .A2(KEYINPUT26), .A3(new_n624), .A4(new_n629), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n660), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n472), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n651), .A2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n218), .A2(new_n219), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n517), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n655), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n526), .B2(new_n677), .ZN(new_n679));
  XOR2_X1   g0479(.A(KEYINPUT88), .B(G330), .Z(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT89), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n554), .A2(new_n675), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT85), .B1(new_n543), .B2(new_n548), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n551), .A2(new_n550), .A3(new_n552), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n563), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n683), .A2(new_n686), .A3(new_n569), .ZN(new_n687));
  INV_X1    g0487(.A(new_n686), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n675), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n656), .A2(new_n675), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n657), .A2(new_n675), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(KEYINPUT90), .A3(new_n694), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n691), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n220), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR4_X1   g0503(.A1(new_n492), .A2(G87), .A3(G107), .A4(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n225), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n686), .A2(new_n656), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n638), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n666), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n676), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n667), .A2(new_n676), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(KEYINPUT29), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n592), .A2(new_n561), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n522), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n590), .A2(new_n591), .B1(new_n566), .B2(new_n519), .ZN(new_n719));
  AOI21_X1  g0519(.A(G179), .B1(new_n719), .B2(KEYINPUT91), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n718), .A2(new_n720), .A3(new_n621), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n617), .A2(new_n590), .A3(new_n591), .A4(new_n620), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n480), .A2(new_n566), .A3(new_n487), .A4(G179), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT30), .B1(new_n722), .B2(new_n724), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n715), .B(new_n676), .C1(new_n721), .C2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n638), .A2(new_n564), .A3(new_n676), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT31), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT92), .B1(new_n721), .B2(new_n729), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n721), .A2(new_n729), .A3(KEYINPUT92), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n675), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n730), .B1(new_n732), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n680), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n714), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n707), .B1(new_n741), .B2(G1), .ZN(G364));
  NAND2_X1  g0542(.A1(new_n219), .A2(G13), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT93), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G45), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G1), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n702), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G303), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n219), .A2(new_n447), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n253), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n383), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G322), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n749), .A2(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G190), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT33), .B(G317), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n265), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n757), .A2(new_n447), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G326), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n219), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n751), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n760), .B(new_n762), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n764), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n756), .B(new_n766), .C1(G329), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n219), .B1(new_n768), .B2(G190), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT98), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT98), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n764), .A2(new_n753), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n771), .B1(new_n557), .B2(new_n775), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT99), .Z(new_n779));
  INV_X1    g0579(.A(new_n754), .ZN(new_n780));
  INV_X1    g0580(.A(new_n777), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G58), .A2(new_n780), .B1(new_n781), .B2(G77), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n782), .B1(new_n600), .B2(new_n752), .C1(new_n360), .C2(new_n765), .ZN(new_n783));
  INV_X1    g0583(.A(new_n758), .ZN(new_n784));
  INV_X1    g0584(.A(new_n761), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n212), .B1(new_n785), .B2(new_n202), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n783), .A2(new_n413), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n324), .B2(new_n775), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n769), .A2(new_n418), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n779), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n227), .B1(G20), .B2(new_n356), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n748), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT95), .Z(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n794), .B1(new_n679), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n798), .A2(new_n793), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n701), .A2(new_n265), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n226), .A2(new_n274), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n248), .C2(new_n274), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n701), .A2(new_n413), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G355), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n804), .B(new_n806), .C1(G116), .C2(new_n220), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n800), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT100), .Z(new_n809));
  OAI211_X1 g0609(.A(new_n682), .B(new_n748), .C1(new_n680), .C2(new_n679), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT94), .Z(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(G396));
  NOR2_X1   g0612(.A1(new_n470), .A2(new_n675), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n378), .A2(new_n380), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n675), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(new_n381), .B1(new_n468), .B2(new_n469), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n713), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n675), .B1(new_n659), .B2(new_n666), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n817), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(new_n739), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n748), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n600), .A2(new_n765), .B1(new_n777), .B2(new_n207), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n265), .B1(new_n758), .B2(G283), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n826), .B1(new_n360), .B2(new_n752), .C1(new_n749), .C2(new_n785), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n825), .B(new_n827), .C1(G311), .C2(new_n770), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n828), .B1(new_n324), .B2(new_n775), .C1(new_n557), .C2(new_n754), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n781), .A2(G159), .B1(G137), .B2(new_n761), .ZN(new_n830));
  INV_X1    g0630(.A(G143), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n831), .B2(new_n754), .C1(new_n293), .C2(new_n784), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n752), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n770), .A2(G132), .B1(G50), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(new_n212), .C2(new_n765), .ZN(new_n837));
  INV_X1    g0637(.A(G58), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n265), .B1(new_n832), .B2(new_n833), .C1(new_n775), .C2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n829), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n793), .A2(new_n795), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n840), .A2(new_n793), .B1(new_n247), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n842), .B(new_n747), .C1(new_n817), .C2(new_n797), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n824), .A2(new_n843), .ZN(G384));
  NAND2_X1  g0644(.A1(new_n347), .A2(new_n675), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n466), .B2(new_n353), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n349), .B(new_n845), .C1(new_n848), .C2(new_n348), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n721), .A2(new_n729), .A3(KEYINPUT92), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n733), .ZN(new_n852));
  AOI22_X1  g0652(.A1(KEYINPUT31), .A2(new_n731), .B1(new_n852), .B2(new_n675), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n736), .A2(new_n715), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n817), .B(new_n850), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  INV_X1    g0656(.A(new_n673), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n436), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n457), .B(new_n438), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n859), .B2(new_n455), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n436), .A2(new_n857), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n436), .A2(new_n453), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT102), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n457), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT37), .B1(new_n457), .B2(new_n864), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n643), .A2(new_n436), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n866), .A2(new_n867), .B1(KEYINPUT37), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n856), .B1(new_n860), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n460), .A2(new_n861), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n412), .A2(new_n864), .A3(new_n436), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n873), .B1(new_n876), .B2(new_n865), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n855), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT105), .ZN(new_n880));
  OR3_X1    g0680(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT40), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n879), .B2(KEYINPUT40), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT103), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n455), .B1(new_n642), .B2(new_n644), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT104), .B1(new_n886), .B2(new_n861), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n643), .A2(KEYINPUT18), .A3(new_n436), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n641), .B1(new_n456), .B2(new_n408), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(new_n889), .B1(new_n454), .B2(new_n451), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n890), .A2(new_n891), .A3(new_n858), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n873), .B(KEYINPUT103), .C1(new_n876), .C2(new_n865), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n885), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n883), .B1(new_n856), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n855), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n881), .A2(new_n882), .B1(new_n897), .B2(KEYINPUT40), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n853), .A2(new_n854), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n311), .A2(new_n320), .A3(new_n358), .A4(new_n381), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n353), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n466), .A2(new_n347), .B1(new_n469), .B2(new_n468), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n901), .A2(new_n455), .A3(new_n859), .A4(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n898), .B(new_n904), .Z(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n680), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n467), .A2(new_n675), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n895), .A2(new_n856), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n910), .A3(new_n878), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n871), .A2(new_n878), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT39), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n813), .B1(new_n820), .B2(new_n817), .ZN(new_n915));
  INV_X1    g0715(.A(new_n850), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n912), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n645), .A2(new_n673), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n650), .B1(new_n714), .B2(new_n472), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n906), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n218), .B2(new_n744), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n575), .A2(new_n579), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n207), .B1(new_n927), .B2(KEYINPUT35), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n928), .B(new_n228), .C1(KEYINPUT35), .C2(new_n927), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT101), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT36), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n421), .A2(G77), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n225), .A2(new_n932), .B1(G50), .B2(new_n212), .ZN(new_n933));
  INV_X1    g0733(.A(G13), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(G1), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n926), .A2(new_n931), .A3(new_n935), .ZN(G367));
  AOI21_X1  g0736(.A(new_n664), .B1(new_n583), .B2(new_n675), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n937), .A2(new_n938), .B1(new_n664), .B2(new_n675), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n693), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT42), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(KEYINPUT107), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n664), .B1(new_n942), .B2(new_n688), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n941), .B1(new_n675), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT108), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT108), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n941), .B(new_n946), .C1(new_n675), .C2(new_n943), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n626), .A2(new_n676), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n624), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(new_n624), .A3(new_n629), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT106), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n949), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT43), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n945), .A2(new_n947), .A3(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n945), .A2(new_n947), .B1(new_n954), .B2(new_n953), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT109), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n690), .A2(new_n942), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n956), .A2(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n958), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n958), .B(new_n959), .C1(new_n956), .C2(new_n957), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n702), .B(KEYINPUT41), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n939), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n699), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT45), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n699), .A2(new_n966), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n690), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(new_n691), .A3(new_n970), .ZN(new_n973));
  INV_X1    g0773(.A(new_n689), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n693), .B1(new_n974), .B2(new_n692), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n682), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n740), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n972), .A2(new_n973), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n965), .B1(new_n978), .B2(new_n741), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n962), .B(new_n963), .C1(new_n979), .C2(new_n746), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n835), .A2(KEYINPUT46), .A3(G116), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n784), .B2(new_n557), .C1(new_n776), .C2(new_n785), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT46), .B1(new_n835), .B2(G116), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n983), .A2(KEYINPUT110), .B1(new_n769), .B2(new_n986), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n413), .B1(new_n765), .B2(new_n501), .C1(new_n763), .C2(new_n777), .ZN(new_n988));
  NOR4_X1   g0788(.A1(new_n982), .A2(new_n985), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n360), .B2(new_n775), .C1(new_n749), .C2(new_n754), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n265), .B1(new_n785), .B2(new_n831), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G159), .B2(new_n758), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n838), .B2(new_n752), .C1(new_n247), .C2(new_n765), .ZN(new_n993));
  INV_X1    g0793(.A(new_n775), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(G68), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G150), .A2(new_n780), .B1(new_n781), .B2(G50), .ZN(new_n996));
  INV_X1    g0796(.A(G137), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n995), .B(new_n996), .C1(new_n997), .C2(new_n769), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n990), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT47), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n793), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n243), .A2(new_n802), .B1(new_n701), .B2(new_n370), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n801), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n953), .A2(new_n798), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1001), .A2(new_n747), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n980), .A2(new_n1005), .ZN(G387));
  INV_X1    g0806(.A(new_n977), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n703), .B1(new_n976), .B2(new_n740), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n793), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n781), .A2(G303), .B1(G322), .B2(new_n761), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n776), .B2(new_n784), .C1(new_n986), .C2(new_n754), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT48), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n763), .B2(new_n775), .C1(new_n557), .C2(new_n752), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT49), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n265), .B1(new_n770), .B2(G326), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n207), .C2(new_n765), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n265), .B1(new_n785), .B2(new_n418), .C1(new_n372), .C2(new_n784), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n752), .A2(new_n247), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G50), .B2(new_n780), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n293), .B2(new_n769), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1018), .B(new_n1021), .C1(G68), .C2(new_n781), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n994), .A2(new_n370), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n324), .C2(new_n765), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1010), .B1(new_n1017), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n239), .A2(G45), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n704), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1026), .A2(new_n802), .B1(new_n1027), .B2(new_n805), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n284), .A2(new_n202), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT111), .Z(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT50), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n704), .B(new_n274), .C1(new_n212), .C2(new_n247), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1028), .A2(new_n1033), .B1(G107), .B2(new_n220), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1025), .B1(new_n801), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n747), .C1(new_n974), .C2(new_n799), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n746), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1009), .B(new_n1036), .C1(new_n1037), .C2(new_n976), .ZN(G393));
  NAND2_X1  g0838(.A1(new_n972), .A2(new_n973), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n703), .B1(new_n1039), .B2(new_n1007), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n978), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n972), .A2(new_n746), .A3(new_n973), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT114), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n780), .A2(G159), .B1(G150), .B2(new_n761), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n265), .B1(new_n212), .B2(new_n752), .C1(new_n1044), .C2(KEYINPUT51), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n994), .A2(G77), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n202), .B2(new_n784), .C1(new_n372), .C2(new_n777), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT113), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n769), .A2(new_n831), .B1(new_n600), .B2(new_n765), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1044), .B2(KEYINPUT51), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1049), .B(new_n1051), .C1(new_n1048), .C2(new_n1047), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n765), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n265), .B1(new_n1053), .B2(G107), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n763), .B2(new_n752), .C1(new_n784), .C2(new_n749), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n785), .A2(new_n986), .B1(new_n754), .B2(new_n776), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  AOI211_X1 g0857(.A(new_n1055), .B(new_n1057), .C1(G322), .C2(new_n770), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n207), .B2(new_n775), .C1(new_n557), .C2(new_n777), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1052), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n748), .B1(new_n1060), .B2(new_n793), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n251), .A2(new_n802), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n801), .B(new_n1062), .C1(new_n220), .C2(new_n501), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT112), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1061), .B(new_n1064), .C1(new_n942), .C2(new_n799), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1042), .A2(new_n1043), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1043), .B1(new_n1042), .B2(new_n1065), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1041), .B1(new_n1067), .B2(new_n1068), .ZN(G390));
  OAI21_X1  g0869(.A(new_n908), .B1(new_n915), .B2(new_n916), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n911), .A2(new_n913), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n909), .A2(new_n878), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n675), .B(new_n816), .C1(new_n709), .C2(new_n666), .ZN(new_n1073));
  OAI21_X1  g0873(.A(KEYINPUT115), .B1(new_n1073), .B2(new_n813), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n816), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n710), .A2(new_n676), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT115), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n813), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1074), .A2(new_n850), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1072), .A2(new_n1080), .A3(new_n908), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n732), .A2(new_n736), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n730), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1084), .A2(new_n680), .A3(new_n817), .A4(new_n850), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n1071), .A2(new_n1081), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT116), .ZN(new_n1088));
  INV_X1    g0888(.A(G330), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n855), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n852), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n818), .B1(new_n1082), .B2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1092), .A2(KEYINPUT116), .A3(G330), .A4(new_n850), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1071), .B2(new_n1081), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1087), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT117), .B1(new_n904), .B2(G330), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT117), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n899), .A2(new_n903), .A3(new_n1098), .A4(new_n1089), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n922), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1073), .A2(KEYINPUT115), .A3(new_n813), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1077), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n680), .B(new_n817), .C1(new_n853), .C2(new_n730), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1101), .A2(new_n1102), .B1(new_n1103), .B2(new_n916), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n850), .B1(new_n1092), .B2(G330), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT118), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1107));
  OAI211_X1 g0907(.A(G330), .B(new_n817), .C1(new_n853), .C2(new_n854), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n916), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT118), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1085), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1103), .A2(new_n916), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1090), .A2(new_n1093), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n915), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1100), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1096), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n702), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n746), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n910), .B1(new_n871), .B2(new_n878), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n896), .B2(new_n910), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n796), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n265), .B1(new_n765), .B2(new_n202), .C1(new_n777), .C2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n752), .A2(new_n293), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT53), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1128), .A2(new_n1129), .B1(G137), .B2(new_n758), .ZN(new_n1130));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1130), .B1(new_n1129), .B2(new_n1128), .C1(new_n1131), .C2(new_n785), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1127), .B(new_n1132), .C1(G125), .C2(new_n770), .ZN(new_n1133));
  INV_X1    g0933(.A(G132), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n754), .C1(new_n418), .C2(new_n775), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n501), .A2(new_n777), .B1(new_n765), .B2(new_n212), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n265), .B1(new_n761), .B2(G283), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n600), .B2(new_n752), .C1(new_n360), .C2(new_n784), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1136), .B(new_n1138), .C1(G294), .C2(new_n770), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1046), .B(new_n1139), .C1(new_n207), .C2(new_n754), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1010), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n372), .B2(new_n841), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1125), .A2(new_n747), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1122), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1121), .A2(new_n1144), .ZN(G378));
  INV_X1    g0945(.A(new_n358), .ZN(new_n1146));
  OR3_X1    g0946(.A1(new_n649), .A2(KEYINPUT120), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT120), .B1(new_n649), .B2(new_n1146), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n312), .A3(new_n857), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n312), .A2(new_n857), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1150), .A2(new_n1154), .A3(new_n1152), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n914), .B2(new_n920), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n917), .A2(new_n912), .B1(new_n645), .B2(new_n673), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(new_n1158), .C1(new_n1124), .C2(new_n908), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n881), .A2(new_n882), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n897), .A2(KEYINPUT40), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(G330), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n898), .A2(new_n1160), .A3(G330), .A4(new_n1162), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1100), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1167), .A2(new_n1168), .B1(new_n1120), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n702), .B1(new_n1170), .B2(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1120), .A2(new_n1169), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1172), .A2(KEYINPUT57), .A3(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT121), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1159), .A2(new_n796), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n841), .A2(new_n202), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n784), .A2(new_n1134), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n754), .A2(new_n1131), .B1(new_n777), .B2(new_n997), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G125), .C2(new_n761), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n752), .B2(new_n1126), .C1(new_n775), .C2(new_n293), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT59), .Z(new_n1183));
  AOI21_X1  g0983(.A(G41), .B1(new_n770), .B2(G124), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G33), .B1(new_n1053), .B2(G159), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n781), .A2(new_n370), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G107), .A2(new_n780), .B1(new_n1053), .B2(G58), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n763), .B2(new_n769), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n413), .B1(new_n784), .B2(new_n324), .C1(new_n207), .C2(new_n785), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1189), .A2(G41), .A3(new_n1190), .A4(new_n1019), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n995), .A2(new_n1187), .A3(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n202), .B1(new_n384), .B2(G41), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1186), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n748), .B1(new_n1196), .B2(new_n793), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1177), .A2(new_n1178), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1172), .B2(new_n746), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1175), .A2(new_n1176), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1176), .B1(new_n1175), .B2(new_n1200), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1202), .A2(new_n1203), .ZN(G375));
  NOR3_X1   g1004(.A1(new_n737), .A2(new_n738), .A3(new_n818), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1205), .A2(new_n850), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1110), .B1(new_n1206), .B2(new_n1109), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1111), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1116), .B(new_n1100), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1118), .A2(new_n964), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1037), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n916), .A2(new_n795), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n752), .A2(new_n418), .B1(new_n777), .B2(new_n293), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1053), .A2(G58), .B1(G132), .B2(new_n761), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1214), .B(new_n265), .C1(new_n784), .C2(new_n1126), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(G128), .C2(new_n770), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n202), .B2(new_n775), .C1(new_n997), .C2(new_n754), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n754), .A2(new_n763), .B1(new_n777), .B2(new_n360), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n265), .B1(new_n758), .B2(G116), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n247), .B2(new_n765), .C1(new_n557), .C2(new_n785), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(G303), .C2(new_n770), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1023), .B(new_n1221), .C1(new_n324), .C2(new_n752), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1010), .B1(new_n1217), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n212), .B2(new_n841), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1212), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1211), .B1(new_n747), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1210), .A2(new_n1226), .ZN(G381));
  NOR2_X1   g1027(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1228));
  INV_X1    g1028(.A(G378), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  OR3_X1    g1030(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1042), .A2(new_n1065), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT114), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1233), .A2(new_n1066), .B1(new_n1040), .B2(new_n978), .ZN(new_n1234));
  INV_X1    g1034(.A(G384), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1005), .A4(new_n980), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1230), .A2(new_n1231), .A3(new_n1236), .ZN(G407));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G343), .C2(new_n1230), .ZN(G409));
  OAI211_X1 g1038(.A(G378), .B(new_n1200), .C1(new_n1171), .C2(new_n1174), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1170), .A2(new_n964), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1172), .A2(new_n746), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1198), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1229), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT122), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1209), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1117), .B1(new_n1246), .B2(KEYINPUT60), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n703), .B1(new_n1209), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1245), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1112), .A2(KEYINPUT60), .A3(new_n1116), .A4(new_n1100), .ZN(new_n1251));
  AND4_X1   g1051(.A1(new_n1245), .A2(new_n1249), .A3(new_n1118), .A4(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1226), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1235), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G384), .B(new_n1226), .C1(new_n1250), .C2(new_n1252), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n674), .A2(G213), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1244), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1258), .A2(KEYINPUT62), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1244), .A2(new_n1257), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT124), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n674), .A2(G213), .A3(G2897), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1254), .A2(new_n1264), .A3(new_n1255), .A4(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1254), .A2(new_n1264), .A3(new_n1255), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1261), .A2(new_n1263), .A3(new_n1266), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1258), .A2(KEYINPUT62), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1259), .A2(new_n1260), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n962), .A2(new_n963), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n978), .A2(new_n741), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n964), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1275), .B2(new_n1037), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1005), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1234), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G390), .A2(new_n980), .A3(new_n1005), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  XOR2_X1   g1080(.A(G393), .B(G396), .Z(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1278), .A2(new_n1279), .A3(new_n1281), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1272), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT125), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1244), .A2(new_n1256), .A3(KEYINPUT63), .A4(new_n1257), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1278), .A2(new_n1279), .A3(new_n1281), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1281), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1270), .A2(new_n1260), .A3(new_n1288), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT123), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1258), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1294), .B1(new_n1258), .B2(new_n1295), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1287), .B1(new_n1293), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1258), .A2(new_n1295), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT123), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1296), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1303), .A2(new_n1292), .A3(KEYINPUT125), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1286), .B1(new_n1300), .B2(new_n1304), .ZN(G405));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G375), .A2(new_n1306), .A3(new_n1229), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT126), .B1(new_n1228), .B2(G378), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1239), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1256), .A2(KEYINPUT127), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1256), .A2(KEYINPUT127), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1285), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1285), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1309), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1312), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1315), .A2(new_n1239), .A3(new_n1308), .A4(new_n1307), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(G402));
endmodule


