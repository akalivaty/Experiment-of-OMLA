//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  XOR2_X1   g000(.A(KEYINPUT73), .B(G217), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G902), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT24), .B(G110), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(G128), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n194), .B(new_n198), .C1(new_n199), .C2(KEYINPUT23), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n197), .B1(new_n200), .B2(G110), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  XOR2_X1   g018(.A(G125), .B(G140), .Z(new_n205));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n206));
  OAI211_X1 g020(.A(G146), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n201), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT75), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n211), .B(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n209), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  INV_X1    g030(.A(G110), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT74), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n217), .B1(new_n200), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n218), .B2(new_n200), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n216), .B(new_n220), .C1(new_n195), .C2(new_n196), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n213), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT22), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT22), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n230), .A3(new_n227), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n229), .A2(new_n231), .A3(G137), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n213), .A2(new_n221), .A3(new_n235), .A4(new_n234), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n190), .B1(new_n240), .B2(KEYINPUT25), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(KEYINPUT25), .B2(new_n240), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n239), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n190), .A2(new_n238), .ZN(new_n245));
  XOR2_X1   g059(.A(new_n245), .B(KEYINPUT77), .Z(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XOR2_X1   g066(.A(new_n252), .B(KEYINPUT27), .Z(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT26), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(G101), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n209), .A2(G143), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n191), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G146), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n209), .A2(KEYINPUT64), .A3(G143), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n265), .A2(new_n266), .B1(new_n264), .B2(G146), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n264), .A2(KEYINPUT65), .A3(G146), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT65), .B1(new_n264), .B2(G146), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n261), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G128), .ZN(new_n272));
  OAI22_X1  g086(.A1(new_n262), .A2(new_n267), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n233), .A2(G134), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(G137), .ZN(new_n279));
  AND2_X1   g093(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G131), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(G137), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n277), .A2(new_n281), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n275), .A2(new_n283), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G131), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n273), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT11), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n280), .B1(new_n279), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n283), .B1(new_n275), .B2(new_n274), .ZN(new_n292));
  OAI21_X1  g106(.A(G131), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n284), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n209), .A2(KEYINPUT64), .A3(G143), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT64), .B1(new_n209), .B2(G143), .ZN(new_n296));
  OAI22_X1  g110(.A1(new_n295), .A2(new_n296), .B1(G143), .B2(new_n209), .ZN(new_n297));
  AND2_X1   g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  NOR2_X1   g112(.A1(KEYINPUT0), .A2(G128), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n264), .A2(G146), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n209), .B2(G143), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n264), .A2(KEYINPUT65), .A3(G146), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n297), .A2(new_n300), .B1(new_n305), .B2(new_n298), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n294), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n287), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT2), .B(G113), .Z(new_n309));
  XNOR2_X1  g123(.A(G116), .B(G119), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT70), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n310), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT2), .B(G113), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(KEYINPUT70), .A3(new_n313), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n308), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n308), .A2(KEYINPUT28), .A3(new_n318), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n284), .A2(new_n286), .ZN(new_n324));
  OAI21_X1  g138(.A(G128), .B1(new_n271), .B2(new_n301), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n297), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n305), .A2(G128), .A3(new_n271), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n307), .A2(KEYINPUT67), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n294), .A2(new_n330), .A3(new_n306), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(new_n318), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n255), .B1(new_n323), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT69), .B1(new_n332), .B2(KEYINPUT30), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n294), .A2(new_n330), .A3(new_n306), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n330), .B1(new_n294), .B2(new_n306), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n287), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT69), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT30), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n308), .A2(KEYINPUT30), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n335), .A2(new_n317), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT31), .ZN(new_n344));
  INV_X1    g158(.A(new_n319), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n255), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n344), .B1(new_n343), .B2(new_n346), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n334), .B(new_n347), .C1(new_n348), .C2(KEYINPUT71), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n350));
  AOI211_X1 g164(.A(new_n350), .B(new_n344), .C1(new_n343), .C2(new_n346), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n250), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n346), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT31), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n350), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n347), .A2(new_n334), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n348), .A2(KEYINPUT71), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT72), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(G472), .A2(G902), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n360), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(new_n362), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n308), .A2(new_n318), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n321), .A2(new_n322), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n255), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT29), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n345), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n343), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n368), .B1(new_n323), .B2(new_n333), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI221_X1 g187(.A(new_n238), .B1(new_n367), .B2(new_n369), .C1(new_n373), .C2(KEYINPUT29), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n359), .A2(new_n365), .B1(G472), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n249), .B1(new_n363), .B2(new_n375), .ZN(new_n376));
  NOR3_X1   g190(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G237), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n223), .A3(G214), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n264), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n282), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n382), .ZN(new_n386));
  AOI21_X1  g200(.A(G143), .B1(new_n251), .B2(G214), .ZN(new_n387));
  OAI21_X1  g201(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n381), .A2(KEYINPUT88), .A3(new_n282), .A4(new_n382), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n208), .A2(KEYINPUT19), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n208), .A2(KEYINPUT19), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n209), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n207), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n205), .A2(G146), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n210), .ZN(new_n396));
  NAND3_X1  g210(.A1(KEYINPUT87), .A2(KEYINPUT18), .A3(G131), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n386), .B2(new_n387), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n381), .A2(new_n382), .A3(new_n397), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G113), .B(G122), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n404), .B(G104), .Z(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(KEYINPUT17), .B(G131), .C1(new_n386), .C2(new_n387), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n215), .A2(new_n207), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT17), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n385), .A2(new_n410), .A3(new_n388), .A4(new_n389), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n405), .A3(new_n402), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n378), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n414), .B(new_n415), .ZN(new_n416));
  AOI211_X1 g230(.A(new_n406), .B(new_n401), .C1(new_n409), .C2(new_n411), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n405), .B1(new_n394), .B2(new_n402), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT89), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n407), .A2(new_n413), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT20), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G475), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n412), .A2(new_n402), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n406), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT91), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n413), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n405), .B1(new_n412), .B2(new_n402), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n431), .B2(KEYINPUT91), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n426), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT92), .B1(new_n425), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n436));
  AOI211_X1 g250(.A(new_n436), .B(new_n433), .C1(new_n416), .C2(new_n424), .ZN(new_n437));
  INV_X1    g251(.A(G122), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n438), .A2(G116), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(G116), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G107), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G128), .B(G143), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT13), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n264), .A2(G128), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n445), .B(G134), .C1(KEYINPUT13), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n278), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT14), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n440), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT93), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n439), .B1(new_n450), .B2(new_n440), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n442), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n444), .B(new_n278), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n441), .A2(new_n442), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n449), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT9), .B(G234), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n187), .A2(G953), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n449), .B(new_n460), .C1(new_n454), .C2(new_n457), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OR3_X1    g279(.A1(new_n458), .A2(new_n463), .A3(new_n461), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n238), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n467), .B(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n223), .A2(G952), .ZN(new_n471));
  NAND2_X1  g285(.A1(G234), .A2(G237), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(G902), .A3(G953), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT21), .B(G898), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR4_X1   g292(.A1(new_n435), .A2(new_n437), .A3(new_n470), .A4(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(KEYINPUT78), .A2(G104), .ZN(new_n480));
  NOR2_X1   g294(.A1(KEYINPUT78), .A2(G104), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n442), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT3), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT3), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n442), .A3(G104), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT79), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT79), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n487), .A2(new_n484), .A3(new_n442), .A4(G104), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G101), .ZN(new_n490));
  OR3_X1    g304(.A1(new_n480), .A2(new_n481), .A3(new_n442), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n483), .A2(new_n489), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n482), .B1(G104), .B2(new_n442), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G101), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT5), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n312), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n193), .A3(G116), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G113), .ZN(new_n499));
  OAI22_X1  g313(.A1(new_n497), .A2(new_n499), .B1(new_n313), .B2(new_n312), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n483), .A2(new_n491), .ZN(new_n503));
  INV_X1    g317(.A(new_n489), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n502), .B(G101), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n317), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n480), .A2(new_n481), .A3(new_n442), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(KEYINPUT3), .B2(new_n482), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n490), .B1(new_n509), .B2(new_n489), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n501), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G110), .B(G122), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n501), .B(new_n513), .C1(new_n506), .C2(new_n511), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(KEYINPUT6), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n297), .A2(new_n300), .ZN(new_n518));
  INV_X1    g332(.A(new_n298), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n518), .B1(new_n270), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G125), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n326), .A2(new_n327), .A3(new_n202), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G224), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(G953), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT85), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n523), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n512), .A2(new_n528), .A3(new_n514), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n517), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n513), .B(KEYINPUT8), .Z(new_n531));
  NAND2_X1  g345(.A1(new_n495), .A2(new_n500), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n501), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT7), .B1(new_n524), .B2(G953), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n523), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n534), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n521), .B2(new_n522), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(G902), .B1(new_n538), .B2(new_n516), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G210), .B1(G237), .B2(G902), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT86), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n542), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G214), .B1(G237), .B2(G902), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT84), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G221), .B1(new_n459), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G469), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(new_n238), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G140), .ZN(new_n553));
  INV_X1    g367(.A(G227), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(G953), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n553), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT80), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n505), .A2(new_n306), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n511), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n520), .B1(new_n510), .B2(new_n502), .ZN(new_n560));
  OAI21_X1  g374(.A(G101), .B1(new_n503), .B2(new_n504), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT4), .A3(new_n492), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(KEYINPUT80), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n294), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n273), .A2(new_n492), .A3(KEYINPUT10), .A4(new_n494), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT82), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT10), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n326), .B2(new_n327), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n570), .A2(KEYINPUT82), .A3(new_n492), .A4(new_n494), .ZN(new_n571));
  OAI21_X1  g385(.A(G128), .B1(new_n301), .B2(new_n256), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n270), .A2(KEYINPUT81), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT81), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n191), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n305), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n576), .A3(new_n327), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(new_n492), .A3(new_n494), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n568), .A2(new_n571), .B1(new_n569), .B2(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n564), .A2(new_n565), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n565), .B1(new_n564), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n556), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n577), .A2(new_n492), .A3(new_n494), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n273), .B1(new_n492), .B2(new_n494), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n294), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT12), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(KEYINPUT12), .B(new_n294), .C1(new_n583), .C2(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n511), .A2(new_n558), .A3(new_n557), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT80), .B1(new_n560), .B2(new_n562), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n579), .B(new_n565), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n556), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n582), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n552), .B1(new_n595), .B2(new_n551), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT83), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n593), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n581), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n593), .B1(new_n589), .B2(new_n592), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n589), .A2(new_n592), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n556), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n579), .B1(new_n590), .B2(new_n591), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n294), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n592), .A3(new_n593), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n606), .A3(KEYINPUT83), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n601), .A2(G469), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n550), .B1(new_n596), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n479), .A2(new_n548), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n376), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  AOI211_X1 g426(.A(new_n249), .B(new_n550), .C1(new_n596), .C2(new_n608), .ZN(new_n613));
  INV_X1    g427(.A(G472), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n352), .B2(new_n358), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n613), .B(new_n361), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT95), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n359), .A2(new_n238), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n620), .A2(KEYINPUT95), .A3(new_n361), .A4(new_n613), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n435), .A2(new_n437), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n478), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n467), .A2(new_n468), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n462), .A2(KEYINPUT33), .A3(new_n464), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n465), .A2(new_n466), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(KEYINPUT33), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n238), .A2(G478), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n540), .A2(new_n541), .ZN(new_n632));
  INV_X1    g446(.A(new_n541), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n530), .B2(new_n539), .ZN(new_n634));
  INV_X1    g448(.A(new_n546), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n624), .A2(new_n625), .A3(new_n631), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n622), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT96), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n638), .B(new_n640), .ZN(G6));
  XOR2_X1   g455(.A(new_n423), .B(KEYINPUT20), .Z(new_n642));
  NAND2_X1  g456(.A1(new_n470), .A2(new_n434), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n636), .A3(new_n625), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n622), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NOR2_X1   g463(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n222), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n247), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n242), .A2(new_n652), .ZN(new_n653));
  AND4_X1   g467(.A1(new_n479), .A2(new_n548), .A3(new_n609), .A4(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n364), .B1(new_n352), .B2(new_n358), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n619), .B2(G472), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AOI21_X1  g473(.A(KEYINPUT71), .B1(new_n353), .B2(KEYINPUT31), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n347), .A2(new_n334), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT72), .B1(new_n662), .B2(new_n357), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n349), .A2(new_n250), .A3(new_n351), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n365), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n374), .A2(G472), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n665), .B(new_n666), .C1(KEYINPUT32), .C2(new_n655), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n636), .A2(new_n653), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n474), .B1(new_n476), .B2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n642), .A2(new_n643), .A3(new_n670), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n668), .A2(new_n609), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT97), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT97), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n667), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XOR2_X1   g492(.A(new_n670), .B(KEYINPUT39), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n609), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT40), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n624), .A2(new_n470), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n545), .B(KEYINPUT38), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n242), .A2(new_n546), .A3(new_n652), .ZN(new_n685));
  NOR4_X1   g499(.A1(new_n681), .A2(new_n682), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(G902), .B1(new_n370), .B2(new_n366), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n255), .B1(new_n343), .B2(new_n319), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n665), .B(new_n690), .C1(KEYINPUT32), .C2(new_n655), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(KEYINPUT98), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(KEYINPUT98), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  INV_X1    g512(.A(new_n670), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n631), .B(new_n699), .C1(new_n435), .C2(new_n437), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n701), .A2(new_n609), .A3(new_n668), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n667), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  INV_X1    g518(.A(new_n249), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n582), .A2(new_n594), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n238), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n593), .B1(new_n605), .B2(new_n592), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n551), .B(new_n238), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n549), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n667), .A2(new_n637), .A3(new_n705), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT41), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G113), .ZN(G15));
  NAND4_X1  g530(.A1(new_n667), .A2(new_n705), .A3(new_n646), .A4(new_n713), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NAND4_X1  g532(.A1(new_n667), .A2(new_n479), .A3(new_n668), .A4(new_n713), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  INV_X1    g534(.A(new_n347), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n367), .A2(new_n255), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n354), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n721), .B1(new_n723), .B2(KEYINPUT100), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT100), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n354), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n364), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n619), .B2(G472), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n636), .B(new_n470), .C1(new_n435), .C2(new_n437), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n729), .A2(new_n478), .A3(new_n712), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(new_n730), .A3(new_n705), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND2_X1  g546(.A1(new_n724), .A2(new_n726), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n360), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n734), .B(new_n653), .C1(new_n615), .C2(new_n614), .ZN(new_n735));
  INV_X1    g549(.A(new_n636), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n712), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n701), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT101), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT101), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n700), .A2(new_n712), .A3(new_n736), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n728), .A2(new_n740), .A3(new_n653), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(new_n552), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n603), .A2(new_n606), .A3(G469), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n711), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n747), .A2(new_n748), .A3(new_n549), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n747), .B2(new_n549), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n543), .A2(new_n546), .A3(new_n544), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n667), .A2(new_n705), .A3(new_n752), .A4(new_n701), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n376), .A2(KEYINPUT42), .A3(new_n701), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT103), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT103), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n282), .ZN(G33));
  AND4_X1   g576(.A1(new_n667), .A2(new_n705), .A3(new_n752), .A4(new_n671), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n278), .ZN(G36));
  AOI21_X1  g578(.A(KEYINPUT45), .B1(new_n601), .B2(new_n607), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n599), .A2(new_n600), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n551), .B(new_n765), .C1(KEYINPUT45), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n552), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT104), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n768), .A2(KEYINPUT46), .B1(new_n551), .B2(new_n595), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n549), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n679), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n623), .A2(new_n631), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT43), .Z(new_n778));
  INV_X1    g592(.A(new_n656), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n653), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n751), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  NAND2_X1  g599(.A1(new_n774), .A2(KEYINPUT47), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n549), .C1(new_n771), .C2(new_n773), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n667), .A2(new_n705), .A3(new_n700), .A4(new_n751), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  INV_X1    g605(.A(new_n694), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n708), .A2(new_n711), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT49), .Z(new_n794));
  NAND3_X1  g608(.A1(new_n705), .A2(new_n547), .A3(new_n549), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n683), .A2(new_n777), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n728), .A2(new_n705), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n778), .A2(new_n474), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n778), .A2(KEYINPUT109), .A3(new_n474), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n751), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n786), .A2(new_n788), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT110), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n708), .A2(new_n550), .A3(new_n711), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n807), .A2(KEYINPUT110), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n712), .A2(new_n751), .A3(new_n249), .A4(new_n473), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n624), .A2(new_n631), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n792), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n802), .A2(new_n803), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n712), .A2(new_n751), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n683), .A2(new_n546), .A3(new_n712), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n804), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(KEYINPUT111), .ZN(new_n821));
  OAI221_X1 g635(.A(new_n815), .B1(new_n735), .B2(new_n818), .C1(new_n821), .C2(KEYINPUT50), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n821), .A2(KEYINPUT50), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n812), .B1(new_n824), .B2(KEYINPUT112), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n822), .A2(new_n826), .A3(new_n823), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n798), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n816), .A2(new_n376), .A3(new_n817), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT48), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n804), .A2(new_n737), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n792), .A2(new_n624), .A3(new_n631), .A4(new_n813), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n830), .A2(new_n471), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n807), .A2(new_n809), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(new_n806), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n833), .B1(new_n824), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n747), .A2(new_n549), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n242), .A2(new_n652), .A3(new_n699), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n729), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n667), .A2(new_n702), .B1(new_n691), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n667), .A2(new_n672), .A3(new_n675), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n675), .B1(new_n667), .B2(new_n672), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n739), .A2(new_n742), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n839), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n677), .A2(KEYINPUT52), .A3(new_n743), .A4(new_n843), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n376), .A2(new_n610), .B1(new_n654), .B2(new_n656), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n548), .A2(new_n625), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n623), .A2(new_n470), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n624), .A2(new_n631), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n618), .A2(new_n621), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n714), .A2(new_n717), .A3(new_n719), .A4(new_n731), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n805), .A2(new_n653), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n642), .A2(new_n470), .A3(new_n433), .A4(new_n670), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n609), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n667), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n749), .A2(new_n750), .A3(new_n700), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n728), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n763), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n859), .A2(new_n759), .A3(new_n760), .A4(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n838), .B1(new_n850), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n867), .A2(KEYINPUT107), .A3(new_n856), .A4(new_n851), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT107), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n376), .A2(new_n671), .A3(new_n752), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n667), .A2(new_n862), .B1(new_n728), .B2(new_n864), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n860), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n872), .B1(new_n857), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n848), .A2(KEYINPUT105), .A3(new_n849), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT105), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n879), .B(new_n839), .C1(new_n846), .C2(new_n847), .ZN(new_n880));
  INV_X1    g694(.A(new_n757), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n881), .A2(new_n838), .A3(new_n858), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n877), .A2(new_n878), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n869), .A2(new_n870), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n850), .A2(new_n868), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT53), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT106), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(KEYINPUT106), .A3(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n878), .A2(new_n880), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n838), .B1(new_n890), .B2(new_n868), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n884), .B1(new_n892), .B2(KEYINPUT54), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n828), .A2(new_n837), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(G952), .A2(G953), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n797), .B1(new_n894), .B2(new_n895), .ZN(G75));
  NOR2_X1   g710(.A1(new_n223), .A2(G952), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT116), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n238), .B1(new_n869), .B2(new_n883), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n899), .B2(G210), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n517), .A2(new_n529), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n527), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT113), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT55), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n898), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n899), .A2(G210), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT114), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n905), .A2(KEYINPUT115), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n905), .A2(KEYINPUT115), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT56), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n906), .B1(new_n908), .B2(new_n911), .ZN(G51));
  NAND2_X1  g726(.A1(new_n869), .A2(new_n883), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n869), .A2(new_n883), .A3(new_n870), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n552), .B(KEYINPUT57), .Z(new_n918));
  OAI21_X1  g732(.A(new_n706), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n899), .A2(new_n767), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n897), .B1(new_n919), .B2(new_n920), .ZN(G54));
  AND3_X1   g735(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n419), .A2(new_n421), .ZN(new_n923));
  OAI22_X1  g737(.A1(new_n922), .A2(new_n923), .B1(G952), .B2(new_n223), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT117), .ZN(G60));
  XNOR2_X1  g740(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n629), .B1(new_n893), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n898), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n629), .A2(new_n929), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n870), .B1(new_n869), .B2(new_n883), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n884), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT119), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n936), .B(new_n932), .C1(new_n884), .C2(new_n933), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n931), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n930), .B1(new_n938), .B2(KEYINPUT120), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n940), .B(new_n931), .C1(new_n935), .C2(new_n937), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT121), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n936), .B1(new_n916), .B2(new_n932), .ZN(new_n943));
  INV_X1    g757(.A(new_n937), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n898), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n938), .A2(KEYINPUT120), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .A4(new_n930), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n942), .A2(new_n949), .ZN(G63));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n898), .B1(new_n951), .B2(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n869), .B2(new_n883), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n955), .B2(new_n651), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n244), .B2(new_n955), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n951), .A2(KEYINPUT61), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G66));
  NOR2_X1   g773(.A1(new_n859), .A2(G953), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT123), .ZN(new_n961));
  OAI21_X1  g775(.A(G953), .B1(new_n477), .B2(new_n524), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n901), .B1(G898), .B2(new_n223), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(G69));
  AOI21_X1  g779(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT126), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(G900), .A2(G953), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n335), .A2(new_n341), .A3(new_n342), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n391), .A2(new_n392), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n729), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n376), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n763), .B1(new_n776), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n677), .A2(new_n703), .A3(new_n743), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n976), .A2(new_n784), .A3(new_n790), .A4(new_n978), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n979), .A2(new_n761), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n969), .B(new_n972), .C1(new_n980), .C2(G953), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT125), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n968), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n854), .A2(new_n853), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n680), .A2(new_n751), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n376), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n784), .A2(new_n790), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n697), .A2(new_n978), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(KEYINPUT62), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n990));
  AOI21_X1  g804(.A(G953), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n972), .B(KEYINPUT124), .Z(new_n992));
  OAI21_X1  g806(.A(new_n981), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n983), .B(new_n993), .Z(G72));
  INV_X1    g808(.A(new_n859), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n980), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n614), .A2(new_n238), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n371), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n689), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n989), .A2(new_n859), .A3(new_n990), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n999), .ZN(new_n1003));
  AND4_X1   g817(.A1(new_n371), .A2(new_n892), .A3(new_n1001), .A4(new_n999), .ZN(new_n1004));
  NOR4_X1   g818(.A1(new_n1000), .A2(new_n1003), .A3(new_n897), .A4(new_n1004), .ZN(G57));
endmodule


