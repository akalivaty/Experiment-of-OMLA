

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601;

  INV_X1 U326 ( .A(KEYINPUT47), .ZN(n400) );
  XNOR2_X1 U327 ( .A(n400), .B(KEYINPUT112), .ZN(n401) );
  XOR2_X1 U328 ( .A(G141GAT), .B(G22GAT), .Z(n449) );
  XNOR2_X1 U329 ( .A(n402), .B(n401), .ZN(n410) );
  XNOR2_X1 U330 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U331 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U332 ( .A(n467), .B(G190GAT), .ZN(n468) );
  XNOR2_X1 U333 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n295) );
  XNOR2_X1 U335 ( .A(G99GAT), .B(G218GAT), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U337 ( .A(G92GAT), .B(KEYINPUT77), .Z(n297) );
  XNOR2_X1 U338 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U340 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U341 ( .A(G43GAT), .B(G134GAT), .Z(n315) );
  XOR2_X1 U342 ( .A(G85GAT), .B(KEYINPUT71), .Z(n354) );
  XOR2_X1 U343 ( .A(G36GAT), .B(G190GAT), .Z(n421) );
  XOR2_X1 U344 ( .A(n354), .B(n421), .Z(n301) );
  NAND2_X1 U345 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n315), .B(n302), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U349 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n306) );
  XNOR2_X1 U350 ( .A(KEYINPUT75), .B(KEYINPUT65), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U352 ( .A(n308), .B(n307), .Z(n312) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n309) );
  XNOR2_X1 U354 ( .A(n309), .B(KEYINPUT7), .ZN(n371) );
  XNOR2_X1 U355 ( .A(G50GAT), .B(KEYINPUT73), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n310), .B(G162GAT), .ZN(n458) );
  XNOR2_X1 U357 ( .A(n371), .B(n458), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n565) );
  XOR2_X1 U359 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n314) );
  XNOR2_X1 U360 ( .A(G176GAT), .B(KEYINPUT83), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n319) );
  XOR2_X1 U362 ( .A(KEYINPUT20), .B(G190GAT), .Z(n317) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G127GAT), .Z(n381) );
  XNOR2_X1 U364 ( .A(n315), .B(n381), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U366 ( .A(n319), .B(n318), .Z(n321) );
  NAND2_X1 U367 ( .A1(G227GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n321), .B(n320), .ZN(n324) );
  XOR2_X1 U369 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n323) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n439) );
  XOR2_X1 U372 ( .A(n324), .B(n439), .Z(n332) );
  XOR2_X1 U373 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n326) );
  XNOR2_X1 U374 ( .A(KEYINPUT85), .B(KEYINPUT17), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U376 ( .A(n327), .B(KEYINPUT86), .Z(n329) );
  XNOR2_X1 U377 ( .A(G169GAT), .B(G183GAT), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n416) );
  XNOR2_X1 U379 ( .A(G99GAT), .B(G71GAT), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n330), .B(G120GAT), .ZN(n351) );
  XNOR2_X1 U381 ( .A(n416), .B(n351), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n532) );
  INV_X1 U383 ( .A(G148GAT), .ZN(n333) );
  NAND2_X1 U384 ( .A1(G78GAT), .A2(n333), .ZN(n336) );
  INV_X1 U385 ( .A(G78GAT), .ZN(n334) );
  NAND2_X1 U386 ( .A1(n334), .A2(G148GAT), .ZN(n335) );
  NAND2_X1 U387 ( .A1(n336), .A2(n335), .ZN(n338) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n448) );
  XNOR2_X1 U390 ( .A(n448), .B(KEYINPUT72), .ZN(n340) );
  AND2_X1 U391 ( .A1(G230GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n343) );
  XOR2_X1 U393 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n342) );
  XNOR2_X1 U394 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n341) );
  XOR2_X1 U395 ( .A(n342), .B(n341), .Z(n344) );
  NAND2_X1 U396 ( .A1(n343), .A2(n344), .ZN(n348) );
  INV_X1 U397 ( .A(n343), .ZN(n346) );
  INV_X1 U398 ( .A(n344), .ZN(n345) );
  NAND2_X1 U399 ( .A1(n346), .A2(n345), .ZN(n347) );
  NAND2_X1 U400 ( .A1(n348), .A2(n347), .ZN(n353) );
  XOR2_X1 U401 ( .A(G64GAT), .B(G92GAT), .Z(n350) );
  XNOR2_X1 U402 ( .A(G176GAT), .B(G204GAT), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n417) );
  XNOR2_X1 U404 ( .A(n351), .B(n417), .ZN(n352) );
  XOR2_X1 U405 ( .A(n353), .B(n352), .Z(n355) );
  XNOR2_X1 U406 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U407 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n382) );
  XNOR2_X1 U408 ( .A(n356), .B(n382), .ZN(n403) );
  XOR2_X1 U409 ( .A(KEYINPUT41), .B(n403), .Z(n560) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G15GAT), .Z(n358) );
  XNOR2_X1 U411 ( .A(G43GAT), .B(G197GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n377) );
  INV_X1 U413 ( .A(G8GAT), .ZN(n359) );
  NAND2_X1 U414 ( .A1(G1GAT), .A2(n359), .ZN(n362) );
  INV_X1 U415 ( .A(G1GAT), .ZN(n360) );
  NAND2_X1 U416 ( .A1(n360), .A2(G8GAT), .ZN(n361) );
  NAND2_X1 U417 ( .A1(n362), .A2(n361), .ZN(n392) );
  XNOR2_X1 U418 ( .A(n449), .B(n392), .ZN(n364) );
  XOR2_X1 U419 ( .A(G50GAT), .B(G36GAT), .Z(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U421 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n366) );
  XNOR2_X1 U422 ( .A(G169GAT), .B(KEYINPUT30), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n370) );
  AND2_X1 U425 ( .A1(G229GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n375) );
  XNOR2_X1 U427 ( .A(n371), .B(KEYINPUT68), .ZN(n373) );
  INV_X1 U428 ( .A(KEYINPUT67), .ZN(n372) );
  XOR2_X1 U429 ( .A(n377), .B(n376), .Z(n569) );
  INV_X1 U430 ( .A(n569), .ZN(n586) );
  NOR2_X1 U431 ( .A1(n560), .A2(n586), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n378), .B(KEYINPUT46), .ZN(n397) );
  XOR2_X1 U433 ( .A(G78GAT), .B(G155GAT), .Z(n380) );
  XNOR2_X1 U434 ( .A(G22GAT), .B(G211GAT), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n396) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n384) );
  NAND2_X1 U437 ( .A1(G231GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U439 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n386) );
  XNOR2_X1 U440 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U442 ( .A(n388), .B(n387), .Z(n394) );
  XOR2_X1 U443 ( .A(G64GAT), .B(KEYINPUT12), .Z(n390) );
  XNOR2_X1 U444 ( .A(G183GAT), .B(G71GAT), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U448 ( .A(n396), .B(n395), .ZN(n577) );
  NOR2_X1 U449 ( .A1(n397), .A2(n577), .ZN(n398) );
  XNOR2_X1 U450 ( .A(n398), .B(KEYINPUT111), .ZN(n399) );
  NOR2_X1 U451 ( .A1(n565), .A2(n399), .ZN(n402) );
  BUF_X1 U452 ( .A(n403), .Z(n591) );
  INV_X1 U453 ( .A(n577), .ZN(n596) );
  XOR2_X1 U454 ( .A(n565), .B(KEYINPUT102), .Z(n404) );
  XNOR2_X1 U455 ( .A(KEYINPUT36), .B(n404), .ZN(n598) );
  NOR2_X1 U456 ( .A1(n596), .A2(n598), .ZN(n406) );
  XNOR2_X1 U457 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n405) );
  XNOR2_X1 U458 ( .A(n406), .B(n405), .ZN(n407) );
  NAND2_X1 U459 ( .A1(n591), .A2(n407), .ZN(n408) );
  NOR2_X1 U460 ( .A1(n408), .A2(n569), .ZN(n409) );
  NOR2_X1 U461 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U462 ( .A(KEYINPUT48), .B(n411), .ZN(n539) );
  XNOR2_X1 U463 ( .A(G211GAT), .B(KEYINPUT89), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n412), .B(KEYINPUT21), .ZN(n413) );
  XOR2_X1 U465 ( .A(n413), .B(KEYINPUT88), .Z(n415) );
  XNOR2_X1 U466 ( .A(G197GAT), .B(G218GAT), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n453) );
  XNOR2_X1 U468 ( .A(n416), .B(n453), .ZN(n425) );
  XOR2_X1 U469 ( .A(n417), .B(KEYINPUT94), .Z(n419) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U472 ( .A(n420), .B(KEYINPUT93), .Z(n423) );
  XNOR2_X1 U473 ( .A(G8GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U475 ( .A(n425), .B(n424), .ZN(n507) );
  XNOR2_X1 U476 ( .A(n507), .B(KEYINPUT119), .ZN(n426) );
  NOR2_X1 U477 ( .A1(n539), .A2(n426), .ZN(n427) );
  XNOR2_X1 U478 ( .A(n427), .B(KEYINPUT54), .ZN(n581) );
  XOR2_X1 U479 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n429) );
  XNOR2_X1 U480 ( .A(G57GAT), .B(KEYINPUT6), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n447) );
  XOR2_X1 U482 ( .A(G148GAT), .B(G134GAT), .Z(n431) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(G141GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U485 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n433) );
  XNOR2_X1 U486 ( .A(G120GAT), .B(G127GAT), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U488 ( .A(n435), .B(n434), .Z(n441) );
  XOR2_X1 U489 ( .A(G85GAT), .B(G162GAT), .Z(n437) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U494 ( .A(n442), .B(KEYINPUT92), .Z(n445) );
  XNOR2_X1 U495 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n443), .B(KEYINPUT2), .ZN(n457) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(n457), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n580) );
  INV_X1 U500 ( .A(n580), .ZN(n504) );
  XOR2_X1 U501 ( .A(n448), .B(G204GAT), .Z(n451) );
  XNOR2_X1 U502 ( .A(n449), .B(KEYINPUT24), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n453), .B(n452), .ZN(n462) );
  XOR2_X1 U505 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n455) );
  NAND2_X1 U506 ( .A1(G228GAT), .A2(G233GAT), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U508 ( .A(n456), .B(KEYINPUT90), .Z(n460) );
  XNOR2_X1 U509 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U510 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U511 ( .A(n462), .B(n461), .ZN(n476) );
  NOR2_X1 U512 ( .A1(n504), .A2(n476), .ZN(n463) );
  AND2_X1 U513 ( .A1(n581), .A2(n463), .ZN(n464) );
  XNOR2_X1 U514 ( .A(n464), .B(KEYINPUT55), .ZN(n465) );
  NOR2_X1 U515 ( .A1(n532), .A2(n465), .ZN(n466) );
  XNOR2_X1 U516 ( .A(KEYINPUT120), .B(n466), .ZN(n578) );
  NAND2_X1 U517 ( .A1(n565), .A2(n578), .ZN(n469) );
  XOR2_X1 U518 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n467) );
  XNOR2_X1 U519 ( .A(n476), .B(KEYINPUT28), .ZN(n543) );
  XOR2_X1 U520 ( .A(n507), .B(KEYINPUT27), .Z(n478) );
  NOR2_X1 U521 ( .A1(n580), .A2(n478), .ZN(n470) );
  XNOR2_X1 U522 ( .A(n470), .B(KEYINPUT95), .ZN(n538) );
  NOR2_X1 U523 ( .A1(n543), .A2(n538), .ZN(n471) );
  XOR2_X1 U524 ( .A(KEYINPUT96), .B(n471), .Z(n473) );
  XNOR2_X1 U525 ( .A(n532), .B(KEYINPUT87), .ZN(n472) );
  NOR2_X1 U526 ( .A1(n473), .A2(n472), .ZN(n483) );
  INV_X1 U527 ( .A(n507), .ZN(n528) );
  NOR2_X1 U528 ( .A1(n532), .A2(n528), .ZN(n474) );
  NOR2_X1 U529 ( .A1(n476), .A2(n474), .ZN(n475) );
  XOR2_X1 U530 ( .A(KEYINPUT25), .B(n475), .Z(n480) );
  NAND2_X1 U531 ( .A1(n476), .A2(n532), .ZN(n477) );
  XNOR2_X1 U532 ( .A(n477), .B(KEYINPUT26), .ZN(n583) );
  NOR2_X1 U533 ( .A1(n583), .A2(n478), .ZN(n479) );
  NOR2_X1 U534 ( .A1(n480), .A2(n479), .ZN(n481) );
  NOR2_X1 U535 ( .A1(n504), .A2(n481), .ZN(n482) );
  NOR2_X1 U536 ( .A1(n483), .A2(n482), .ZN(n498) );
  NOR2_X1 U537 ( .A1(n565), .A2(n596), .ZN(n484) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U539 ( .A1(n498), .A2(n485), .ZN(n486) );
  XOR2_X1 U540 ( .A(KEYINPUT97), .B(n486), .Z(n516) );
  AND2_X1 U541 ( .A1(n569), .A2(n591), .ZN(n502) );
  NAND2_X1 U542 ( .A1(n516), .A2(n502), .ZN(n487) );
  XNOR2_X1 U543 ( .A(KEYINPUT98), .B(n487), .ZN(n495) );
  NOR2_X1 U544 ( .A1(n495), .A2(n580), .ZN(n491) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(KEYINPUT100), .ZN(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT99), .B(n489), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  NOR2_X1 U549 ( .A1(n495), .A2(n528), .ZN(n492) );
  XOR2_X1 U550 ( .A(G8GAT), .B(n492), .Z(G1325GAT) );
  XNOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n494) );
  NOR2_X1 U552 ( .A1(n532), .A2(n495), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n497) );
  INV_X1 U555 ( .A(n543), .ZN(n535) );
  NOR2_X1 U556 ( .A1(n535), .A2(n495), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .Z(n506) );
  NOR2_X1 U559 ( .A1(n598), .A2(n498), .ZN(n499) );
  NAND2_X1 U560 ( .A1(n596), .A2(n499), .ZN(n500) );
  XNOR2_X1 U561 ( .A(KEYINPUT103), .B(n500), .ZN(n501) );
  XOR2_X1 U562 ( .A(KEYINPUT37), .B(n501), .Z(n526) );
  NAND2_X1 U563 ( .A1(n526), .A2(n502), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT38), .B(n503), .Z(n514) );
  NAND2_X1 U565 ( .A1(n504), .A2(n514), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n514), .A2(n507), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n508), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n510) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(n513) );
  INV_X1 U572 ( .A(n532), .ZN(n540) );
  NAND2_X1 U573 ( .A1(n514), .A2(n540), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(KEYINPUT104), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(G1330GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n543), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n515), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U578 ( .A(n560), .B(KEYINPUT107), .ZN(n574) );
  AND2_X1 U579 ( .A1(n586), .A2(n574), .ZN(n525) );
  NAND2_X1 U580 ( .A1(n516), .A2(n525), .ZN(n521) );
  NOR2_X1 U581 ( .A1(n580), .A2(n521), .ZN(n517) );
  XOR2_X1 U582 ( .A(KEYINPUT42), .B(n517), .Z(n518) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(n518), .ZN(G1332GAT) );
  NOR2_X1 U584 ( .A1(n528), .A2(n521), .ZN(n519) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n519), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n532), .A2(n521), .ZN(n520) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n535), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n534) );
  NOR2_X1 U593 ( .A1(n580), .A2(n534), .ZN(n527) );
  XOR2_X1 U594 ( .A(G85GAT), .B(n527), .Z(G1336GAT) );
  NOR2_X1 U595 ( .A1(n528), .A2(n534), .ZN(n530) );
  XNOR2_X1 U596 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  NOR2_X1 U599 ( .A1(n532), .A2(n534), .ZN(n533) );
  XOR2_X1 U600 ( .A(G99GAT), .B(n533), .Z(G1338GAT) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(n536), .Z(n537) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n545) );
  NOR2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n557) );
  NAND2_X1 U606 ( .A1(n557), .A2(n540), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT113), .B(n541), .Z(n542) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n569), .A2(n553), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n547) );
  NAND2_X1 U612 ( .A1(n553), .A2(n574), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT115), .Z(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n551) );
  NAND2_X1 U617 ( .A1(n553), .A2(n577), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U620 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n565), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  INV_X1 U623 ( .A(n583), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n566) );
  NOR2_X1 U625 ( .A1(n586), .A2(n566), .ZN(n558) );
  XOR2_X1 U626 ( .A(G141GAT), .B(n558), .Z(n559) );
  XNOR2_X1 U627 ( .A(KEYINPUT118), .B(n559), .ZN(G1344GAT) );
  NOR2_X1 U628 ( .A1(n560), .A2(n566), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  NOR2_X1 U632 ( .A1(n596), .A2(n566), .ZN(n564) );
  XOR2_X1 U633 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  INV_X1 U634 ( .A(n565), .ZN(n567) );
  NOR2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U636 ( .A(G162GAT), .B(n568), .Z(G1347GAT) );
  NAND2_X1 U637 ( .A1(n578), .A2(n569), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n570), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n572) );
  XNOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U642 ( .A(KEYINPUT121), .B(n573), .Z(n576) );
  NAND2_X1 U643 ( .A1(n574), .A2(n578), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n576), .B(n575), .ZN(G1349GAT) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U647 ( .A(KEYINPUT124), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n599) );
  NOR2_X1 U651 ( .A1(n586), .A2(n599), .ZN(n590) );
  XOR2_X1 U652 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n588) );
  XNOR2_X1 U653 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1352GAT) );
  NOR2_X1 U656 ( .A1(n591), .A2(n599), .ZN(n595) );
  XOR2_X1 U657 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n593) );
  XNOR2_X1 U658 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n592) );
  XNOR2_X1 U659 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U660 ( .A(n595), .B(n594), .ZN(G1353GAT) );
  NOR2_X1 U661 ( .A1(n596), .A2(n599), .ZN(n597) );
  XOR2_X1 U662 ( .A(G211GAT), .B(n597), .Z(G1354GAT) );
  NOR2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U664 ( .A(KEYINPUT62), .B(n600), .Z(n601) );
  XNOR2_X1 U665 ( .A(G218GAT), .B(n601), .ZN(G1355GAT) );
endmodule

